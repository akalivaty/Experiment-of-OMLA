//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT32), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT11), .A2(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT65), .A2(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT11), .A2(G134), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT11), .A2(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G137), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n197), .A2(new_n198), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT65), .A2(G137), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT65), .A2(G137), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n203), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n198), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT71), .B1(new_n202), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n197), .A2(new_n201), .A3(new_n198), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT71), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n194), .A2(new_n196), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n207), .B1(new_n213), .B2(new_n203), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n211), .B(new_n212), .C1(new_n214), .C2(new_n198), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT64), .A2(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(G143), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n220), .A2(G128), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT68), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n225), .B1(new_n220), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n217), .A2(G143), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n218), .A2(new_n219), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(new_n222), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n224), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n210), .A2(new_n215), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n220), .A2(new_n238), .A3(new_n223), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT0), .B(G128), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT64), .A2(G146), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT64), .A2(G146), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n222), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n243), .B2(new_n232), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n198), .A2(KEYINPUT66), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n197), .B2(new_n201), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n197), .A2(new_n246), .A3(new_n201), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G119), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT70), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n253), .A3(G116), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G113), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT2), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G113), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n254), .A2(new_n256), .A3(new_n262), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n237), .A2(new_n249), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT67), .B1(new_n202), .B2(new_n209), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n211), .B(new_n271), .C1(new_n214), .C2(new_n198), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n236), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n267), .B1(new_n273), .B2(new_n249), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT28), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n237), .A2(new_n249), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n237), .B2(new_n249), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n278), .A2(new_n279), .A3(new_n266), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n275), .B1(new_n280), .B2(KEYINPUT28), .ZN(new_n281));
  NOR2_X1   g095(.A1(G237), .A2(G953), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G210), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT27), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G101), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT75), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n237), .A2(new_n249), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n266), .B1(new_n289), .B2(KEYINPUT74), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT28), .B1(new_n290), .B2(new_n277), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n273), .A2(new_n249), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n266), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n294), .B2(new_n268), .ZN(new_n295));
  OAI211_X1 g109(.A(KEYINPUT75), .B(new_n287), .C1(new_n291), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n288), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n237), .A2(new_n249), .A3(KEYINPUT30), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n237), .A2(new_n249), .A3(KEYINPUT72), .A4(KEYINPUT30), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n293), .A2(KEYINPUT69), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT69), .B1(new_n293), .B2(new_n304), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n303), .B(new_n266), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n268), .A2(KEYINPUT73), .A3(new_n286), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(KEYINPUT31), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n293), .A2(new_n304), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n314), .A2(new_n305), .B1(new_n301), .B2(new_n302), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n309), .B1(new_n315), .B2(new_n266), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n191), .B1(new_n298), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n289), .A2(new_n266), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n292), .B1(new_n320), .B2(new_n268), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n291), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n287), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(G902), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n275), .B(new_n286), .C1(new_n280), .C2(KEYINPUT28), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n323), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n286), .B1(new_n308), .B2(new_n268), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G472), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n309), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n308), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n333), .A2(KEYINPUT31), .B1(new_n308), .B2(new_n310), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n287), .B1(new_n291), .B2(new_n295), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n296), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT32), .B1(new_n339), .B2(new_n188), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n187), .B1(new_n331), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n188), .B1(new_n298), .B2(new_n318), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n190), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n339), .A2(new_n191), .B1(new_n329), .B2(G472), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT76), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  INV_X1    g160(.A(G953), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n347), .A2(G221), .A3(G234), .ZN(new_n348));
  XOR2_X1   g162(.A(new_n346), .B(new_n348), .Z(new_n349));
  INV_X1    g163(.A(G140), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G125), .ZN(new_n351));
  INV_X1    g165(.A(G125), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G140), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n354), .A2(new_n218), .A3(new_n219), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT78), .ZN(new_n356));
  OR3_X1    g170(.A1(new_n352), .A2(KEYINPUT78), .A3(G140), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT16), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT16), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n351), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n355), .B1(new_n361), .B2(G146), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT23), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT70), .B(G119), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(G128), .ZN(new_n365));
  INV_X1    g179(.A(G110), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n251), .A2(new_n253), .A3(G128), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n225), .A2(KEYINPUT23), .A3(G119), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n365), .A2(new_n366), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(G119), .B2(new_n225), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n367), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n364), .A2(new_n370), .A3(G128), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT24), .B(G110), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n362), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n362), .A2(new_n376), .A3(KEYINPUT79), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n361), .A2(G146), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n358), .A2(new_n217), .A3(new_n360), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n372), .A2(new_n373), .ZN(new_n385));
  INV_X1    g199(.A(new_n374), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G110), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n349), .B1(new_n381), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n362), .A2(new_n376), .A3(KEYINPUT79), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT79), .B1(new_n362), .B2(new_n376), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n390), .B(new_n349), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  INV_X1    g211(.A(G902), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(G234), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n404));
  INV_X1    g218(.A(new_n349), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n398), .A3(new_n394), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT25), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT81), .B1(new_n407), .B2(new_n408), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT81), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n396), .A2(new_n413), .A3(KEYINPUT25), .A4(new_n398), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(KEYINPUT80), .A3(new_n408), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n411), .A2(new_n412), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n403), .B1(new_n399), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n341), .A2(new_n345), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G214), .B1(G237), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G210), .B1(G237), .B2(G902), .ZN(new_n421));
  OR2_X1    g235(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n254), .A2(new_n256), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n364), .A2(G116), .A3(new_n422), .A4(new_n423), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G113), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n428));
  INV_X1    g242(.A(G104), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(G107), .ZN(new_n430));
  INV_X1    g244(.A(G107), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT3), .A3(G104), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G101), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n431), .B2(G104), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(KEYINPUT83), .A3(G107), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n433), .A2(new_n434), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n429), .A2(G107), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n431), .A2(G104), .ZN(new_n440));
  OAI21_X1  g254(.A(G101), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n427), .A2(new_n265), .A3(new_n438), .A4(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n430), .A2(new_n432), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n436), .A2(new_n437), .ZN(new_n444));
  OAI21_X1  g258(.A(G101), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n445), .A2(KEYINPUT4), .A3(new_n438), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT4), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(G101), .C1(new_n443), .C2(new_n444), .ZN(new_n448));
  INV_X1    g262(.A(new_n265), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n262), .B1(new_n254), .B2(new_n256), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n442), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G122), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT87), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n445), .A2(KEYINPUT4), .A3(new_n438), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n266), .A3(new_n448), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n454), .B1(new_n459), .B2(new_n442), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n453), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G125), .B1(new_n239), .B2(new_n244), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n352), .B(new_n224), .C1(new_n231), .C2(new_n235), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT88), .B(G125), .C1(new_n239), .C2(new_n244), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n347), .A2(G224), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n436), .A2(new_n437), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n434), .B1(new_n473), .B2(new_n433), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n447), .A2(new_n474), .B1(new_n264), .B2(new_n265), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n438), .A2(new_n265), .A3(new_n441), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n475), .A2(new_n458), .B1(new_n477), .B2(new_n427), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n453), .B1(new_n478), .B2(new_n454), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n452), .A2(new_n455), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n454), .B(new_n442), .C1(new_n446), .C2(new_n451), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT6), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n483), .A2(KEYINPUT86), .A3(new_n460), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n463), .B(new_n471), .C1(new_n481), .C2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n454), .B(KEYINPUT8), .ZN(new_n486));
  OAI21_X1  g300(.A(G113), .B1(new_n254), .B2(new_n424), .ZN(new_n487));
  INV_X1    g301(.A(new_n257), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(KEYINPUT5), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(new_n476), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n427), .A2(new_n265), .B1(new_n438), .B2(new_n441), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n466), .A2(new_n467), .A3(new_n470), .A4(new_n468), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n464), .A2(new_n467), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n470), .B1(KEYINPUT89), .B2(KEYINPUT7), .ZN(new_n498));
  AND2_X1   g312(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n496), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  AOI211_X1 g316(.A(KEYINPUT90), .B(new_n500), .C1(new_n464), .C2(new_n467), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT91), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n497), .A2(new_n501), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT90), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n496), .A3(new_n501), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n468), .A2(new_n467), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n512), .A2(KEYINPUT7), .A3(new_n470), .A4(new_n466), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n509), .A2(new_n510), .A3(new_n513), .A4(new_n492), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n505), .A2(new_n514), .A3(new_n482), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n485), .A2(new_n515), .A3(new_n398), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n421), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT86), .B1(new_n483), .B2(new_n460), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n480), .A2(new_n472), .A3(KEYINPUT6), .A4(new_n482), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n519), .A2(new_n520), .B1(new_n457), .B2(new_n462), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n521), .B2(new_n471), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(KEYINPUT92), .A3(new_n515), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n485), .A2(new_n515), .A3(new_n398), .A4(new_n421), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n420), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n282), .A2(G143), .A3(G214), .ZN(new_n529));
  AOI21_X1  g343(.A(G143), .B1(new_n282), .B2(G214), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT93), .ZN(new_n532));
  INV_X1    g346(.A(G237), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n347), .A3(G214), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n222), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n282), .A2(G143), .A3(G214), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT93), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(G131), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n528), .B1(new_n532), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n527), .B1(new_n384), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n538), .B1(new_n537), .B2(G131), .ZN(new_n542));
  AOI211_X1 g356(.A(KEYINPUT93), .B(new_n198), .C1(new_n535), .C2(new_n536), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT17), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n544), .A2(KEYINPUT94), .A3(new_n382), .A4(new_n383), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n537), .A2(G131), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n528), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n541), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G113), .B(G122), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(new_n429), .ZN(new_n551));
  NAND2_X1  g365(.A1(KEYINPUT18), .A2(G131), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n537), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n356), .A2(new_n357), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(new_n217), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n355), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n549), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n551), .B1(new_n549), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n398), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(KEYINPUT96), .B(new_n398), .C1(new_n557), .C2(new_n558), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(G475), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n255), .A2(G122), .ZN(new_n564));
  INV_X1    g378(.A(G122), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G116), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT97), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n567), .B1(new_n564), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n431), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n565), .A2(G116), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n255), .A2(G122), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT97), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(G107), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n222), .A2(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n225), .A2(G143), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n203), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n222), .A2(KEYINPUT13), .A3(G128), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n580), .A2(new_n578), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  AOI211_X1 g398(.A(KEYINPUT98), .B(KEYINPUT13), .C1(new_n222), .C2(G128), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G134), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n576), .A2(new_n579), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n573), .A2(new_n574), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n577), .A2(new_n578), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G134), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n589), .A2(new_n431), .B1(new_n579), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT14), .B1(new_n565), .B2(G116), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT99), .B1(new_n593), .B2(new_n571), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT14), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n255), .B2(G122), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n564), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n564), .B2(KEYINPUT14), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n571), .A2(KEYINPUT100), .A3(new_n595), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n594), .A2(new_n598), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G107), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n592), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n588), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT9), .B(G234), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n606), .A2(new_n397), .A3(G953), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n588), .A2(new_n604), .A3(new_n607), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n605), .A2(KEYINPUT101), .A3(new_n608), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n612), .A2(new_n613), .A3(new_n398), .A4(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT15), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n615), .A2(new_n616), .A3(G478), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(G478), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n398), .A3(new_n614), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT102), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n615), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G952), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(G953), .ZN(new_n624));
  NAND2_X1  g438(.A1(G234), .A2(G237), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(G902), .A3(G953), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT21), .B(G898), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n549), .A2(new_n551), .A3(new_n556), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n354), .A2(KEYINPUT19), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n554), .B2(KEYINPUT19), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n382), .B1(new_n635), .B2(new_n234), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n556), .B1(new_n636), .B2(new_n547), .ZN(new_n637));
  INV_X1    g451(.A(new_n551), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(G475), .A2(G902), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT95), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT20), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT20), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n640), .A2(new_n645), .A3(new_n642), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n563), .A2(new_n622), .A3(new_n632), .A4(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(G221), .B1(new_n606), .B2(G902), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(G110), .B(G140), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n347), .A2(G227), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n248), .A2(new_n247), .ZN(new_n655));
  INV_X1    g469(.A(new_n224), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n225), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n220), .B2(new_n223), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n438), .B(new_n441), .C1(new_n656), .C2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n458), .A2(new_n245), .A3(new_n448), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n438), .A2(KEYINPUT10), .A3(new_n441), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n236), .ZN(new_n664));
  AND4_X1   g478(.A1(new_n655), .A2(new_n661), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n659), .A2(new_n660), .B1(new_n663), .B2(new_n236), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n655), .B1(new_n666), .B2(new_n662), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n654), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n438), .A2(new_n441), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n669), .B(new_n224), .C1(new_n235), .C2(new_n231), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n659), .ZN(new_n671));
  INV_X1    g485(.A(new_n655), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT12), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT12), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n671), .A2(new_n675), .A3(new_n672), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n666), .A2(new_n655), .A3(new_n662), .ZN(new_n677));
  INV_X1    g491(.A(new_n654), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n674), .A2(new_n676), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(G469), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n398), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT84), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(G902), .B1(new_n668), .B2(new_n679), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(KEYINPUT84), .A3(new_n681), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n654), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n672), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n677), .A3(new_n678), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n681), .B1(new_n693), .B2(new_n398), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n651), .B1(new_n687), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n526), .A2(new_n649), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n418), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n434), .ZN(G3));
  NAND2_X1  g513(.A1(new_n563), .A2(new_n647), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT33), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n612), .A2(new_n701), .A3(new_n614), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n609), .A2(KEYINPUT33), .A3(new_n611), .ZN(new_n703));
  INV_X1    g517(.A(G478), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(G902), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n702), .A2(KEYINPUT103), .A3(new_n703), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n619), .A2(new_n704), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n700), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n421), .B1(new_n522), .B2(new_n515), .ZN(new_n714));
  INV_X1    g528(.A(new_n525), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n419), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n713), .A2(new_n716), .A3(new_n631), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n416), .A2(new_n399), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n401), .B(KEYINPUT82), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND4_X1   g534(.A1(KEYINPUT84), .A2(new_n680), .A3(new_n681), .A4(new_n398), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT84), .B1(new_n685), .B2(new_n681), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n650), .B1(new_n723), .B2(new_n694), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n339), .A2(new_n398), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n726), .A2(G472), .B1(new_n188), .B2(new_n339), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n717), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT34), .B(G104), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G6));
  NAND2_X1  g544(.A1(new_n621), .A2(new_n618), .ZN(new_n731));
  INV_X1    g545(.A(new_n617), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n563), .A3(new_n647), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n631), .B(KEYINPUT104), .Z(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n716), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n725), .A2(new_n737), .A3(new_n727), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT35), .B(G107), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G9));
  NOR2_X1   g554(.A1(new_n405), .A2(KEYINPUT36), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n404), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n400), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n416), .B2(new_n399), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n648), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n727), .A2(new_n746), .A3(new_n526), .A4(new_n696), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT37), .B(G110), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G12));
  INV_X1    g563(.A(G900), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n629), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n626), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n733), .A2(new_n563), .A3(new_n647), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT105), .ZN(new_n754));
  INV_X1    g568(.A(G475), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n549), .A2(new_n556), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n638), .ZN(new_n757));
  AOI21_X1  g571(.A(G902), .B1(new_n757), .B2(new_n633), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n755), .B1(new_n758), .B2(KEYINPUT96), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n759), .A2(new_n561), .B1(new_n644), .B2(new_n646), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n733), .A4(new_n752), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n724), .A2(new_n716), .A3(new_n745), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n341), .A3(new_n345), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G128), .ZN(G30));
  XNOR2_X1  g580(.A(new_n752), .B(KEYINPUT39), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n696), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT107), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT40), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n524), .A2(new_n525), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT38), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n700), .A2(new_n733), .A3(new_n419), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n287), .B1(new_n308), .B2(new_n268), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n320), .A2(new_n268), .A3(new_n287), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n398), .ZN(new_n779));
  OAI21_X1  g593(.A(G472), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n343), .A3(new_n319), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n718), .A2(new_n743), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n769), .A2(new_n770), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n771), .A2(new_n776), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G143), .ZN(G45));
  INV_X1    g603(.A(new_n752), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n713), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n764), .A2(new_n341), .A3(new_n345), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G146), .ZN(G48));
  AOI21_X1  g607(.A(new_n681), .B1(new_n680), .B2(new_n398), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n687), .A2(new_n650), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n720), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n341), .A2(new_n717), .A3(new_n345), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT41), .B(G113), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G15));
  NAND4_X1  g614(.A1(new_n341), .A2(new_n345), .A3(new_n737), .A4(new_n797), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G116), .ZN(G18));
  NAND3_X1  g616(.A1(new_n341), .A2(new_n345), .A3(new_n746), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n651), .B(new_n794), .C1(new_n684), .C2(new_n686), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n805));
  INV_X1    g619(.A(new_n421), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n516), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n420), .B1(new_n807), .B2(new_n525), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n804), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n805), .B1(new_n804), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n803), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G119), .ZN(G21));
  NOR2_X1   g627(.A1(new_n714), .A2(new_n715), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n775), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n322), .A2(new_n286), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n188), .B1(new_n318), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(G902), .B1(new_n334), .B2(new_n338), .ZN(new_n818));
  INV_X1    g632(.A(G472), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n796), .A2(new_n736), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n815), .A2(new_n821), .A3(new_n822), .A4(new_n417), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G122), .ZN(G24));
  NOR2_X1   g638(.A1(new_n820), .A2(new_n745), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n825), .B(new_n791), .C1(new_n809), .C2(new_n810), .ZN(new_n826));
  XOR2_X1   g640(.A(KEYINPUT109), .B(G125), .Z(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(G27));
  OAI21_X1  g642(.A(new_n417), .B1(new_n331), .B2(new_n340), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n525), .A2(new_n419), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n518), .B2(new_n523), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n692), .A2(KEYINPUT110), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n691), .A2(new_n833), .A3(new_n677), .A4(new_n678), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n689), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n398), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(G469), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n651), .B1(new_n687), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n563), .A2(new_n647), .B1(new_n711), .B2(new_n708), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n831), .A2(new_n838), .A3(new_n839), .A4(new_n752), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT42), .B1(new_n829), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n831), .A2(new_n838), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT42), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n791), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n841), .B1(new_n418), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n198), .ZN(G33));
  NAND2_X1  g660(.A1(new_n763), .A2(new_n842), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n418), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(new_n203), .ZN(G36));
  INV_X1    g663(.A(KEYINPUT45), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n835), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n693), .A2(new_n850), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(G469), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(G469), .A2(G902), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(KEYINPUT111), .A3(KEYINPUT46), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n854), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT46), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n723), .B1(new_n858), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n650), .A3(new_n767), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT112), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n727), .A2(new_n745), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT113), .Z(new_n867));
  NAND2_X1  g681(.A1(new_n760), .A2(new_n712), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT43), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT43), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n760), .A2(new_n870), .A3(new_n712), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT44), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n865), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  INV_X1    g690(.A(new_n830), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n524), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(G137), .ZN(G39));
  NAND2_X1  g695(.A1(new_n791), .A2(new_n720), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n341), .B2(new_n345), .ZN(new_n883));
  INV_X1    g697(.A(new_n862), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n860), .B2(new_n856), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT47), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(new_n651), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT47), .B1(new_n863), .B2(new_n650), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n831), .B(new_n883), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(G140), .ZN(G42));
  NAND3_X1  g704(.A1(new_n417), .A2(new_n419), .A3(new_n650), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n687), .A2(new_n795), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n868), .B(new_n891), .C1(KEYINPUT49), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(KEYINPUT49), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT114), .Z(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n784), .A3(new_n774), .A4(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n341), .A2(new_n345), .A3(new_n696), .A4(new_n785), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n760), .A2(new_n622), .A3(new_n752), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT115), .B1(new_n878), .B2(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n700), .A2(new_n733), .A3(new_n790), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT115), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n831), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n418), .A2(new_n847), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT116), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n726), .A2(G472), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n785), .A3(new_n817), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n907), .B2(new_n840), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n825), .A2(new_n842), .A3(KEYINPUT116), .A4(new_n791), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n904), .A2(new_n910), .A3(new_n845), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n798), .B1(new_n418), .B2(new_n697), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n801), .B1(new_n803), .B2(new_n811), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n736), .B1(new_n713), .B2(new_n734), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n725), .A2(new_n914), .A3(new_n727), .A4(new_n526), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(new_n823), .A3(new_n747), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n912), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n765), .A2(new_n826), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT52), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n838), .A2(new_n752), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n783), .A2(new_n921), .A3(new_n815), .A4(new_n745), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n919), .A2(new_n920), .A3(new_n792), .A4(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n765), .A2(new_n792), .A3(new_n826), .A4(new_n922), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT52), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT53), .ZN(new_n926));
  INV_X1    g740(.A(new_n919), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(KEYINPUT52), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n918), .A2(new_n923), .A3(new_n925), .A4(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n911), .A2(new_n923), .A3(new_n917), .A4(new_n925), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n926), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT51), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n886), .B1(new_n885), .B2(new_n651), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n863), .A2(KEYINPUT47), .A3(new_n650), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n687), .A2(new_n651), .A3(new_n795), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n821), .A2(new_n417), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n869), .A2(new_n627), .A3(new_n871), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n878), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n831), .A2(new_n804), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n783), .A2(new_n946), .A3(new_n720), .A4(new_n626), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n700), .A2(new_n712), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n941), .A2(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n825), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n804), .A2(new_n420), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n773), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n942), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT50), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(KEYINPUT50), .A3(new_n942), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT117), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n945), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n952), .ZN(new_n962));
  INV_X1    g776(.A(new_n958), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT50), .B1(new_n954), .B2(new_n942), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n962), .B(new_n960), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n935), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n947), .A2(new_n839), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n968), .B(new_n624), .C1(new_n811), .C2(new_n943), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n941), .A2(new_n829), .A3(new_n946), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT48), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n935), .B1(new_n939), .B2(new_n944), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n969), .B(new_n971), .C1(new_n972), .C2(new_n959), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT53), .B1(new_n927), .B2(KEYINPUT52), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n931), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n930), .B1(new_n976), .B2(new_n932), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n934), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n623), .A2(new_n347), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT118), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n896), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT119), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT119), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n983), .B(new_n896), .C1(new_n978), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G75));
  AND2_X1   g799(.A1(new_n931), .A2(new_n926), .ZN(new_n986));
  INV_X1    g800(.A(new_n928), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n931), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n398), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(KEYINPUT120), .A3(G210), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT56), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n521), .B(new_n471), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT55), .Z(new_n994));
  NAND3_X1  g808(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT120), .B1(new_n990), .B2(G210), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n623), .A2(G953), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT121), .Z(new_n999));
  AOI21_X1  g813(.A(KEYINPUT56), .B1(new_n990), .B2(G210), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n994), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n997), .A2(new_n1001), .ZN(G51));
  INV_X1    g816(.A(new_n680), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT54), .B1(new_n986), .B2(new_n988), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n933), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n854), .B(KEYINPUT57), .Z(new_n1006));
  AOI21_X1  g820(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n853), .ZN(new_n1008));
  OAI211_X1 g822(.A(G902), .B(new_n1008), .C1(new_n986), .C2(new_n988), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT122), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n929), .A2(new_n932), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1012), .A2(KEYINPUT122), .A3(G902), .A4(new_n1008), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n999), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT123), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g831(.A(KEYINPUT123), .B(new_n999), .C1(new_n1007), .C2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(G54));
  INV_X1    g833(.A(new_n999), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n990), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1021));
  OR2_X1    g835(.A1(new_n1021), .A2(new_n640), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n640), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(G60));
  NAND2_X1  g838(.A1(new_n702), .A2(new_n703), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT124), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n934), .A2(new_n977), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G478), .A2(G902), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT59), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1026), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1005), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1030), .A2(new_n1020), .A3(new_n1031), .ZN(G63));
  NAND2_X1  g846(.A1(G217), .A2(G902), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT60), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n989), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n742), .ZN(new_n1036));
  OAI22_X1  g850(.A1(new_n989), .A2(new_n1034), .B1(new_n395), .B2(new_n391), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1036), .A2(new_n999), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT61), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(G66));
  INV_X1    g854(.A(G224), .ZN(new_n1041));
  OAI21_X1  g855(.A(G953), .B1(new_n630), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n917), .B2(G953), .ZN(new_n1043));
  INV_X1    g857(.A(new_n521), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1044), .B1(G898), .B2(new_n347), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n1043), .B(new_n1045), .ZN(G69));
  NOR3_X1   g860(.A1(new_n829), .A2(new_n814), .A3(new_n775), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n865), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(KEYINPUT125), .ZN(new_n1049));
  INV_X1    g863(.A(KEYINPUT125), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n865), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(new_n889), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n765), .A2(new_n792), .A3(new_n826), .ZN(new_n1054));
  NOR4_X1   g868(.A1(new_n1053), .A2(new_n845), .A3(new_n848), .A4(new_n1054), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n1052), .A2(new_n347), .A3(new_n1055), .A4(new_n880), .ZN(new_n1056));
  XOR2_X1   g870(.A(new_n315), .B(new_n635), .Z(new_n1057));
  OAI211_X1 g871(.A(new_n1056), .B(new_n1057), .C1(new_n750), .C2(new_n347), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n713), .A2(new_n734), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n769), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1059), .B1(new_n418), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g876(.A1(new_n875), .A2(new_n879), .B1(new_n831), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g877(.A(new_n1054), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n788), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT62), .Z(new_n1066));
  AOI21_X1  g880(.A(G953), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1058), .B1(new_n1067), .B2(new_n1057), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n347), .B1(G227), .B2(G900), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g884(.A(new_n1069), .ZN(new_n1071));
  OAI211_X1 g885(.A(new_n1058), .B(new_n1071), .C1(new_n1067), .C2(new_n1057), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1070), .A2(new_n1072), .ZN(G72));
  NAND3_X1  g887(.A1(new_n1063), .A2(new_n1066), .A3(new_n917), .ZN(new_n1074));
  NAND2_X1  g888(.A1(G472), .A2(G902), .ZN(new_n1075));
  XOR2_X1   g889(.A(new_n1075), .B(KEYINPUT63), .Z(new_n1076));
  NAND2_X1  g890(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g891(.A(new_n1020), .B1(new_n1077), .B2(new_n777), .ZN(new_n1078));
  NAND2_X1  g892(.A1(new_n976), .A2(new_n932), .ZN(new_n1079));
  INV_X1    g893(.A(new_n777), .ZN(new_n1080));
  NAND3_X1  g894(.A1(new_n308), .A2(new_n268), .A3(new_n287), .ZN(new_n1081));
  NAND4_X1  g895(.A1(new_n1079), .A2(new_n1080), .A3(new_n1076), .A4(new_n1081), .ZN(new_n1082));
  NAND4_X1  g896(.A1(new_n1052), .A2(new_n880), .A3(new_n1055), .A4(new_n917), .ZN(new_n1083));
  INV_X1    g897(.A(KEYINPUT126), .ZN(new_n1084));
  NAND3_X1  g898(.A1(new_n1083), .A2(new_n1084), .A3(new_n1076), .ZN(new_n1085));
  XNOR2_X1  g899(.A(new_n1081), .B(KEYINPUT127), .ZN(new_n1086));
  NAND2_X1  g900(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g901(.A(new_n1084), .B1(new_n1083), .B2(new_n1076), .ZN(new_n1088));
  OAI211_X1 g902(.A(new_n1078), .B(new_n1082), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g903(.A(new_n1089), .ZN(G57));
endmodule


