

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757;

  NAND2_X1 U373 ( .A1(n578), .A2(n664), .ZN(n660) );
  XNOR2_X1 U374 ( .A(n432), .B(n507), .ZN(n525) );
  INV_X1 U375 ( .A(G953), .ZN(n741) );
  NAND2_X1 U376 ( .A1(n392), .A2(n387), .ZN(n549) );
  XNOR2_X1 U377 ( .A(KEYINPUT110), .B(KEYINPUT63), .ZN(n351) );
  XOR2_X1 U378 ( .A(n636), .B(n635), .Z(n352) );
  XNOR2_X1 U379 ( .A(KEYINPUT62), .B(n641), .ZN(n353) );
  XNOR2_X1 U380 ( .A(n386), .B(n564), .ZN(n724) );
  BUF_X2 U381 ( .A(n382), .Z(n714) );
  NOR2_X2 U382 ( .A1(n702), .A2(n719), .ZN(n704) );
  XNOR2_X1 U383 ( .A(n408), .B(n438), .ZN(n751) );
  NOR2_X2 U384 ( .A1(n580), .A2(n565), .ZN(n431) );
  XOR2_X2 U385 ( .A(KEYINPUT38), .B(n611), .Z(n676) );
  XNOR2_X2 U386 ( .A(n583), .B(KEYINPUT1), .ZN(n661) );
  XNOR2_X2 U387 ( .A(n516), .B(n515), .ZN(n583) );
  NAND2_X1 U388 ( .A1(n436), .A2(n434), .ZN(n688) );
  INV_X1 U389 ( .A(KEYINPUT69), .ZN(n418) );
  INV_X1 U390 ( .A(KEYINPUT60), .ZN(n356) );
  XNOR2_X1 U391 ( .A(n358), .B(n351), .ZN(G57) );
  XNOR2_X1 U392 ( .A(n357), .B(n356), .ZN(G60) );
  XNOR2_X1 U393 ( .A(n713), .B(n712), .ZN(n355) );
  XNOR2_X1 U394 ( .A(n362), .B(KEYINPUT83), .ZN(n361) );
  NOR2_X1 U395 ( .A1(n563), .A2(n643), .ZN(n364) );
  XNOR2_X1 U396 ( .A(n428), .B(KEYINPUT40), .ZN(n640) );
  NAND2_X1 U397 ( .A1(n429), .A2(n653), .ZN(n428) );
  OR2_X1 U398 ( .A1(n689), .A2(n585), .ZN(n586) );
  AND2_X1 U399 ( .A1(n399), .A2(n442), .ZN(n398) );
  XNOR2_X1 U400 ( .A(n471), .B(n378), .ZN(n544) );
  AND2_X1 U401 ( .A1(n430), .A2(n579), .ZN(n572) );
  XNOR2_X1 U402 ( .A(n580), .B(n420), .ZN(n424) );
  XNOR2_X1 U403 ( .A(n506), .B(n505), .ZN(n739) );
  XNOR2_X1 U404 ( .A(n482), .B(KEYINPUT4), .ZN(n736) );
  XNOR2_X1 U405 ( .A(n369), .B(n374), .ZN(n531) );
  INV_X1 U406 ( .A(n719), .ZN(n354) );
  XNOR2_X1 U407 ( .A(G116), .B(G113), .ZN(n521) );
  INV_X1 U408 ( .A(G146), .ZN(n444) );
  XNOR2_X1 U409 ( .A(KEYINPUT79), .B(KEYINPUT17), .ZN(n448) );
  INV_X1 U410 ( .A(G125), .ZN(n445) );
  XOR2_X1 U411 ( .A(G113), .B(G104), .Z(n493) );
  XOR2_X1 U412 ( .A(G128), .B(G137), .Z(n374) );
  NOR2_X1 U413 ( .A1(n355), .A2(n719), .ZN(G63) );
  NAND2_X1 U414 ( .A1(n359), .A2(n354), .ZN(n357) );
  NAND2_X1 U415 ( .A1(n360), .A2(n354), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n637), .B(n352), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n642), .B(n353), .ZN(n360) );
  NAND2_X1 U418 ( .A1(n365), .A2(n361), .ZN(n386) );
  NAND2_X1 U419 ( .A1(n364), .A2(n363), .ZN(n362) );
  NAND2_X1 U420 ( .A1(n549), .A2(KEYINPUT44), .ZN(n363) );
  NAND2_X1 U421 ( .A1(n366), .A2(n548), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n547), .B(n542), .ZN(n366) );
  NOR2_X2 U423 ( .A1(n751), .A2(n754), .ZN(n547) );
  XNOR2_X1 U424 ( .A(n367), .B(n368), .ZN(n702) );
  NAND2_X1 U425 ( .A1(n705), .A2(G210), .ZN(n367) );
  XOR2_X1 U426 ( .A(n701), .B(n381), .Z(n368) );
  INV_X1 U427 ( .A(n656), .ZN(n403) );
  INV_X1 U428 ( .A(n437), .ZN(n407) );
  INV_X1 U429 ( .A(n424), .ZN(n419) );
  AND2_X1 U430 ( .A1(n402), .A2(n373), .ZN(n563) );
  NOR2_X1 U431 ( .A1(n577), .A2(n575), .ZN(n501) );
  XOR2_X1 U432 ( .A(G110), .B(G119), .Z(n369) );
  XOR2_X1 U433 ( .A(KEYINPUT98), .B(KEYINPUT9), .Z(n477) );
  XNOR2_X1 U434 ( .A(n736), .B(n454), .ZN(n507) );
  NOR2_X1 U435 ( .A1(n424), .A2(n546), .ZN(n435) );
  XNOR2_X1 U436 ( .A(n458), .B(n481), .ZN(n720) );
  XNOR2_X1 U437 ( .A(n456), .B(n518), .ZN(n458) );
  XNOR2_X1 U438 ( .A(n489), .B(KEYINPUT10), .ZN(n737) );
  XNOR2_X1 U439 ( .A(n739), .B(G146), .ZN(n432) );
  XNOR2_X1 U440 ( .A(n576), .B(KEYINPUT41), .ZN(n689) );
  NOR2_X1 U441 ( .A1(n575), .A2(n678), .ZN(n576) );
  NAND2_X1 U442 ( .A1(n591), .A2(n419), .ZN(n592) );
  XNOR2_X1 U443 ( .A(n443), .B(n538), .ZN(n539) );
  NOR2_X1 U444 ( .A1(n715), .A2(G902), .ZN(n414) );
  INV_X1 U445 ( .A(G137), .ZN(n504) );
  XOR2_X1 U446 ( .A(KEYINPUT78), .B(KEYINPUT18), .Z(n451) );
  XNOR2_X1 U447 ( .A(n431), .B(KEYINPUT30), .ZN(n430) );
  INV_X1 U448 ( .A(KEYINPUT22), .ZN(n426) );
  INV_X1 U449 ( .A(KEYINPUT6), .ZN(n420) );
  XNOR2_X1 U450 ( .A(n525), .B(n524), .ZN(n641) );
  NAND2_X1 U451 ( .A1(n631), .A2(n385), .ZN(n740) );
  XNOR2_X1 U452 ( .A(n417), .B(n416), .ZN(n532) );
  INV_X1 U453 ( .A(KEYINPUT8), .ZN(n416) );
  NAND2_X1 U454 ( .A1(n741), .A2(G234), .ZN(n417) );
  XNOR2_X1 U455 ( .A(KEYINPUT23), .B(KEYINPUT89), .ZN(n529) );
  XOR2_X1 U456 ( .A(G116), .B(G107), .Z(n457) );
  XNOR2_X1 U457 ( .A(G134), .B(KEYINPUT7), .ZN(n476) );
  XOR2_X1 U458 ( .A(KEYINPUT72), .B(G110), .Z(n512) );
  XNOR2_X1 U459 ( .A(G107), .B(G104), .ZN(n508) );
  XOR2_X1 U460 ( .A(G140), .B(KEYINPUT77), .Z(n509) );
  INV_X1 U461 ( .A(n659), .ZN(n427) );
  XNOR2_X1 U462 ( .A(n497), .B(n496), .ZN(n636) );
  XNOR2_X1 U463 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U464 ( .A(n490), .B(n737), .ZN(n497) );
  AND2_X1 U465 ( .A1(n638), .A2(G953), .ZN(n719) );
  NAND2_X1 U466 ( .A1(n603), .A2(n584), .ZN(n585) );
  INV_X1 U467 ( .A(n601), .ZN(n584) );
  AND2_X1 U468 ( .A1(n421), .A2(n560), .ZN(n595) );
  XNOR2_X1 U469 ( .A(n422), .B(KEYINPUT36), .ZN(n421) );
  AND2_X1 U470 ( .A1(n395), .A2(n393), .ZN(n392) );
  NOR2_X1 U471 ( .A1(n391), .A2(n389), .ZN(n388) );
  XNOR2_X1 U472 ( .A(n404), .B(KEYINPUT31), .ZN(n656) );
  NAND2_X1 U473 ( .A1(n406), .A2(n405), .ZN(n404) );
  INV_X1 U474 ( .A(KEYINPUT104), .ZN(n438) );
  INV_X1 U475 ( .A(n578), .ZN(n439) );
  AND2_X1 U476 ( .A1(n558), .A2(n557), .ZN(n437) );
  XNOR2_X1 U477 ( .A(n554), .B(KEYINPUT88), .ZN(n556) );
  AND2_X1 U478 ( .A1(G214), .A2(n519), .ZN(n370) );
  XOR2_X1 U479 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n371) );
  XOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT76), .Z(n372) );
  XOR2_X1 U481 ( .A(n679), .B(KEYINPUT80), .Z(n373) );
  XNOR2_X1 U482 ( .A(KEYINPUT3), .B(G119), .ZN(n518) );
  AND2_X1 U483 ( .A1(n661), .A2(n580), .ZN(n375) );
  NOR2_X1 U484 ( .A1(n578), .A2(n577), .ZN(n376) );
  XNOR2_X1 U485 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n377) );
  XOR2_X1 U486 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n378) );
  XNOR2_X1 U487 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n546) );
  NOR2_X1 U488 ( .A1(n659), .A2(n632), .ZN(n379) );
  NAND2_X1 U489 ( .A1(KEYINPUT2), .A2(KEYINPUT74), .ZN(n380) );
  XOR2_X1 U490 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n381) );
  INV_X1 U491 ( .A(n594), .ZN(n423) );
  XNOR2_X2 U492 ( .A(n634), .B(KEYINPUT65), .ZN(n382) );
  XNOR2_X1 U493 ( .A(n634), .B(KEYINPUT65), .ZN(n705) );
  NAND2_X2 U494 ( .A1(n633), .A2(n379), .ZN(n634) );
  NAND2_X1 U495 ( .A1(n425), .A2(n375), .ZN(n411) );
  XNOR2_X1 U496 ( .A(n503), .B(n426), .ZN(n425) );
  NAND2_X1 U497 ( .A1(n446), .A2(n447), .ZN(n383) );
  NAND2_X1 U498 ( .A1(n446), .A2(n447), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n573), .B(KEYINPUT75), .ZN(n614) );
  XNOR2_X2 U500 ( .A(n384), .B(n380), .ZN(n633) );
  NOR2_X2 U501 ( .A1(n724), .A2(n740), .ZN(n384) );
  XNOR2_X1 U502 ( .A(n621), .B(n620), .ZN(n385) );
  NAND2_X1 U503 ( .A1(n388), .A2(n400), .ZN(n387) );
  NAND2_X1 U504 ( .A1(n397), .A2(n390), .ZN(n389) );
  INV_X1 U505 ( .A(KEYINPUT35), .ZN(n390) );
  INV_X1 U506 ( .A(n398), .ZN(n391) );
  NAND2_X1 U507 ( .A1(n394), .A2(KEYINPUT35), .ZN(n393) );
  NAND2_X1 U508 ( .A1(n398), .A2(n397), .ZN(n394) );
  NAND2_X1 U509 ( .A1(n396), .A2(KEYINPUT35), .ZN(n395) );
  INV_X1 U510 ( .A(n400), .ZN(n396) );
  NAND2_X1 U511 ( .A1(n556), .A2(KEYINPUT34), .ZN(n397) );
  NAND2_X1 U512 ( .A1(n688), .A2(KEYINPUT34), .ZN(n399) );
  NAND2_X1 U513 ( .A1(n558), .A2(n401), .ZN(n400) );
  NOR2_X1 U514 ( .A1(n688), .A2(KEYINPUT34), .ZN(n401) );
  INV_X1 U515 ( .A(n612), .ZN(n442) );
  NAND2_X1 U516 ( .A1(n407), .A2(n403), .ZN(n402) );
  INV_X1 U517 ( .A(n554), .ZN(n405) );
  INV_X1 U518 ( .A(n670), .ZN(n406) );
  NAND2_X1 U519 ( .A1(n409), .A2(n439), .ZN(n408) );
  XNOR2_X1 U520 ( .A(n411), .B(n410), .ZN(n409) );
  INV_X1 U521 ( .A(KEYINPUT66), .ZN(n410) );
  INV_X1 U522 ( .A(n429), .ZN(n622) );
  XNOR2_X2 U523 ( .A(n412), .B(n377), .ZN(n429) );
  NAND2_X1 U524 ( .A1(n614), .A2(n676), .ZN(n412) );
  NAND2_X1 U525 ( .A1(n415), .A2(n413), .ZN(n570) );
  INV_X1 U526 ( .A(n660), .ZN(n413) );
  XNOR2_X2 U527 ( .A(n414), .B(n539), .ZN(n578) );
  INV_X1 U528 ( .A(n583), .ZN(n415) );
  XNOR2_X2 U529 ( .A(n418), .B(G131), .ZN(n506) );
  NAND2_X1 U530 ( .A1(n545), .A2(n419), .ZN(n433) );
  AND2_X1 U531 ( .A1(n625), .A2(n423), .ZN(n422) );
  AND2_X1 U532 ( .A1(n425), .A2(n424), .ZN(n562) );
  XNOR2_X1 U533 ( .A(n441), .B(n448), .ZN(n449) );
  NOR2_X2 U534 ( .A1(n600), .A2(n470), .ZN(n471) );
  NAND2_X1 U535 ( .A1(n633), .A2(n427), .ZN(n694) );
  NAND2_X1 U536 ( .A1(n574), .A2(n675), .ZN(n589) );
  NAND2_X1 U537 ( .A1(n640), .A2(n748), .ZN(n588) );
  XNOR2_X2 U538 ( .A(n528), .B(n527), .ZN(n580) );
  XNOR2_X2 U539 ( .A(G143), .B(G128), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n433), .A2(n546), .ZN(n436) );
  NAND2_X1 U541 ( .A1(n545), .A2(n435), .ZN(n434) );
  NAND2_X1 U542 ( .A1(n437), .A2(n655), .ZN(n645) );
  NAND2_X1 U543 ( .A1(n437), .A2(n653), .ZN(n644) );
  XNOR2_X2 U544 ( .A(n440), .B(n461), .ZN(n574) );
  NAND2_X1 U545 ( .A1(n700), .A2(n632), .ZN(n440) );
  XNOR2_X1 U546 ( .A(n459), .B(n720), .ZN(n700) );
  XNOR2_X1 U547 ( .A(n383), .B(G140), .ZN(n489) );
  AND2_X1 U548 ( .A1(G217), .A2(n537), .ZN(n443) );
  INV_X1 U549 ( .A(n544), .ZN(n554) );
  INV_X1 U550 ( .A(KEYINPUT45), .ZN(n564) );
  INV_X1 U551 ( .A(KEYINPUT19), .ZN(n463) );
  NAND2_X1 U552 ( .A1(n618), .A2(n617), .ZN(n621) );
  XNOR2_X1 U553 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U554 ( .A(n481), .B(n480), .ZN(n486) );
  NAND2_X1 U555 ( .A1(n444), .A2(G125), .ZN(n447) );
  NAND2_X1 U556 ( .A1(G146), .A2(n445), .ZN(n446) );
  XNOR2_X1 U557 ( .A(n449), .B(n512), .ZN(n453) );
  NAND2_X1 U558 ( .A1(G224), .A2(n741), .ZN(n450) );
  XNOR2_X1 U559 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U560 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U561 ( .A(KEYINPUT68), .B(G101), .ZN(n454) );
  XNOR2_X1 U562 ( .A(n455), .B(n507), .ZN(n459) );
  XNOR2_X1 U563 ( .A(KEYINPUT16), .B(n493), .ZN(n456) );
  XOR2_X1 U564 ( .A(G122), .B(n457), .Z(n481) );
  XNOR2_X1 U565 ( .A(KEYINPUT15), .B(G902), .ZN(n632) );
  INV_X1 U566 ( .A(G902), .ZN(n526) );
  INV_X1 U567 ( .A(G237), .ZN(n460) );
  NAND2_X1 U568 ( .A1(n526), .A2(n460), .ZN(n462) );
  AND2_X1 U569 ( .A1(n462), .A2(G210), .ZN(n461) );
  NAND2_X1 U570 ( .A1(n462), .A2(G214), .ZN(n675) );
  XNOR2_X1 U571 ( .A(n589), .B(n463), .ZN(n600) );
  NAND2_X1 U572 ( .A1(G234), .A2(G237), .ZN(n464) );
  XNOR2_X1 U573 ( .A(n464), .B(KEYINPUT14), .ZN(n466) );
  NAND2_X1 U574 ( .A1(n466), .A2(G952), .ZN(n465) );
  XNOR2_X1 U575 ( .A(n465), .B(KEYINPUT84), .ZN(n687) );
  NOR2_X1 U576 ( .A1(n687), .A2(G953), .ZN(n569) );
  NAND2_X1 U577 ( .A1(n466), .A2(G902), .ZN(n467) );
  XNOR2_X1 U578 ( .A(KEYINPUT86), .B(n467), .ZN(n566) );
  XNOR2_X1 U579 ( .A(KEYINPUT85), .B(G898), .ZN(n727) );
  NAND2_X1 U580 ( .A1(G953), .A2(n727), .ZN(n723) );
  NOR2_X1 U581 ( .A1(n566), .A2(n723), .ZN(n468) );
  XOR2_X1 U582 ( .A(KEYINPUT87), .B(n468), .Z(n469) );
  NOR2_X1 U583 ( .A1(n569), .A2(n469), .ZN(n470) );
  NAND2_X1 U584 ( .A1(n632), .A2(G234), .ZN(n473) );
  XNOR2_X1 U585 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n472) );
  XNOR2_X1 U586 ( .A(n473), .B(n472), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n537), .A2(G221), .ZN(n474) );
  XNOR2_X1 U588 ( .A(n474), .B(KEYINPUT21), .ZN(n475) );
  XNOR2_X1 U589 ( .A(n475), .B(KEYINPUT91), .ZN(n664) );
  INV_X1 U590 ( .A(n664), .ZN(n577) );
  XNOR2_X1 U591 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U592 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n478) );
  NAND2_X1 U593 ( .A1(G217), .A2(n532), .ZN(n484) );
  XNOR2_X1 U594 ( .A(n482), .B(KEYINPUT97), .ZN(n483) );
  XNOR2_X1 U595 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n486), .B(n485), .ZN(n712) );
  NOR2_X1 U597 ( .A1(n712), .A2(G902), .ZN(n487) );
  XNOR2_X1 U598 ( .A(G478), .B(n487), .ZN(n550) );
  XNOR2_X1 U599 ( .A(G143), .B(n506), .ZN(n488) );
  XNOR2_X1 U600 ( .A(n488), .B(G122), .ZN(n490) );
  XNOR2_X1 U601 ( .A(KEYINPUT11), .B(KEYINPUT94), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n371), .B(n491), .ZN(n492) );
  NOR2_X1 U603 ( .A1(G953), .A2(G237), .ZN(n519) );
  XNOR2_X1 U604 ( .A(n492), .B(n370), .ZN(n495) );
  XNOR2_X1 U605 ( .A(n493), .B(KEYINPUT95), .ZN(n494) );
  NOR2_X1 U606 ( .A1(G902), .A2(n636), .ZN(n499) );
  XNOR2_X1 U607 ( .A(KEYINPUT13), .B(G475), .ZN(n498) );
  XNOR2_X1 U608 ( .A(n499), .B(n498), .ZN(n551) );
  INV_X1 U609 ( .A(n551), .ZN(n500) );
  NAND2_X1 U610 ( .A1(n550), .A2(n500), .ZN(n575) );
  XNOR2_X1 U611 ( .A(n501), .B(KEYINPUT102), .ZN(n502) );
  NAND2_X1 U612 ( .A1(n544), .A2(n502), .ZN(n503) );
  XNOR2_X1 U613 ( .A(n504), .B(G134), .ZN(n505) );
  XNOR2_X1 U614 ( .A(n509), .B(n508), .ZN(n511) );
  NAND2_X1 U615 ( .A1(n741), .A2(G227), .ZN(n510) );
  XNOR2_X1 U616 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U617 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U618 ( .A(n525), .B(n514), .ZN(n708) );
  NAND2_X1 U619 ( .A1(n708), .A2(n526), .ZN(n516) );
  XNOR2_X1 U620 ( .A(KEYINPUT71), .B(G469), .ZN(n515) );
  XNOR2_X1 U621 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n518), .B(n517), .ZN(n523) );
  NAND2_X1 U623 ( .A1(G210), .A2(n519), .ZN(n520) );
  XNOR2_X1 U624 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U625 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U626 ( .A1(n641), .A2(n526), .ZN(n528) );
  XNOR2_X1 U627 ( .A(G472), .B(KEYINPUT93), .ZN(n527) );
  XNOR2_X1 U628 ( .A(n372), .B(n529), .ZN(n530) );
  XNOR2_X1 U629 ( .A(n531), .B(n530), .ZN(n534) );
  NAND2_X1 U630 ( .A1(G221), .A2(n532), .ZN(n533) );
  XNOR2_X1 U631 ( .A(n534), .B(n533), .ZN(n536) );
  INV_X1 U632 ( .A(n737), .ZN(n535) );
  XNOR2_X1 U633 ( .A(n536), .B(n535), .ZN(n715) );
  INV_X1 U634 ( .A(KEYINPUT25), .ZN(n538) );
  XNOR2_X1 U635 ( .A(KEYINPUT103), .B(n578), .ZN(n559) );
  INV_X1 U636 ( .A(n559), .ZN(n663) );
  NOR2_X1 U637 ( .A1(n661), .A2(n663), .ZN(n540) );
  AND2_X1 U638 ( .A1(n562), .A2(n540), .ZN(n541) );
  XNOR2_X1 U639 ( .A(n541), .B(KEYINPUT32), .ZN(n754) );
  INV_X1 U640 ( .A(KEYINPUT44), .ZN(n542) );
  INV_X1 U641 ( .A(n550), .ZN(n543) );
  NAND2_X1 U642 ( .A1(n543), .A2(n551), .ZN(n612) );
  NOR2_X1 U643 ( .A1(n661), .A2(n660), .ZN(n545) );
  NAND2_X1 U644 ( .A1(n547), .A2(n549), .ZN(n548) );
  INV_X1 U645 ( .A(KEYINPUT101), .ZN(n553) );
  OR2_X1 U646 ( .A1(n551), .A2(n550), .ZN(n623) );
  INV_X1 U647 ( .A(n623), .ZN(n655) );
  AND2_X1 U648 ( .A1(n551), .A2(n550), .ZN(n653) );
  NOR2_X1 U649 ( .A1(n655), .A2(n653), .ZN(n552) );
  XNOR2_X1 U650 ( .A(n553), .B(n552), .ZN(n679) );
  INV_X1 U651 ( .A(n661), .ZN(n560) );
  NOR2_X1 U652 ( .A1(n580), .A2(n660), .ZN(n555) );
  NAND2_X1 U653 ( .A1(n560), .A2(n555), .ZN(n670) );
  INV_X1 U654 ( .A(n556), .ZN(n558) );
  INV_X1 U655 ( .A(n580), .ZN(n666) );
  NOR2_X1 U656 ( .A1(n666), .A2(n570), .ZN(n557) );
  NOR2_X1 U657 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U658 ( .A1(n562), .A2(n561), .ZN(n643) );
  INV_X1 U659 ( .A(n675), .ZN(n565) );
  OR2_X1 U660 ( .A1(n566), .A2(n741), .ZN(n567) );
  NOR2_X1 U661 ( .A1(n567), .A2(G900), .ZN(n568) );
  OR2_X1 U662 ( .A1(n569), .A2(n568), .ZN(n579) );
  XNOR2_X1 U663 ( .A(n570), .B(KEYINPUT105), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n572), .A2(n571), .ZN(n573) );
  BUF_X1 U665 ( .A(n574), .Z(n611) );
  NAND2_X1 U666 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U667 ( .A1(n579), .A2(n376), .ZN(n590) );
  OR2_X1 U668 ( .A1(n580), .A2(n590), .ZN(n582) );
  XNOR2_X1 U669 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n581) );
  XNOR2_X1 U670 ( .A(n582), .B(n581), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n583), .B(KEYINPUT106), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n586), .B(KEYINPUT42), .ZN(n748) );
  XOR2_X1 U673 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n587) );
  XNOR2_X1 U674 ( .A(n588), .B(n587), .ZN(n618) );
  BUF_X1 U675 ( .A(n589), .Z(n594) );
  INV_X1 U676 ( .A(n653), .ZN(n593) );
  INV_X1 U677 ( .A(n590), .ZN(n591) );
  NOR2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n625) );
  XNOR2_X1 U679 ( .A(n595), .B(KEYINPUT108), .ZN(n756) );
  INV_X1 U680 ( .A(n679), .ZN(n607) );
  NOR2_X1 U681 ( .A1(KEYINPUT80), .A2(n607), .ZN(n599) );
  INV_X1 U682 ( .A(KEYINPUT47), .ZN(n596) );
  NAND2_X1 U683 ( .A1(KEYINPUT80), .A2(n596), .ZN(n597) );
  NOR2_X1 U684 ( .A1(n679), .A2(n597), .ZN(n598) );
  NOR2_X1 U685 ( .A1(n599), .A2(n598), .ZN(n606) );
  BUF_X1 U686 ( .A(n600), .Z(n602) );
  NOR2_X1 U687 ( .A1(n602), .A2(n601), .ZN(n604) );
  AND2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n651) );
  INV_X1 U689 ( .A(n651), .ZN(n605) );
  OR2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n651), .A2(n607), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n608), .A2(KEYINPUT47), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n615) );
  INV_X1 U694 ( .A(n611), .ZN(n628) );
  NOR2_X1 U695 ( .A1(n628), .A2(n612), .ZN(n613) );
  AND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n639) );
  OR2_X1 U697 ( .A1(n615), .A2(n639), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n756), .A2(n616), .ZN(n617) );
  XNOR2_X1 U699 ( .A(KEYINPUT81), .B(KEYINPUT48), .ZN(n619) );
  XNOR2_X1 U700 ( .A(n619), .B(KEYINPUT70), .ZN(n620) );
  NOR2_X1 U701 ( .A1(n622), .A2(n623), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n624), .B(KEYINPUT109), .ZN(n750) );
  INV_X1 U703 ( .A(n750), .ZN(n630) );
  AND2_X1 U704 ( .A1(n675), .A2(n625), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n661), .A2(n626), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n627), .B(KEYINPUT43), .ZN(n629) );
  AND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n658) );
  NOR2_X1 U708 ( .A1(n630), .A2(n658), .ZN(n631) );
  NOR2_X1 U709 ( .A1(KEYINPUT2), .A2(KEYINPUT74), .ZN(n659) );
  NAND2_X1 U710 ( .A1(n382), .A2(G475), .ZN(n637) );
  INV_X1 U711 ( .A(KEYINPUT59), .ZN(n635) );
  INV_X1 U712 ( .A(G952), .ZN(n638) );
  XOR2_X1 U713 ( .A(G143), .B(n639), .Z(G45) );
  XNOR2_X1 U714 ( .A(n640), .B(G131), .ZN(G33) );
  NAND2_X1 U715 ( .A1(n382), .A2(G472), .ZN(n642) );
  XOR2_X1 U716 ( .A(G101), .B(n643), .Z(G3) );
  XNOR2_X1 U717 ( .A(n644), .B(G104), .ZN(G6) );
  XOR2_X1 U718 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n646) );
  XNOR2_X1 U719 ( .A(n646), .B(n645), .ZN(n648) );
  XOR2_X1 U720 ( .A(G107), .B(KEYINPUT26), .Z(n647) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(G9) );
  XOR2_X1 U722 ( .A(G128), .B(KEYINPUT29), .Z(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n655), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(G30) );
  NAND2_X1 U725 ( .A1(n651), .A2(n653), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n652), .B(G146), .ZN(G48) );
  NAND2_X1 U727 ( .A1(n656), .A2(n653), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(G113), .ZN(G15) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(G116), .ZN(G18) );
  XOR2_X1 U731 ( .A(G140), .B(n658), .Z(G42) );
  XNOR2_X1 U732 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n699) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n662), .B(KEYINPUT50), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U736 ( .A(KEYINPUT49), .B(n665), .Z(n667) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U740 ( .A(KEYINPUT114), .B(n672), .ZN(n673) );
  XNOR2_X1 U741 ( .A(n673), .B(KEYINPUT51), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n689), .A2(n674), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n575), .A2(n677), .ZN(n681) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n682), .A2(n688), .ZN(n683) );
  NOR2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U749 ( .A(n685), .B(KEYINPUT52), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U752 ( .A(n690), .B(KEYINPUT115), .Z(n691) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  AND2_X1 U754 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U755 ( .A(KEYINPUT116), .B(n695), .ZN(n696) );
  NAND2_X1 U756 ( .A1(n696), .A2(n741), .ZN(n697) );
  XNOR2_X1 U757 ( .A(n697), .B(KEYINPUT53), .ZN(n698) );
  XNOR2_X1 U758 ( .A(n699), .B(n698), .ZN(G75) );
  BUF_X1 U759 ( .A(n700), .Z(n701) );
  XOR2_X1 U760 ( .A(KEYINPUT56), .B(KEYINPUT119), .Z(n703) );
  XNOR2_X1 U761 ( .A(n704), .B(n703), .ZN(G51) );
  NAND2_X1 U762 ( .A1(n714), .A2(G469), .ZN(n710) );
  XOR2_X1 U763 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n706) );
  XOR2_X1 U764 ( .A(n706), .B(KEYINPUT120), .Z(n707) );
  XNOR2_X1 U765 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U766 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U767 ( .A1(n719), .A2(n711), .ZN(G54) );
  NAND2_X1 U768 ( .A1(n714), .A2(G478), .ZN(n713) );
  NAND2_X1 U769 ( .A1(n714), .A2(G217), .ZN(n717) );
  XOR2_X1 U770 ( .A(n715), .B(KEYINPUT121), .Z(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(G66) );
  XNOR2_X1 U773 ( .A(G101), .B(n720), .ZN(n721) );
  XNOR2_X1 U774 ( .A(n721), .B(G110), .ZN(n722) );
  NAND2_X1 U775 ( .A1(n723), .A2(n722), .ZN(n734) );
  NOR2_X1 U776 ( .A1(G953), .A2(n724), .ZN(n731) );
  XOR2_X1 U777 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n726) );
  NAND2_X1 U778 ( .A1(G224), .A2(G953), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U781 ( .A(KEYINPUT123), .B(n729), .Z(n730) );
  NOR2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U783 ( .A(KEYINPUT125), .B(n732), .Z(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U785 ( .A(KEYINPUT124), .B(n735), .ZN(G69) );
  XNOR2_X1 U786 ( .A(n737), .B(n736), .ZN(n738) );
  XOR2_X1 U787 ( .A(n739), .B(n738), .Z(n743) );
  XNOR2_X1 U788 ( .A(n740), .B(n743), .ZN(n742) );
  NAND2_X1 U789 ( .A1(n742), .A2(n741), .ZN(n747) );
  XNOR2_X1 U790 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(G953), .ZN(n746) );
  NAND2_X1 U793 ( .A1(n747), .A2(n746), .ZN(G72) );
  XNOR2_X1 U794 ( .A(G137), .B(n748), .ZN(n749) );
  XNOR2_X1 U795 ( .A(n749), .B(KEYINPUT126), .ZN(G39) );
  XNOR2_X1 U796 ( .A(G134), .B(n750), .ZN(G36) );
  BUF_X1 U797 ( .A(n751), .Z(n752) );
  XOR2_X1 U798 ( .A(G110), .B(KEYINPUT112), .Z(n753) );
  XNOR2_X1 U799 ( .A(n752), .B(n753), .ZN(G12) );
  XOR2_X1 U800 ( .A(G122), .B(n549), .Z(G24) );
  XOR2_X1 U801 ( .A(G119), .B(n754), .Z(G21) );
  XOR2_X1 U802 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n755) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U804 ( .A(G125), .B(n757), .ZN(G27) );
endmodule

