//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  AOI21_X1  g001(.A(new_n202), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR3_X1   g004(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  OAI221_X1 g006(.A(new_n203), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(KEYINPUT15), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n209), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT17), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT95), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  INV_X1    g016(.A(G8gat), .ZN(new_n218));
  OAI221_X1 g017(.A(new_n217), .B1(KEYINPUT94), .B2(new_n218), .C1(G1gat), .C2(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT94), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n210), .A2(KEYINPUT93), .A3(new_n211), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT93), .B1(new_n210), .B2(new_n211), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n214), .A2(new_n222), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT96), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n230), .B(new_n221), .C1(new_n225), .C2(new_n226), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n226), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n224), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n230), .B1(new_n234), .B2(new_n221), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n228), .B(new_n229), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT97), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(KEYINPUT18), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n221), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT96), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n231), .ZN(new_n242));
  INV_X1    g041(.A(new_n238), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n242), .A2(new_n229), .A3(new_n228), .A4(new_n243), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n235), .A2(new_n232), .B1(new_n221), .B2(new_n234), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n229), .B(KEYINPUT13), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n239), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G197gat), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT11), .B(G169gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n252), .B(KEYINPUT12), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n244), .A3(new_n247), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT80), .ZN(new_n260));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT2), .ZN(new_n262));
  INV_X1    g061(.A(G141gat), .ZN(new_n263));
  INV_X1    g062(.A(G148gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G155gat), .B(G162gat), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n260), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G141gat), .B(G148gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(G155gat), .B2(G162gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n269), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n268), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(KEYINPUT80), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G134gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G127gat), .ZN(new_n282));
  INV_X1    g081(.A(G127gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G134gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G113gat), .B2(G120gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n285), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(KEYINPUT73), .A2(G113gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT73), .A2(G113gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT1), .B1(new_n286), .B2(new_n287), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n282), .A3(new_n284), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n291), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n272), .A2(new_n280), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n279), .ZN(new_n299));
  INV_X1    g098(.A(new_n296), .ZN(new_n300));
  INV_X1    g099(.A(new_n294), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n295), .B1(new_n286), .B2(new_n287), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n300), .A2(new_n301), .B1(new_n302), .B2(new_n285), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n259), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n272), .A2(new_n280), .A3(KEYINPUT3), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n303), .B1(new_n299), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT4), .A4(new_n299), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n304), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n312), .A2(new_n306), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n308), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G1gat), .B(G29gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT0), .ZN(new_n322));
  XNOR2_X1  g121(.A(G57gat), .B(G85gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n322), .B(new_n323), .Z(new_n324));
  NAND4_X1  g123(.A1(new_n313), .A2(new_n315), .A3(new_n317), .A4(new_n299), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n304), .A2(KEYINPUT4), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n327), .A2(new_n259), .A3(new_n306), .A4(new_n312), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n320), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT82), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n320), .A2(new_n328), .ZN(new_n332));
  INV_X1    g131(.A(new_n324), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT6), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n320), .A2(KEYINPUT82), .A3(new_n324), .A4(new_n328), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n331), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT83), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n334), .B2(new_n335), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n324), .B1(new_n320), .B2(new_n328), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G197gat), .B(G204gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344));
  INV_X1    g143(.A(G218gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346));
  INV_X1    g145(.A(G211gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n343), .B(new_n344), .C1(new_n350), .C2(KEYINPUT22), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n354));
  OAI21_X1  g153(.A(G218gat), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT22), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n344), .B1(new_n357), .B2(new_n343), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  AND2_X1   g159(.A1(KEYINPUT69), .A2(KEYINPUT24), .ZN(new_n361));
  NOR2_X1   g160(.A1(KEYINPUT69), .A2(KEYINPUT24), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(G190gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT70), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT70), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n369), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n363), .A2(new_n366), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n373), .A2(KEYINPUT25), .ZN(new_n374));
  NAND2_X1  g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT67), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT67), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(G169gat), .B2(G176gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(KEYINPUT23), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n382), .A3(KEYINPUT68), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT68), .B1(new_n377), .B2(new_n382), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n371), .B(new_n374), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT64), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n375), .B1(new_n378), .B2(KEYINPUT23), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n372), .A2(G169gat), .A3(G176gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n378), .A2(KEYINPUT23), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n391), .A2(new_n373), .A3(KEYINPUT64), .A4(new_n375), .ZN(new_n392));
  INV_X1    g191(.A(new_n360), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n366), .B(new_n367), .C1(new_n393), .C2(KEYINPUT24), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n395), .A2(KEYINPUT65), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT65), .B1(new_n395), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n386), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT26), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n379), .A2(new_n400), .A3(new_n381), .ZN(new_n401));
  INV_X1    g200(.A(new_n375), .ZN(new_n402));
  INV_X1    g201(.A(new_n378), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(KEYINPUT26), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n393), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT71), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n408), .A2(new_n364), .A3(KEYINPUT27), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n409), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT27), .B1(new_n408), .B2(new_n364), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT27), .B(G183gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n365), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n410), .A2(new_n411), .B1(new_n413), .B2(KEYINPUT28), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n406), .A2(new_n407), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n399), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n399), .A2(new_n415), .B1(new_n418), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n359), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n418), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n371), .A2(new_n374), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT68), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n379), .A2(KEYINPUT23), .A3(new_n381), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n375), .B(KEYINPUT66), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n422), .B1(new_n383), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n395), .A2(new_n396), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT65), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n395), .A2(KEYINPUT65), .A3(new_n396), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n406), .A2(new_n407), .A3(new_n414), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n421), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n359), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n399), .A2(new_n415), .A3(new_n416), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G8gat), .B(G36gat), .Z(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT78), .ZN(new_n439));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n420), .A2(new_n437), .A3(KEYINPUT30), .A4(new_n441), .ZN(new_n445));
  INV_X1    g244(.A(new_n441), .ZN(new_n446));
  INV_X1    g245(.A(new_n437), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n435), .B1(new_n434), .B2(new_n436), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n444), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n342), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n310), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n278), .B2(new_n279), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n359), .B1(new_n456), .B2(KEYINPUT29), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n457), .B2(KEYINPUT86), .ZN(new_n458));
  INV_X1    g257(.A(new_n299), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n343), .B1(new_n350), .B2(KEYINPUT22), .ZN(new_n460));
  INV_X1    g259(.A(new_n344), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT29), .B1(new_n462), .B2(new_n351), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n459), .B1(new_n463), .B2(new_n455), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT85), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n359), .B(new_n466), .C1(new_n456), .C2(KEYINPUT29), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n468), .B(new_n459), .C1(new_n463), .C2(new_n455), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n458), .A2(new_n465), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n272), .A2(new_n280), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n457), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n454), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n470), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n470), .B2(new_n474), .ZN(new_n478));
  XOR2_X1   g277(.A(G78gat), .B(G106gat), .Z(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(G50gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(G22gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n477), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n469), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n457), .A2(KEYINPUT86), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n453), .A3(new_n467), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n474), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n475), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n474), .A3(new_n476), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n452), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n444), .A2(new_n445), .A3(new_n449), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n306), .B1(new_n327), .B2(new_n312), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT39), .B1(new_n305), .B2(new_n307), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT39), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n333), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(KEYINPUT40), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT40), .B1(new_n496), .B2(new_n498), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(new_n340), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n493), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n337), .A2(new_n339), .A3(new_n341), .A4(new_n442), .ZN(new_n503));
  XOR2_X1   g302(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n504));
  NAND3_X1  g303(.A1(new_n420), .A2(new_n437), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n441), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n448), .B1(new_n510), .B2(new_n437), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n510), .B2(new_n437), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT38), .B1(new_n512), .B2(KEYINPUT37), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n503), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT37), .B1(new_n447), .B2(new_n448), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n508), .A2(new_n507), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT38), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n502), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n492), .B1(new_n518), .B2(new_n491), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n313), .A2(new_n315), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n432), .B2(new_n433), .ZN(new_n521));
  NAND2_X1  g320(.A1(G227gat), .A2(G233gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n520), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n399), .A2(new_n523), .A3(new_n415), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n522), .B2(KEYINPUT76), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n525), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT32), .ZN(new_n529));
  INV_X1    g328(.A(new_n522), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n399), .A2(new_n523), .A3(new_n415), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n523), .B1(new_n399), .B2(new_n415), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT75), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n521), .A2(new_n524), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT75), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n530), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n529), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G43gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(G71gat), .B(G99gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT33), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n528), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n536), .B1(new_n535), .B2(new_n530), .ZN(new_n546));
  AOI211_X1 g345(.A(KEYINPUT75), .B(new_n522), .C1(new_n521), .C2(new_n524), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT32), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  INV_X1    g348(.A(new_n541), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n528), .ZN(new_n553));
  OAI211_X1 g352(.A(KEYINPUT32), .B(new_n544), .C1(new_n546), .C2(new_n547), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT36), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n545), .A2(new_n551), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n537), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n541), .B1(new_n559), .B2(KEYINPUT32), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n560), .A2(new_n548), .B1(new_n538), .B2(new_n544), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n557), .B(new_n558), .C1(new_n561), .C2(new_n553), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n519), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n483), .A2(new_n490), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n553), .A2(new_n554), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n568), .A2(new_n555), .A3(new_n451), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n555), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n491), .B1(new_n551), .B2(new_n545), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n452), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(KEYINPUT91), .A3(KEYINPUT35), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n568), .A2(new_n555), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n451), .A2(KEYINPUT90), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n342), .A2(new_n450), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n576), .A2(new_n570), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n571), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n258), .B1(new_n563), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G120gat), .B(G148gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT103), .ZN(new_n584));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT7), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n588), .B2(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G99gat), .B(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n593), .A2(new_n597), .A3(new_n595), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT9), .ZN(new_n607));
  XNOR2_X1  g406(.A(G57gat), .B(G64gat), .ZN(new_n608));
  OAI221_X1 g407(.A(new_n605), .B1(new_n603), .B2(new_n604), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(G57gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT99), .A2(G57gat), .A3(G64gat), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n602), .A2(KEYINPUT9), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n606), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n599), .A2(new_n609), .A3(new_n616), .A4(new_n600), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT102), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n601), .A2(new_n621), .A3(new_n617), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT10), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n587), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n587), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n620), .A2(new_n627), .A3(new_n622), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n586), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n626), .A2(new_n628), .A3(new_n586), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n630), .A2(KEYINPUT104), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT104), .B1(new_n630), .B2(new_n631), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  XNOR2_X1  g437(.A(G127gat), .B(G155gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT100), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G183gat), .B(G211gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n643), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n222), .B1(new_n635), .B2(new_n617), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n644), .B2(new_n645), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n214), .A2(new_n227), .A3(new_n601), .ZN(new_n652));
  XOR2_X1   g451(.A(G190gat), .B(G218gat), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n601), .ZN(new_n655));
  AND2_X1   g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n234), .A2(new_n655), .B1(KEYINPUT41), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n652), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n654), .B1(new_n652), .B2(new_n657), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n656), .A2(KEYINPUT41), .ZN(new_n660));
  XNOR2_X1  g459(.A(G134gat), .B(G162gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OR3_X1    g462(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(new_n658), .B2(new_n659), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n634), .A2(new_n651), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n582), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n342), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n493), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n674), .A2(KEYINPUT105), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n674), .A2(new_n677), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(KEYINPUT42), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n218), .B1(new_n670), .B2(new_n493), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n682), .A2(new_n675), .B1(new_n674), .B2(new_n677), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n678), .B1(new_n681), .B2(new_n683), .ZN(G1325gat));
  NAND2_X1  g483(.A1(new_n556), .A2(new_n562), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n556), .A2(new_n562), .A3(KEYINPUT106), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G15gat), .B1(new_n669), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n552), .A2(new_n555), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(new_n669), .B2(new_n694), .ZN(G1326gat));
  NOR2_X1   g494(.A1(new_n669), .A2(new_n565), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n651), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n634), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n666), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n582), .A2(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(G29gat), .A3(new_n342), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT45), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n563), .A2(new_n581), .ZN(new_n705));
  INV_X1    g504(.A(new_n666), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n706), .A2(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n700), .A2(new_n258), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n519), .A2(new_n687), .A3(new_n688), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n666), .B1(new_n710), .B2(new_n581), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n708), .B(new_n709), .C1(KEYINPUT44), .C2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(KEYINPUT107), .A3(new_n342), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT107), .B1(new_n712), .B2(new_n342), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G29gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n704), .B1(new_n713), .B2(new_n715), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n702), .A2(G36gat), .A3(new_n450), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n712), .B2(new_n450), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n702), .B2(new_n693), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n689), .A2(G43gat), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n722), .B(new_n723), .C1(new_n712), .C2(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n725), .A2(KEYINPUT109), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n722), .B1(new_n712), .B2(new_n724), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT47), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(KEYINPUT109), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n712), .B2(new_n565), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT48), .B1(new_n731), .B2(KEYINPUT111), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n565), .A2(G50gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT110), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n731), .B1(new_n702), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  OAI221_X1 g536(.A(new_n731), .B1(KEYINPUT111), .B2(KEYINPUT48), .C1(new_n702), .C2(new_n735), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1331gat));
  NAND2_X1  g538(.A1(new_n710), .A2(new_n581), .ZN(new_n740));
  NOR4_X1   g539(.A1(new_n699), .A2(new_n634), .A3(new_n257), .A4(new_n706), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n342), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n612), .ZN(G1332gat));
  AND2_X1   g543(.A1(new_n740), .A2(new_n741), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n450), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT112), .ZN(new_n748));
  OR2_X1    g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1333gat));
  OR3_X1    g549(.A1(new_n742), .A2(G71gat), .A3(new_n693), .ZN(new_n751));
  OAI21_X1  g550(.A(G71gat), .B1(new_n742), .B2(new_n690), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g553(.A1(new_n745), .A2(new_n491), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n634), .A2(G85gat), .A3(new_n342), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n257), .A2(new_n651), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT113), .ZN(new_n759));
  AND4_X1   g558(.A1(KEYINPUT51), .A2(new_n740), .A3(new_n706), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT51), .B1(new_n711), .B2(new_n759), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n760), .A2(new_n761), .A3(KEYINPUT114), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n740), .A2(new_n706), .A3(new_n759), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n759), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n757), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n634), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n759), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n708), .B(new_n771), .C1(KEYINPUT44), .C2(new_n711), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n342), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n772), .B2(new_n450), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n634), .A2(G92gat), .A3(new_n450), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n760), .B2(new_n761), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT52), .ZN(G1337gat));
  NOR3_X1   g578(.A1(new_n693), .A2(G99gat), .A3(new_n634), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n762), .B2(new_n768), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782));
  OAI21_X1  g581(.A(G99gat), .B1(new_n772), .B2(new_n690), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n780), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT114), .B1(new_n760), .B2(new_n761), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n763), .A3(new_n767), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n783), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT115), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n784), .A2(new_n790), .ZN(G1338gat));
  OAI21_X1  g590(.A(G106gat), .B1(new_n772), .B2(new_n565), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n634), .A2(G106gat), .A3(new_n565), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT116), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n760), .B2(new_n761), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g596(.A1(new_n667), .A2(new_n257), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n620), .A2(new_n622), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n624), .ZN(new_n801));
  INV_X1    g600(.A(new_n625), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n627), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n626), .A3(KEYINPUT54), .ZN(new_n804));
  INV_X1    g603(.A(new_n586), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n806), .B(new_n587), .C1(new_n623), .C2(new_n625), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n631), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n803), .A2(new_n626), .A3(KEYINPUT54), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n805), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n257), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n229), .B1(new_n242), .B2(new_n228), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n245), .A2(new_n246), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n252), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n256), .B(new_n817), .C1(new_n632), .C2(new_n633), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n666), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n813), .A2(new_n631), .A3(new_n808), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n256), .A2(new_n817), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n699), .B1(new_n823), .B2(new_n666), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n799), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n826), .A3(new_n565), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n821), .A2(new_n822), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n651), .B1(new_n828), .B2(new_n706), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n798), .B1(new_n829), .B2(new_n819), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT117), .B1(new_n830), .B2(new_n491), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n342), .A2(new_n493), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n827), .A2(new_n831), .A3(new_n692), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n258), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n825), .A2(new_n671), .A3(new_n576), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT118), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n493), .B1(new_n835), .B2(KEYINPUT118), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT119), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n257), .A2(new_n292), .A3(new_n293), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n834), .B1(new_n839), .B2(new_n840), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n833), .B2(new_n634), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n770), .A2(new_n287), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n839), .B2(new_n843), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n833), .B2(new_n699), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n651), .A2(new_n283), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n838), .B2(new_n846), .ZN(G1342gat));
  NAND2_X1  g646(.A1(new_n706), .A2(new_n281), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n838), .A2(KEYINPUT56), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n833), .B2(new_n666), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT56), .B1(new_n838), .B2(new_n848), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G1343gat));
  OR3_X1    g651(.A1(new_n830), .A2(KEYINPUT57), .A3(new_n565), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT57), .B1(new_n830), .B2(new_n565), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n690), .A3(new_n832), .A4(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G141gat), .B1(new_n855), .B2(new_n258), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n830), .A2(new_n342), .A3(new_n493), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n689), .A2(new_n565), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n263), .A3(new_n257), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g662(.A1(new_n860), .A2(new_n264), .A3(new_n770), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  INV_X1    g664(.A(new_n855), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n770), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(G148gat), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n865), .B(G148gat), .C1(new_n855), .C2(new_n634), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n864), .B1(new_n868), .B2(new_n870), .ZN(G1345gat));
  AOI21_X1  g670(.A(G155gat), .B1(new_n860), .B2(new_n651), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n651), .A2(G155gat), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT120), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n866), .B2(new_n874), .ZN(G1346gat));
  OR3_X1    g674(.A1(new_n859), .A2(G162gat), .A3(new_n666), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(KEYINPUT121), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(KEYINPUT121), .ZN(new_n878));
  OAI21_X1  g677(.A(G162gat), .B1(new_n855), .B2(new_n666), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(G1347gat));
  NOR2_X1   g679(.A1(new_n671), .A2(new_n450), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n827), .A2(new_n831), .A3(new_n692), .A4(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(G169gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n882), .A2(new_n883), .A3(new_n258), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n825), .B2(new_n342), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n830), .A2(KEYINPUT122), .A3(new_n671), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n568), .A2(new_n555), .A3(new_n450), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n257), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n884), .B1(new_n891), .B2(new_n883), .ZN(G1348gat));
  INV_X1    g691(.A(G176gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n893), .A3(new_n770), .ZN(new_n894));
  OAI21_X1  g693(.A(G176gat), .B1(new_n882), .B2(new_n634), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1349gat));
  OAI21_X1  g695(.A(G183gat), .B1(new_n882), .B2(new_n699), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n651), .A2(new_n412), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n889), .B(new_n899), .C1(new_n886), .C2(new_n887), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT123), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT60), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n365), .A3(new_n706), .ZN(new_n909));
  OAI21_X1  g708(.A(G190gat), .B1(new_n882), .B2(new_n666), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(G1351gat));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n853), .A2(new_n690), .A3(new_n854), .A4(new_n881), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n258), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G197gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n916), .A2(new_n915), .A3(new_n258), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n689), .A2(new_n565), .A3(new_n450), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n888), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n258), .A2(G197gat), .ZN(new_n924));
  OAI22_X1  g723(.A1(new_n918), .A2(new_n919), .B1(new_n923), .B2(new_n924), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n634), .A2(G204gat), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n888), .A2(new_n921), .A3(new_n922), .A4(new_n926), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n916), .A2(KEYINPUT127), .A3(new_n634), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT127), .B1(new_n916), .B2(new_n634), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G204gat), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n928), .B(new_n929), .C1(new_n930), .C2(new_n932), .ZN(G1353gat));
  OR2_X1    g732(.A1(new_n916), .A2(new_n699), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT63), .B1(new_n934), .B2(G211gat), .ZN(new_n935));
  OAI211_X1 g734(.A(KEYINPUT63), .B(G211gat), .C1(new_n916), .C2(new_n699), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n651), .A2(new_n348), .A3(new_n349), .ZN(new_n938));
  OAI22_X1  g737(.A1(new_n935), .A2(new_n937), .B1(new_n923), .B2(new_n938), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n916), .B2(new_n666), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n706), .A2(new_n345), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n923), .B2(new_n941), .ZN(G1355gat));
endmodule


