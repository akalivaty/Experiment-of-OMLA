//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  XNOR2_X1  g001(.A(G183gat), .B(G211gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G15gat), .ZN(new_n206));
  INV_X1    g005(.A(G22gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G15gat), .A2(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G1gat), .ZN(new_n212));
  INV_X1    g011(.A(G1gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n213), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(G8gat), .B1(new_n214), .B2(KEYINPUT89), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT93), .ZN(new_n218));
  INV_X1    g017(.A(G57gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n219), .A2(KEYINPUT92), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(KEYINPUT92), .ZN(new_n221));
  OAI21_X1  g020(.A(G64gat), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G64gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G57gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G71gat), .A2(G78gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT9), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n222), .A2(new_n224), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n226), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n225), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n219), .A2(G64gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n230), .B1(new_n232), .B2(KEYINPUT9), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n218), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT92), .B(G57gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n224), .B1(new_n235), .B2(new_n223), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n225), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n232), .A2(KEYINPUT9), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n225), .A3(new_n229), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT93), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT21), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n217), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G127gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n242), .B2(new_n243), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(new_n247), .A3(new_n244), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n205), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT94), .B(G155gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G231gat), .A2(G233gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  NAND3_X1  g056(.A1(new_n250), .A2(new_n252), .A3(new_n205), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n254), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G190gat), .B(G218gat), .Z(new_n262));
  INV_X1    g061(.A(KEYINPUT96), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G85gat), .A2(G92gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT7), .ZN(new_n266));
  XNOR2_X1  g065(.A(G99gat), .B(G106gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G99gat), .A2(G106gat), .ZN(new_n268));
  INV_X1    g067(.A(G85gat), .ZN(new_n269));
  INV_X1    g068(.A(G92gat), .ZN(new_n270));
  AOI22_X1  g069(.A1(KEYINPUT8), .A2(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n266), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n267), .B1(new_n266), .B2(new_n271), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT17), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT14), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n276), .A2(G29gat), .A3(G36gat), .ZN(new_n277));
  OR2_X1    g076(.A1(G29gat), .A2(G36gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G29gat), .A2(G36gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT14), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G43gat), .B(G50gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT15), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT15), .ZN(new_n284));
  INV_X1    g083(.A(G43gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(G50gat), .ZN(new_n286));
  INV_X1    g085(.A(G50gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(G43gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n281), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n280), .A2(new_n278), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT15), .B(new_n282), .C1(new_n291), .C2(new_n277), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT88), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT88), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n275), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n290), .B2(new_n292), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n283), .A2(new_n289), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT88), .B1(new_n299), .B2(new_n281), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT17), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n274), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT95), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n262), .A2(new_n263), .ZN(new_n304));
  AND3_X1   g103(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n294), .A2(new_n296), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n272), .A2(new_n273), .ZN(new_n307));
  AOI211_X1 g106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n294), .A2(new_n275), .A3(new_n296), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT17), .B1(new_n298), .B2(new_n300), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT95), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n274), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n303), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G134gat), .B(G162gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n315), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n319), .A3(new_n308), .A4(new_n313), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n316), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n318), .B1(new_n316), .B2(new_n320), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n264), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n312), .B1(new_n311), .B2(new_n274), .ZN(new_n324));
  AOI211_X1 g123(.A(KEYINPUT95), .B(new_n307), .C1(new_n309), .C2(new_n310), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n319), .B1(new_n326), .B2(new_n308), .ZN(new_n327));
  INV_X1    g126(.A(new_n320), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n317), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n264), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n316), .A2(new_n318), .A3(new_n320), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n261), .B1(new_n323), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G141gat), .B(G148gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(KEYINPUT2), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT74), .B(G162gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(G155gat), .ZN(new_n343));
  INV_X1    g142(.A(G141gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(G148gat), .ZN(new_n345));
  INV_X1    g144(.A(G148gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(G141gat), .ZN(new_n347));
  OAI22_X1  g146(.A1(new_n345), .A2(new_n347), .B1(new_n336), .B2(new_n337), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n340), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT75), .B1(new_n349), .B2(KEYINPUT3), .ZN(new_n350));
  INV_X1    g149(.A(G162gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT74), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G162gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n354), .A3(G155gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT2), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n346), .A2(G141gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(G148gat), .ZN(new_n358));
  INV_X1    g157(.A(G155gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n351), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n357), .A2(new_n358), .B1(new_n360), .B2(new_n335), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n341), .B1(new_n345), .B2(new_n347), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n356), .A2(new_n361), .B1(new_n362), .B2(new_n338), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n350), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G197gat), .B(G204gat), .ZN(new_n368));
  INV_X1    g167(.A(G211gat), .ZN(new_n369));
  INV_X1    g168(.A(G218gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(KEYINPUT22), .B2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G211gat), .B(G218gat), .Z(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n375), .A2(KEYINPUT82), .ZN(new_n376));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n377), .B(KEYINPUT31), .Z(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n376), .A2(G228gat), .A3(G233gat), .A4(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(G228gat), .B(G233gat), .C1(new_n375), .C2(KEYINPUT82), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n374), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n365), .B1(new_n384), .B2(KEYINPUT29), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n349), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n367), .B2(new_n374), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G22gat), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n386), .B(new_n207), .C1(new_n367), .C2(new_n374), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n388), .A2(new_n287), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n287), .B1(new_n388), .B2(new_n389), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n383), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n389), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G50gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n388), .A2(new_n287), .A3(new_n389), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n394), .A2(new_n395), .B1(new_n380), .B2(new_n382), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399));
  OR3_X1    g198(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT67), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT67), .B1(new_n398), .B2(new_n399), .ZN(new_n401));
  INV_X1    g200(.A(new_n399), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n400), .B(new_n401), .C1(KEYINPUT26), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT66), .ZN(new_n404));
  OR2_X1    g203(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n404), .B(KEYINPUT28), .C1(new_n408), .C2(G190gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT28), .ZN(new_n411));
  AOI21_X1  g210(.A(G190gat), .B1(new_n405), .B2(new_n406), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(KEYINPUT66), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n403), .A2(new_n409), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G169gat), .ZN(new_n415));
  INV_X1    g214(.A(G176gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT65), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT65), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT23), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n417), .B1(new_n422), .B2(new_n402), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n399), .A2(KEYINPUT23), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n410), .A2(KEYINPUT24), .ZN(new_n425));
  OR2_X1    g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(KEYINPUT24), .A3(new_n410), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(new_n424), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n423), .A2(KEYINPUT64), .A3(new_n425), .A4(new_n427), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT25), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n430), .B2(new_n429), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n414), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G120gat), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT70), .B1(new_n434), .B2(G113gat), .ZN(new_n435));
  INV_X1    g234(.A(G113gat), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT69), .B1(new_n436), .B2(G120gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n436), .A3(G120gat), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT69), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(new_n434), .A3(G113gat), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n435), .A2(new_n437), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT1), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT1), .ZN(new_n446));
  INV_X1    g245(.A(G134gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n246), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G127gat), .A2(G134gat), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n444), .A2(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n442), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(KEYINPUT68), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G134gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n454), .A3(G127gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G113gat), .B(G120gat), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n455), .B(new_n448), .C1(KEYINPUT1), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n433), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G227gat), .ZN(new_n461));
  INV_X1    g260(.A(G233gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n458), .B(new_n414), .C1(new_n431), .C2(new_n432), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G43gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(G71gat), .ZN(new_n470));
  INV_X1    g269(.A(G99gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n465), .B(KEYINPUT32), .C1(new_n467), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(KEYINPUT72), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n480));
  INV_X1    g279(.A(new_n463), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n480), .A2(new_n481), .B1(KEYINPUT72), .B2(new_n477), .ZN(new_n482));
  INV_X1    g281(.A(new_n478), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n473), .A2(new_n483), .A3(new_n475), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n482), .ZN(new_n486));
  INV_X1    g285(.A(new_n484), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n473), .B2(new_n475), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT35), .B(new_n397), .C1(new_n485), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G8gat), .B(G36gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(new_n223), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(new_n270), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT29), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n433), .A2(new_n494), .B1(G226gat), .B2(G233gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n414), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(new_n424), .C1(KEYINPUT64), .C2(KEYINPUT25), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(G226gat), .A2(G233gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n495), .A2(new_n502), .A3(new_n384), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n500), .B2(KEYINPUT29), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n433), .A2(G226gat), .A3(G233gat), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n374), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n493), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n384), .B1(new_n495), .B2(new_n502), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n374), .A3(new_n505), .ZN(new_n509));
  INV_X1    g308(.A(new_n493), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(KEYINPUT30), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n508), .A2(new_n509), .A3(new_n513), .A4(new_n510), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n350), .A2(new_n366), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n458), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n458), .B2(new_n349), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT77), .B1(new_n458), .B2(new_n349), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT77), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n363), .A2(new_n522), .A3(new_n457), .A4(new_n451), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(KEYINPUT4), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n518), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G225gat), .A2(G233gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OR3_X1    g326(.A1(new_n525), .A2(KEYINPUT5), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n521), .A2(new_n519), .A3(new_n523), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT4), .B1(new_n458), .B2(new_n349), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT76), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT76), .B(KEYINPUT4), .C1(new_n458), .C2(new_n349), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n526), .A3(new_n518), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT5), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n523), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n458), .A2(new_n349), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n536), .B1(new_n539), .B2(new_n527), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n535), .A2(KEYINPUT78), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT78), .B1(new_n535), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n528), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G57gat), .B(G85gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G1gat), .B(G29gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n546), .B(new_n547), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT6), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n540), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT78), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n535), .A2(KEYINPUT78), .A3(new_n540), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT80), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n548), .A4(new_n528), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n548), .B(new_n528), .C1(new_n541), .C2(new_n542), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT80), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n550), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n548), .B1(new_n555), .B2(new_n528), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT6), .ZN(new_n562));
  AOI211_X1 g361(.A(KEYINPUT85), .B(new_n515), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT85), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n562), .ZN(new_n565));
  INV_X1    g364(.A(new_n515), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n490), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n562), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT81), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n560), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n550), .A2(new_n559), .A3(new_n557), .A4(KEYINPUT81), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n392), .A2(new_n396), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n487), .A2(new_n488), .A3(new_n486), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n482), .B1(new_n479), .B2(new_n484), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n573), .A2(new_n515), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n568), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n397), .B1(new_n573), .B2(new_n515), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n489), .A2(new_n485), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n489), .A2(new_n485), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n539), .A2(new_n527), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT39), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n590), .A2(KEYINPUT83), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n525), .A2(new_n527), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT83), .B1(new_n590), .B2(new_n591), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n593), .A2(KEYINPUT39), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n595), .A2(new_n549), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT40), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n561), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n598), .B(new_n515), .C1(new_n600), .C2(new_n597), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n503), .B2(new_n506), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT37), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n510), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n560), .B(new_n562), .C1(new_n602), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n511), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n601), .B(new_n574), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n581), .A2(new_n589), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n334), .B1(new_n580), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n416), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(G204gat), .Z(new_n615));
  AOI21_X1  g414(.A(new_n307), .B1(new_n234), .B2(new_n241), .ZN(new_n616));
  NOR4_X1   g415(.A1(new_n272), .A2(new_n228), .A3(new_n273), .A4(new_n233), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT10), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n242), .A2(new_n619), .A3(new_n274), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT100), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n622), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n616), .B2(new_n617), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n615), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT101), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n228), .A2(new_n218), .A3(new_n233), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT93), .B1(new_n238), .B2(new_n240), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n274), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n307), .A2(new_n238), .A3(new_n240), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n619), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n632), .A2(new_n633), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(KEYINPUT10), .A3(new_n307), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT97), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT97), .B1(new_n636), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n622), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT98), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n618), .B2(new_n620), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT97), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n647), .A3(new_n622), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n629), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n615), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n298), .A2(new_n300), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT90), .B1(new_n653), .B2(new_n217), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n215), .B(new_n216), .Z(new_n655));
  INV_X1    g454(.A(KEYINPUT90), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n306), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT91), .B1(new_n653), .B2(new_n217), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n653), .A2(KEYINPUT91), .A3(new_n217), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G229gat), .A2(G233gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT13), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n311), .A2(new_n217), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n653), .A2(new_n217), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT18), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n666), .B1(new_n311), .B2(new_n217), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(KEYINPUT18), .A3(new_n662), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n664), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT87), .ZN(new_n674));
  XNOR2_X1  g473(.A(G113gat), .B(G141gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G197gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT11), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n415), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  AND3_X1   g479(.A1(new_n673), .A2(new_n674), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n673), .B2(new_n674), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n652), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n612), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n573), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n213), .ZN(G1324gat));
  INV_X1    g487(.A(new_n685), .ZN(new_n689));
  INV_X1    g488(.A(G8gat), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n689), .B(new_n515), .C1(new_n211), .C2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n689), .B2(new_n515), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT42), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n691), .B2(new_n692), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1325gat));
  NOR3_X1   g497(.A1(new_n685), .A2(new_n206), .A3(new_n589), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n689), .A2(new_n582), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n206), .B2(new_n700), .ZN(G1326gat));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n574), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT43), .B(G22gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  NAND2_X1  g503(.A1(new_n580), .A2(new_n611), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n321), .A2(new_n322), .A3(new_n264), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n330), .B1(new_n329), .B2(new_n331), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n708), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n580), .B2(new_n611), .ZN(new_n712));
  INV_X1    g511(.A(new_n709), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n710), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n684), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n261), .B(KEYINPUT103), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(new_n573), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G29gat), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n712), .A2(new_n573), .A3(new_n684), .A4(new_n261), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n722), .A2(KEYINPUT102), .A3(G29gat), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT102), .B1(new_n722), .B2(G29gat), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n723), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(G1328gat));
  AOI211_X1 g527(.A(new_n717), .B(new_n711), .C1(new_n580), .C2(new_n611), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n261), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(G36gat), .A3(new_n566), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n515), .A3(new_n719), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G36gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1329gat));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  AOI21_X1  g535(.A(G43gat), .B1(new_n489), .B2(new_n485), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n712), .A2(new_n684), .A3(new_n261), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT47), .ZN(new_n739));
  INV_X1    g538(.A(new_n589), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n715), .B1(new_n705), .B2(new_n708), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n711), .B(new_n713), .C1(new_n580), .C2(new_n611), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n740), .B(new_n719), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n736), .B(new_n739), .C1(new_n743), .C2(G43gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(G43gat), .ZN(new_n745));
  INV_X1    g544(.A(new_n739), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT106), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n738), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n729), .A2(KEYINPUT105), .A3(new_n261), .A4(new_n737), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(G43gat), .B2(new_n743), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n744), .A2(new_n747), .B1(new_n752), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g552(.A1(new_n716), .A2(G50gat), .A3(new_n397), .A4(new_n719), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n287), .B1(new_n730), .B2(new_n574), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g556(.A1(new_n259), .A2(new_n260), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n683), .B(new_n758), .C1(new_n706), .C2(new_n707), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n580), .B2(new_n611), .ZN(new_n760));
  INV_X1    g559(.A(new_n652), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n686), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n235), .B(KEYINPUT107), .Z(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1332gat));
  NOR2_X1   g564(.A1(new_n761), .A2(new_n566), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  NAND4_X1  g569(.A1(new_n760), .A2(G71gat), .A3(new_n652), .A4(new_n740), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n760), .A2(new_n652), .A3(new_n582), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(G71gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g573(.A1(new_n760), .A2(new_n652), .A3(new_n397), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT108), .B(G78gat), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1335gat));
  INV_X1    g576(.A(new_n680), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n664), .A2(new_n670), .A3(new_n672), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(KEYINPUT87), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n673), .A2(new_n674), .A3(new_n680), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n758), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n712), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n708), .A4(new_n783), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n712), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n783), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n762), .A2(new_n269), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT110), .Z(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n783), .ZN(new_n795));
  INV_X1    g594(.A(new_n741), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n710), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n762), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n799), .B2(new_n269), .ZN(G1336gat));
  NAND2_X1  g599(.A1(new_n766), .A2(new_n270), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n791), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n652), .B(new_n783), .C1(new_n741), .C2(new_n742), .ZN(new_n804));
  OAI21_X1  g603(.A(G92gat), .B1(new_n804), .B2(new_n566), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT112), .B1(new_n712), .B2(new_n783), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(new_n785), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n801), .B(KEYINPUT111), .Z(new_n810));
  NAND4_X1  g609(.A1(new_n716), .A2(new_n652), .A3(new_n515), .A4(new_n783), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(G92gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n812), .B2(new_n806), .ZN(G1337gat));
  NAND4_X1  g612(.A1(new_n797), .A2(KEYINPUT113), .A3(new_n652), .A4(new_n740), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n804), .B2(new_n589), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n816), .A3(G99gat), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n791), .A2(new_n471), .A3(new_n652), .A4(new_n582), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1338gat));
  NOR3_X1   g618(.A1(new_n761), .A2(G106gat), .A3(new_n574), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n791), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G106gat), .B1(new_n804), .B2(new_n574), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n716), .A2(new_n652), .A3(new_n397), .A4(new_n783), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n809), .A2(new_n820), .B1(new_n825), .B2(G106gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n826), .B2(new_n823), .ZN(G1339gat));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n621), .B2(new_n624), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n647), .B1(new_n646), .B2(new_n622), .ZN(new_n830));
  AOI211_X1 g629(.A(KEYINPUT98), .B(new_n626), .C1(new_n644), .C2(new_n645), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n650), .B1(new_n625), .B2(new_n828), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n323), .A2(new_n834), .A3(new_n651), .A4(new_n332), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  INV_X1    g635(.A(new_n829), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n642), .B2(new_n648), .ZN(new_n838));
  INV_X1    g637(.A(new_n833), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n661), .A2(new_n663), .B1(new_n662), .B2(new_n671), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n678), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n673), .B2(new_n680), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT115), .B1(new_n835), .B2(new_n845), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n615), .B(new_n629), .C1(new_n642), .C2(new_n648), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n838), .A2(new_n839), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n833), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n843), .B1(new_n850), .B2(new_n836), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n708), .A2(new_n849), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n782), .A2(new_n840), .A3(new_n651), .A4(new_n834), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n652), .A2(new_n844), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n711), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n718), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n759), .B2(new_n652), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n333), .A2(new_n761), .A3(KEYINPUT114), .A4(new_n683), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n686), .ZN(new_n865));
  INV_X1    g664(.A(new_n577), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n566), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n683), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(new_n436), .ZN(G1340gat));
  NOR2_X1   g668(.A1(new_n867), .A2(new_n761), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(new_n434), .ZN(G1341gat));
  INV_X1    g670(.A(new_n718), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n867), .A2(new_n246), .A3(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n867), .A2(new_n261), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n246), .ZN(G1342gat));
  NOR2_X1   g674(.A1(new_n867), .A2(new_n711), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n452), .A2(new_n454), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n880));
  INV_X1    g679(.A(new_n876), .ZN(new_n881));
  INV_X1    g680(.A(new_n878), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT56), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(G134gat), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n876), .A2(new_n885), .A3(new_n877), .A4(new_n878), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n880), .A2(new_n883), .A3(new_n884), .A4(new_n886), .ZN(G1343gat));
  OAI21_X1  g686(.A(KEYINPUT117), .B1(new_n838), .B2(new_n839), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n832), .A2(new_n889), .A3(new_n833), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n890), .A3(new_n836), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n849), .A3(new_n782), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n856), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n711), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n758), .B1(new_n894), .B2(new_n854), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n397), .B1(new_n895), .B2(new_n863), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT57), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n861), .A2(new_n862), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n846), .A2(new_n853), .B1(new_n857), .B2(new_n711), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n718), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n397), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n740), .A2(new_n686), .A3(new_n515), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n897), .A2(new_n782), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(G141gat), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n864), .B2(new_n686), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n740), .A2(new_n574), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n900), .A2(KEYINPUT118), .A3(new_n573), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR4_X1   g709(.A1(new_n910), .A2(G141gat), .A3(new_n683), .A4(new_n515), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT58), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n683), .A2(G141gat), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n907), .A2(KEYINPUT119), .A3(new_n908), .A4(new_n909), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n914), .A2(new_n566), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT58), .B1(new_n904), .B2(G141gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n912), .A2(new_n919), .ZN(G1344gat));
  NOR2_X1   g719(.A1(new_n761), .A2(G148gat), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n914), .A2(new_n566), .A3(new_n916), .A4(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n900), .A2(new_n397), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT57), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n708), .B1(new_n892), .B2(new_n856), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n835), .A2(new_n845), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n261), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n759), .A2(new_n652), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT57), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n397), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n925), .A2(new_n652), .A3(new_n903), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n346), .B1(new_n933), .B2(KEYINPUT120), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n924), .A2(KEYINPUT57), .B1(new_n931), .B2(new_n397), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n935), .A2(new_n936), .A3(new_n652), .A4(new_n903), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n923), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n897), .A2(new_n902), .A3(new_n903), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n923), .B1(new_n939), .B2(new_n761), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(new_n346), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n922), .B1(new_n938), .B2(new_n941), .ZN(G1345gat));
  NOR3_X1   g741(.A1(new_n939), .A2(new_n359), .A3(new_n872), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n914), .A2(new_n566), .A3(new_n758), .A4(new_n916), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n359), .ZN(G1346gat));
  AND2_X1   g744(.A1(new_n897), .A2(new_n903), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n946), .A2(KEYINPUT121), .A3(new_n708), .A4(new_n902), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n948), .B1(new_n939), .B2(new_n711), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n342), .A3(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n914), .A2(new_n566), .A3(new_n708), .A4(new_n916), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n342), .ZN(G1347gat));
  NAND4_X1  g751(.A1(new_n900), .A2(new_n686), .A3(new_n515), .A4(new_n866), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(new_n683), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(new_n415), .ZN(G1348gat));
  NAND4_X1  g754(.A1(new_n900), .A2(new_n686), .A3(new_n866), .A4(new_n766), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n957), .A3(G176gat), .ZN(new_n958));
  XOR2_X1   g757(.A(KEYINPUT122), .B(G176gat), .Z(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n956), .B2(new_n959), .ZN(G1349gat));
  OAI211_X1 g759(.A(new_n686), .B(new_n866), .C1(new_n859), .C2(new_n863), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(new_n566), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(KEYINPUT124), .A3(new_n718), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(new_n953), .B2(new_n872), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(new_n965), .A3(G183gat), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n961), .A2(new_n408), .A3(new_n566), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(new_n758), .ZN(new_n971));
  NOR4_X1   g770(.A1(new_n953), .A2(KEYINPUT123), .A3(new_n408), .A4(new_n261), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT60), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n962), .A2(new_n407), .A3(new_n758), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT123), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n970), .A2(new_n969), .A3(new_n758), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT60), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n978), .A2(new_n967), .A3(new_n979), .A4(new_n966), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n974), .A2(new_n980), .ZN(G1350gat));
  XNOR2_X1  g780(.A(KEYINPUT61), .B(G190gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n953), .A2(new_n711), .ZN(new_n984));
  MUX2_X1   g783(.A(new_n982), .B(new_n983), .S(new_n984), .Z(G1351gat));
  NOR3_X1   g784(.A1(new_n740), .A2(new_n573), .A3(new_n566), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n935), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(KEYINPUT126), .A3(new_n782), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n935), .A2(new_n782), .A3(new_n986), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n988), .A2(new_n991), .A3(G197gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n986), .A2(new_n900), .A3(new_n397), .ZN(new_n993));
  OR3_X1    g792(.A1(new_n993), .A2(G197gat), .A3(new_n683), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(G1352gat));
  NAND2_X1  g794(.A1(new_n908), .A2(new_n766), .ZN(new_n996));
  NOR4_X1   g795(.A1(new_n996), .A2(new_n864), .A3(G204gat), .A4(new_n573), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT62), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n935), .A2(new_n652), .A3(new_n986), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G204gat), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1000), .ZN(G1353gat));
  NAND4_X1  g800(.A1(new_n925), .A2(new_n758), .A3(new_n932), .A4(new_n986), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(G211gat), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT63), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1002), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(new_n993), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1008), .A2(new_n369), .A3(new_n758), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1003), .A2(new_n1010), .A3(new_n1004), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1011), .ZN(G1354gat));
  AOI21_X1  g811(.A(G218gat), .B1(new_n1008), .B2(new_n708), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n711), .A2(new_n370), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1013), .B1(new_n987), .B2(new_n1014), .ZN(G1355gat));
endmodule


