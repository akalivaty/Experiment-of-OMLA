//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT68), .B(G116), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G119), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT2), .A2(G113), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT2), .A2(G113), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT67), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT2), .A2(G113), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT69), .B1(new_n191), .B2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT68), .A2(G116), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT68), .A2(G116), .ZN(new_n204));
  OAI21_X1  g018(.A(G119), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(new_n188), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n194), .A4(new_n200), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n191), .A2(new_n197), .A3(new_n199), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n202), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G104), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT3), .B1(new_n214), .B2(G107), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(G107), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G101), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n219), .B(new_n213), .C1(new_n215), .C2(new_n216), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n222), .A3(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT85), .B1(new_n210), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(G110), .B(G122), .Z(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n221), .A2(new_n223), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n202), .A2(new_n208), .A3(new_n209), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n212), .A2(G104), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n216), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n220), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT5), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n196), .B1(new_n189), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n206), .B2(new_n236), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n238), .A3(new_n209), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n225), .A2(new_n227), .A3(new_n231), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT86), .ZN(new_n241));
  INV_X1    g055(.A(new_n239), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n228), .A2(new_n230), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(KEYINPUT85), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n227), .A4(new_n231), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n238), .A2(new_n209), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n234), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n239), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n226), .B(KEYINPUT8), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G224), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT7), .B1(new_n254), .B2(G953), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n260), .A2(KEYINPUT1), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n258), .B2(G146), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n258), .C2(G146), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(G128), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n262), .B1(new_n260), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G125), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n272), .A2(new_n257), .A3(new_n259), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(KEYINPUT0), .B2(G128), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT0), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n261), .A3(KEYINPUT64), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n260), .A2(new_n271), .A3(new_n276), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G125), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n255), .B1(new_n270), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n270), .A2(new_n281), .A3(new_n255), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n253), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n247), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n284), .B1(new_n241), .B2(new_n246), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT88), .B1(new_n290), .B2(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n227), .B1(new_n244), .B2(new_n231), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n293), .A2(KEYINPUT6), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n241), .B2(new_n246), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n270), .A2(new_n281), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n254), .A2(G953), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(KEYINPUT87), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n298), .B(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G210), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n292), .A2(new_n305), .A3(new_n303), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n305), .B1(new_n292), .B2(new_n303), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT89), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT78), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G221), .B1(new_n317), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(new_n288), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n278), .A2(new_n276), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n272), .B1(new_n257), .B2(new_n259), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n273), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n221), .A2(new_n324), .A3(new_n223), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT79), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n221), .A2(new_n327), .A3(new_n324), .A4(new_n223), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G137), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT65), .B1(new_n330), .B2(G134), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT11), .ZN(new_n332));
  OAI22_X1  g146(.A1(new_n331), .A2(new_n332), .B1(G134), .B2(new_n330), .ZN(new_n333));
  AOI211_X1 g147(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n330), .C2(G134), .ZN(new_n334));
  OAI21_X1  g148(.A(G131), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n330), .A2(G134), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT65), .ZN(new_n337));
  INV_X1    g151(.A(G134), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(G137), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n336), .B1(new_n339), .B2(KEYINPUT11), .ZN(new_n340));
  INV_X1    g154(.A(G131), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n331), .A2(new_n332), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n263), .A2(G128), .B1(new_n257), .B2(new_n259), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n220), .B(new_n233), .C1(new_n262), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n234), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n266), .A2(G128), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT66), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n260), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n257), .A2(new_n259), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G128), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n353), .A2(KEYINPUT71), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT71), .B1(new_n353), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n329), .A2(new_n345), .A3(new_n349), .A4(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G110), .B(G140), .ZN(new_n361));
  INV_X1    g175(.A(G953), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(G227), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n361), .B(new_n363), .Z(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(KEYINPUT83), .A3(new_n364), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n353), .A2(new_n356), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n347), .B1(new_n370), .B2(new_n235), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT12), .A3(new_n344), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT12), .B1(new_n371), .B2(new_n344), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n374), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT82), .A3(new_n372), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n367), .A2(new_n368), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n365), .A2(new_n366), .B1(new_n375), .B2(new_n377), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT84), .A3(new_n368), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n326), .A2(new_n328), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n359), .A2(new_n349), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n344), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT80), .B(new_n344), .C1(new_n385), .C2(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n360), .ZN(new_n392));
  INV_X1    g206(.A(new_n364), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(G902), .B1(new_n384), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n321), .B1(new_n395), .B2(new_n320), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n360), .A3(new_n364), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n360), .B1(new_n373), .B2(new_n374), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n393), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n397), .A2(KEYINPUT81), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT81), .B1(new_n397), .B2(new_n399), .ZN(new_n401));
  OAI21_X1  g215(.A(G469), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n319), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n362), .A2(G952), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(G234), .B2(G237), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI211_X1 g220(.A(new_n288), .B(new_n362), .C1(G234), .C2(G237), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT21), .B(G898), .Z(new_n409));
  OAI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G214), .B1(G237), .B2(G902), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n190), .A2(G122), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT97), .B1(new_n413), .B2(KEYINPUT14), .ZN(new_n414));
  INV_X1    g228(.A(G122), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G116), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT94), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(KEYINPUT14), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n413), .A2(KEYINPUT97), .A3(KEYINPUT14), .ZN(new_n420));
  OAI21_X1  g234(.A(G107), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n212), .A3(new_n413), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n258), .A2(KEYINPUT95), .A3(G128), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT95), .B1(new_n258), .B2(G128), .ZN(new_n424));
  OAI22_X1  g238(.A1(new_n423), .A2(new_n424), .B1(G128), .B2(new_n258), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G134), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n425), .A2(G134), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n421), .B(new_n422), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n423), .A2(new_n424), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n429), .A2(KEYINPUT13), .B1(new_n261), .B2(G143), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT96), .B1(new_n429), .B2(KEYINPUT13), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n429), .A2(KEYINPUT96), .A3(KEYINPUT13), .ZN(new_n433));
  OAI21_X1  g247(.A(G134), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n417), .A2(new_n413), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G107), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n426), .B1(new_n436), .B2(new_n422), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G217), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n317), .A2(new_n440), .A3(G953), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n428), .A2(new_n438), .A3(new_n441), .ZN(new_n444));
  AOI21_X1  g258(.A(G902), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G478), .ZN(new_n446));
  OAI22_X1  g260(.A1(new_n445), .A2(KEYINPUT98), .B1(KEYINPUT15), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT98), .ZN(new_n448));
  INV_X1    g262(.A(new_n445), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n445), .B(KEYINPUT98), .C1(KEYINPUT15), .C2(new_n446), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G237), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n362), .A3(G214), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n258), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G131), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT18), .ZN(new_n457));
  OR3_X1    g271(.A1(new_n456), .A2(KEYINPUT90), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT90), .B1(new_n456), .B2(new_n457), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n454), .B(G143), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  XNOR2_X1  g275(.A(G125), .B(G140), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G146), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n256), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n460), .A2(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n458), .A2(new_n459), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n462), .A2(KEYINPUT16), .ZN(new_n468));
  OR3_X1    g282(.A1(new_n269), .A2(KEYINPUT16), .A3(G140), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(G146), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(G146), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n455), .A2(KEYINPUT17), .A3(G131), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n460), .A2(new_n341), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n456), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n473), .B(new_n474), .C1(new_n476), .C2(KEYINPUT17), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G113), .B(G122), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(new_n214), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT92), .Z(new_n481));
  NOR2_X1   g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT19), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  MUX2_X1   g301(.A(new_n485), .B(new_n487), .S(new_n462), .Z(new_n488));
  OAI211_X1 g302(.A(new_n476), .B(new_n470), .C1(G146), .C2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n480), .B1(new_n467), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(G475), .A2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OR3_X1    g307(.A1(new_n491), .A2(KEYINPUT20), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT20), .B1(new_n491), .B2(new_n493), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n480), .B1(new_n467), .B2(new_n477), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n288), .B1(new_n482), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT93), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n478), .A2(new_n481), .ZN(new_n500));
  INV_X1    g314(.A(new_n497), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n504), .A3(G475), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n452), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n314), .A2(new_n403), .A3(new_n412), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n453), .A2(new_n362), .A3(G210), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n219), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n511));
  XOR2_X1   g325(.A(new_n510), .B(new_n511), .Z(new_n512));
  INV_X1    g326(.A(KEYINPUT72), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n210), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n230), .A2(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n333), .A2(G131), .A3(new_n334), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n341), .B1(new_n340), .B2(new_n342), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n324), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT70), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n344), .A2(new_n521), .A3(new_n324), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n338), .A2(G137), .ZN(new_n524));
  OAI21_X1  g338(.A(G131), .B1(new_n524), .B2(new_n336), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n343), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n357), .B2(new_n358), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n516), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n268), .A2(new_n526), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n280), .B1(new_n343), .B2(new_n335), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT30), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n520), .A3(new_n522), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n533), .B2(KEYINPUT30), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n512), .B(new_n529), .C1(new_n534), .C2(new_n210), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT73), .B1(new_n535), .B2(KEYINPUT31), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(KEYINPUT73), .A3(KEYINPUT31), .ZN(new_n539));
  INV_X1    g353(.A(new_n515), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n230), .A2(KEYINPUT72), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n528), .B(new_n519), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT28), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n528), .A2(new_n520), .A3(new_n522), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n519), .B1(new_n268), .B2(new_n526), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n545), .A2(new_n516), .B1(new_n230), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n544), .B1(new_n547), .B2(new_n543), .ZN(new_n548));
  INV_X1    g362(.A(new_n512), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n538), .A2(new_n539), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G472), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n288), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT32), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n551), .A2(KEYINPUT32), .A3(new_n552), .A4(new_n288), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n534), .A2(new_n210), .ZN(new_n557));
  INV_X1    g371(.A(new_n529), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n549), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT29), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n512), .B(new_n544), .C1(new_n547), .C2(new_n543), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT74), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n559), .A2(new_n561), .A3(KEYINPUT74), .A4(new_n560), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n544), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n549), .A2(new_n560), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n531), .B1(new_n514), .B2(new_n515), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT28), .B1(new_n569), .B2(new_n528), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n533), .A2(new_n515), .A3(new_n514), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n529), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n572), .B2(KEYINPUT28), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n567), .B(new_n568), .C1(new_n573), .C2(new_n566), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n564), .A2(new_n288), .A3(new_n565), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G472), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n555), .A2(new_n556), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n440), .B1(G234), .B2(new_n288), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(G119), .B2(new_n261), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n187), .A2(KEYINPUT23), .A3(G128), .ZN(new_n582));
  OAI22_X1  g396(.A1(new_n581), .A2(new_n582), .B1(G119), .B2(new_n261), .ZN(new_n583));
  XNOR2_X1  g397(.A(G119), .B(G128), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT24), .B(G110), .Z(new_n585));
  OAI22_X1  g399(.A1(new_n583), .A2(G110), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n465), .A3(new_n470), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT76), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n586), .A2(new_n589), .A3(new_n465), .A4(new_n470), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n583), .A2(G110), .B1(new_n584), .B2(new_n585), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n471), .B2(new_n472), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT22), .B(G137), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n362), .A2(G221), .A3(G234), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n588), .A2(new_n592), .A3(new_n590), .A4(new_n596), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n288), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n598), .A2(KEYINPUT25), .A3(new_n288), .A4(new_n599), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n579), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n598), .A2(new_n599), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n578), .A2(G902), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT77), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n577), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n508), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n219), .ZN(G3));
  INV_X1    g426(.A(new_n411), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n307), .B2(new_n309), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n614), .A2(new_n410), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n552), .B1(new_n551), .B2(new_n288), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n553), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(new_n403), .A3(new_n609), .ZN(new_n621));
  INV_X1    g435(.A(new_n506), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n443), .A2(new_n444), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT33), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n446), .A2(G902), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n449), .A2(KEYINPUT100), .A3(new_n446), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n445), .B2(G478), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n629), .A2(new_n630), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NOR4_X1   g448(.A1(new_n616), .A2(new_n621), .A3(new_n622), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT34), .B(G104), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND2_X1  g451(.A1(new_n622), .A2(new_n452), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n621), .A2(new_n616), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n212), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NAND4_X1  g456(.A1(new_n314), .A2(new_n403), .A3(new_n412), .A4(new_n620), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n602), .A2(new_n603), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n578), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n597), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n593), .B(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n648), .A2(G902), .A3(new_n578), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n644), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n604), .A2(new_n649), .A3(KEYINPUT102), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n507), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n643), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT37), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NOR2_X1   g470(.A1(new_n651), .A2(new_n652), .ZN(new_n657));
  AOI211_X1 g471(.A(new_n613), .B(new_n657), .C1(new_n307), .C2(new_n309), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n405), .B1(new_n407), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n638), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n403), .A2(new_n658), .A3(new_n577), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n314), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n314), .A2(new_n664), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n452), .A2(new_n506), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n668), .A2(new_n613), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n604), .A2(new_n649), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n535), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n549), .B2(new_n572), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n674), .B2(G902), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n555), .A2(new_n556), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n403), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n660), .B(KEYINPUT39), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n681));
  AOI211_X1 g495(.A(new_n672), .B(new_n677), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n670), .B(new_n682), .C1(new_n681), .C2(new_n680), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  INV_X1    g498(.A(new_n660), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n631), .A2(new_n633), .ZN(new_n686));
  INV_X1    g500(.A(new_n630), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n627), .B2(new_n628), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n506), .B(new_n685), .C1(new_n686), .C2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n403), .A2(new_n658), .A3(new_n577), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NOR2_X1   g506(.A1(new_n622), .A2(new_n634), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n615), .A2(new_n609), .A3(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n381), .A2(new_n383), .B1(new_n392), .B2(new_n393), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n379), .A2(new_n380), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT84), .B1(new_n382), .B2(new_n368), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n394), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n320), .A3(new_n288), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n696), .A2(new_n700), .A3(new_n318), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n696), .A2(new_n700), .A3(KEYINPUT104), .A4(new_n318), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n703), .A2(new_n577), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n694), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n615), .A2(new_n577), .A3(new_n703), .A4(new_n704), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n609), .A2(new_n622), .A3(new_n452), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(G116), .Z(G18));
  NOR2_X1   g526(.A1(new_n709), .A2(new_n653), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n187), .ZN(G21));
  NAND4_X1  g528(.A1(new_n614), .A2(new_n410), .A3(new_n506), .A4(new_n452), .ZN(new_n715));
  NOR2_X1   g529(.A1(G472), .A2(G902), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n567), .B1(new_n573), .B2(new_n566), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT105), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n720), .B(new_n567), .C1(new_n573), .C2(new_n566), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n549), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n535), .B(KEYINPUT31), .Z(new_n723));
  AOI21_X1  g537(.A(new_n717), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n608), .A3(new_n618), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n715), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n703), .A2(new_n704), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NOR4_X1   g544(.A1(new_n724), .A2(new_n689), .A3(new_n617), .A4(new_n671), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(KEYINPUT106), .A3(new_n614), .A4(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n703), .A2(new_n614), .A3(new_n704), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n724), .A2(new_n617), .A3(new_n671), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n690), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n733), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n292), .A2(new_n305), .A3(new_n303), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n311), .A3(KEYINPUT89), .ZN(new_n742));
  INV_X1    g556(.A(new_n312), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n411), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n610), .ZN(new_n747));
  INV_X1    g561(.A(new_n321), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n397), .A2(new_n399), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(G469), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n700), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n700), .A2(KEYINPUT107), .A3(new_n748), .A4(new_n751), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n319), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n313), .A2(KEYINPUT108), .A3(new_n411), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n746), .A2(new_n747), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n740), .B1(new_n758), .B2(new_n689), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n689), .A2(new_n740), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n577), .A2(new_n608), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n746), .A2(new_n761), .A3(new_n757), .A4(new_n756), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  INV_X1    g580(.A(new_n661), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n338), .ZN(G36));
  NOR2_X1   g583(.A1(new_n634), .A2(new_n506), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT43), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n634), .B2(new_n506), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n619), .A3(new_n672), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT44), .Z(new_n776));
  NAND2_X1  g590(.A1(new_n746), .A2(new_n757), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT45), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n320), .B1(new_n750), .B2(KEYINPUT45), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n321), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT46), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n781), .B2(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n700), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n318), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n679), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n778), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT111), .B(G137), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G39));
  NAND2_X1  g605(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT108), .B1(new_n313), .B2(new_n411), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n745), .B(new_n613), .C1(new_n310), .C2(new_n312), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n786), .A2(new_n796), .A3(new_n318), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n577), .A2(new_n609), .A3(new_n689), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n792), .A2(new_n795), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  AND4_X1   g614(.A1(new_n608), .A2(new_n770), .A3(new_n318), .A4(new_n411), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n696), .A2(new_n700), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n801), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n668), .A3(new_n677), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n666), .A2(new_n667), .A3(new_n411), .ZN(new_n810));
  INV_X1    g624(.A(new_n728), .ZN(new_n811));
  INV_X1    g625(.A(new_n726), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n406), .B1(new_n771), .B2(new_n773), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n810), .A2(KEYINPUT50), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT50), .B1(new_n810), .B2(new_n815), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT116), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n818), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n777), .A2(new_n811), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n813), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(KEYINPUT117), .A3(new_n813), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n735), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n609), .A2(new_n824), .A3(new_n405), .A4(new_n677), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n622), .A3(new_n634), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n823), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT118), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n777), .A2(new_n814), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n792), .A2(new_n797), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT115), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n696), .A2(new_n700), .A3(new_n319), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n837), .A2(KEYINPUT115), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n834), .A2(KEYINPUT118), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n809), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n553), .A2(new_n693), .A3(new_n618), .A4(new_n609), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n314), .A3(new_n403), .A4(new_n412), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n508), .B2(new_n610), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT113), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n848), .B(new_n851), .C1(new_n508), .C2(new_n610), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n709), .A2(new_n643), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n653), .A2(new_n710), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n694), .A2(new_n705), .B1(new_n728), .B2(new_n727), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n403), .A2(new_n577), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n653), .A2(new_n660), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n859), .A2(new_n860), .B1(new_n756), .B2(new_n731), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n861), .A2(new_n777), .B1(new_n758), .B2(new_n767), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n765), .A2(new_n853), .A3(new_n858), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n662), .A2(new_n691), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n614), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n867), .A2(new_n660), .A3(new_n669), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n671), .A3(new_n676), .A4(new_n756), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n738), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT52), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n865), .B1(new_n732), .B2(new_n737), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n869), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n846), .B1(new_n864), .B2(new_n875), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n873), .A2(new_n738), .A3(new_n866), .A4(new_n869), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n873), .B1(new_n872), .B2(new_n869), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n856), .A2(new_n857), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n850), .B2(new_n852), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT109), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n795), .A2(new_n883), .A3(new_n756), .A4(new_n761), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n862), .B1(new_n885), .B2(new_n759), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n879), .A2(KEYINPUT53), .A3(new_n881), .A4(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n876), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT114), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n876), .A2(new_n891), .A3(new_n887), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT114), .B(new_n846), .C1(new_n864), .C2(new_n875), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT54), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n837), .A2(new_n839), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT119), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n837), .A2(new_n898), .A3(new_n839), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n836), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n809), .B1(new_n820), .B2(new_n816), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n831), .A3(new_n833), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n577), .A2(new_n608), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n827), .B2(new_n829), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT48), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n904), .B2(new_n905), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n814), .A2(new_n734), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n404), .B(new_n910), .C1(new_n832), .C2(new_n693), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n906), .A2(new_n908), .ZN(new_n912));
  AND4_X1   g726(.A1(new_n902), .A2(new_n909), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n845), .A2(new_n895), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n808), .B1(new_n914), .B2(new_n915), .ZN(G75));
  NAND2_X1  g730(.A1(new_n892), .A2(new_n893), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n288), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(G210), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n297), .B(new_n301), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n362), .A2(G952), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G51));
  AND3_X1   g740(.A1(new_n892), .A2(KEYINPUT54), .A3(new_n893), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n894), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n321), .B(KEYINPUT57), .Z(new_n929));
  OAI21_X1  g743(.A(new_n699), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n918), .A2(new_n779), .A3(new_n780), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n933), .A2(new_n491), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n491), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n925), .ZN(G60));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  INV_X1    g751(.A(new_n629), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n917), .A2(new_n889), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n892), .A2(KEYINPUT54), .A3(new_n893), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n937), .B1(new_n945), .B2(new_n925), .ZN(new_n946));
  INV_X1    g760(.A(new_n925), .ZN(new_n947));
  OAI211_X1 g761(.A(KEYINPUT121), .B(new_n947), .C1(new_n928), .C2(new_n942), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n938), .B1(new_n895), .B2(new_n940), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n892), .A2(new_n893), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n954), .A2(new_n605), .ZN(new_n955));
  NOR2_X1   g769(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n925), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n954), .B2(new_n648), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G66));
  INV_X1    g775(.A(new_n409), .ZN(new_n962));
  OAI21_X1  g776(.A(G953), .B1(new_n962), .B2(new_n254), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n881), .B2(G953), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  INV_X1    g779(.A(new_n297), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(G898), .B2(new_n362), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  AOI21_X1  g782(.A(new_n362), .B1(G227), .B2(G900), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n903), .A2(new_n867), .A3(new_n669), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n788), .B1(new_n778), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n768), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n973), .A2(new_n974), .A3(new_n799), .A4(new_n872), .ZN(new_n975));
  INV_X1    g789(.A(new_n765), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n362), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n659), .A2(G953), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n977), .B2(new_n979), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n534), .B(new_n488), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n683), .A2(new_n872), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n638), .B1(new_n622), .B2(new_n634), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n795), .A2(new_n747), .A3(new_n680), .A4(new_n988), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT124), .Z(new_n990));
  AND3_X1   g804(.A1(new_n990), .A2(new_n789), .A3(new_n799), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n982), .B1(new_n992), .B2(new_n362), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n970), .B(new_n971), .C1(new_n984), .C2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n981), .A2(new_n983), .ZN(new_n995));
  INV_X1    g809(.A(new_n980), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n993), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT126), .A4(new_n969), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n994), .A2(new_n999), .ZN(G72));
  NOR2_X1   g814(.A1(new_n557), .A2(new_n558), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT127), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n987), .A2(new_n881), .A3(new_n991), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  AOI211_X1 g819(.A(new_n549), .B(new_n1002), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1005), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n1007), .B(new_n888), .C1(new_n535), .C2(new_n559), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n975), .A2(new_n976), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1007), .B1(new_n1009), .B2(new_n881), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1002), .A2(new_n549), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n947), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1006), .A2(new_n1008), .A3(new_n1012), .ZN(G57));
endmodule


