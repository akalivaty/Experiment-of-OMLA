

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U547 ( .A1(n902), .A2(n728), .ZN(n727) );
  BUF_X1 U548 ( .A(n861), .Z(n512) );
  NOR2_X1 U549 ( .A1(n519), .A2(G2105), .ZN(n861) );
  NOR2_X1 U550 ( .A1(n533), .A2(n532), .ZN(G160) );
  AND2_X1 U551 ( .A1(G2105), .A2(n519), .ZN(n864) );
  NOR2_X1 U552 ( .A1(n525), .A2(n524), .ZN(G164) );
  NAND2_X1 U553 ( .A1(n752), .A2(G1341), .ZN(n513) );
  INV_X1 U554 ( .A(KEYINPUT101), .ZN(n745) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n702) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n514) );
  XNOR2_X2 U558 ( .A(n514), .B(KEYINPUT65), .ZN(n866) );
  NAND2_X1 U559 ( .A1(n866), .A2(G114), .ZN(n515) );
  XOR2_X1 U560 ( .A(KEYINPUT87), .B(n515), .Z(n517) );
  XOR2_X1 U561 ( .A(KEYINPUT64), .B(G2104), .Z(n519) );
  NAND2_X1 U562 ( .A1(n864), .A2(G126), .ZN(n516) );
  NAND2_X1 U563 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U564 ( .A(n518), .B(KEYINPUT88), .ZN(n525) );
  NAND2_X1 U565 ( .A1(n512), .A2(G102), .ZN(n523) );
  XNOR2_X1 U566 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n521) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XNOR2_X1 U568 ( .A(n521), .B(n520), .ZN(n860) );
  NAND2_X1 U569 ( .A1(n860), .A2(G138), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U571 ( .A1(G113), .A2(n866), .ZN(n526) );
  XNOR2_X1 U572 ( .A(n526), .B(KEYINPUT66), .ZN(n529) );
  NAND2_X1 U573 ( .A1(G101), .A2(n861), .ZN(n527) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n527), .Z(n528) );
  NAND2_X1 U575 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U576 ( .A1(G125), .A2(n864), .ZN(n531) );
  NAND2_X1 U577 ( .A1(G137), .A2(n860), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U579 ( .A(G651), .ZN(n537) );
  NOR2_X1 U580 ( .A1(G543), .A2(n537), .ZN(n534) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n534), .Z(n637) );
  NAND2_X1 U582 ( .A1(G64), .A2(n637), .ZN(n536) );
  XOR2_X1 U583 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  NOR2_X2 U584 ( .A1(G651), .A2(n622), .ZN(n646) );
  NAND2_X1 U585 ( .A1(G52), .A2(n646), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n542) );
  NOR2_X1 U587 ( .A1(n622), .A2(n537), .ZN(n641) );
  NAND2_X1 U588 ( .A1(G77), .A2(n641), .ZN(n539) );
  NAND2_X1 U589 ( .A1(G90), .A2(n638), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U592 ( .A1(n542), .A2(n541), .ZN(G171) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U594 ( .A1(G123), .A2(n864), .ZN(n543) );
  XNOR2_X1 U595 ( .A(n543), .B(KEYINPUT18), .ZN(n550) );
  NAND2_X1 U596 ( .A1(G111), .A2(n866), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G135), .A2(n860), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G99), .A2(n512), .ZN(n546) );
  XNOR2_X1 U600 ( .A(KEYINPUT79), .B(n546), .ZN(n547) );
  NOR2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U603 ( .A(KEYINPUT80), .B(n551), .ZN(n956) );
  XNOR2_X1 U604 ( .A(n956), .B(G2096), .ZN(n552) );
  OR2_X1 U605 ( .A1(G2100), .A2(n552), .ZN(G156) );
  INV_X1 U606 ( .A(G57), .ZN(G237) );
  INV_X1 U607 ( .A(G132), .ZN(G219) );
  INV_X1 U608 ( .A(G82), .ZN(G220) );
  XOR2_X1 U609 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n554) );
  NAND2_X1 U610 ( .A1(G7), .A2(G661), .ZN(n553) );
  XNOR2_X1 U611 ( .A(n554), .B(n553), .ZN(G223) );
  INV_X1 U612 ( .A(G223), .ZN(n820) );
  NAND2_X1 U613 ( .A1(n820), .A2(G567), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  NAND2_X1 U615 ( .A1(G56), .A2(n637), .ZN(n556) );
  XOR2_X1 U616 ( .A(KEYINPUT14), .B(n556), .Z(n562) );
  NAND2_X1 U617 ( .A1(n638), .A2(G81), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT12), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G68), .A2(n641), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U621 ( .A(KEYINPUT13), .B(n560), .Z(n561) );
  NOR2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n646), .A2(G43), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n921) );
  INV_X1 U625 ( .A(G860), .ZN(n598) );
  OR2_X1 U626 ( .A1(n921), .A2(n598), .ZN(G153) );
  INV_X1 U627 ( .A(G171), .ZN(G301) );
  NAND2_X1 U628 ( .A1(G868), .A2(G301), .ZN(n574) );
  NAND2_X1 U629 ( .A1(G92), .A2(n638), .ZN(n571) );
  NAND2_X1 U630 ( .A1(G66), .A2(n637), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G79), .A2(n641), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n646), .A2(G54), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT76), .B(n567), .Z(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT15), .ZN(n902) );
  OR2_X1 U638 ( .A1(n902), .A2(G868), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(G284) );
  NAND2_X1 U640 ( .A1(G63), .A2(n637), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G51), .A2(n646), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT6), .B(n577), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n638), .A2(G89), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT4), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G76), .A2(n641), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(KEYINPUT5), .B(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(KEYINPUT77), .B(n582), .ZN(n583) );
  NOR2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT7), .B(n585), .Z(G168) );
  XOR2_X1 U652 ( .A(G168), .B(KEYINPUT8), .Z(n586) );
  XNOR2_X1 U653 ( .A(KEYINPUT78), .B(n586), .ZN(G286) );
  NAND2_X1 U654 ( .A1(n646), .A2(G53), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT72), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G65), .A2(n637), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT73), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G78), .A2(n641), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G91), .A2(n638), .ZN(n593) );
  XNOR2_X1 U662 ( .A(KEYINPUT71), .B(n593), .ZN(n594) );
  NOR2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n920) );
  XOR2_X1 U664 ( .A(n920), .B(KEYINPUT74), .Z(G299) );
  NAND2_X1 U665 ( .A1(G868), .A2(G286), .ZN(n597) );
  INV_X1 U666 ( .A(G868), .ZN(n658) );
  NAND2_X1 U667 ( .A1(G299), .A2(n658), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n599), .A2(n902), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n921), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G868), .A2(n902), .ZN(n601) );
  NOR2_X1 U674 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U675 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G559), .A2(n902), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(n921), .ZN(n654) );
  NOR2_X1 U678 ( .A1(n654), .A2(G860), .ZN(n612) );
  NAND2_X1 U679 ( .A1(G67), .A2(n637), .ZN(n606) );
  NAND2_X1 U680 ( .A1(G55), .A2(n646), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G80), .A2(n641), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G93), .A2(n638), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U685 ( .A(KEYINPUT81), .B(n609), .Z(n610) );
  OR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n657) );
  XOR2_X1 U687 ( .A(n612), .B(n657), .Z(G145) );
  NAND2_X1 U688 ( .A1(n637), .A2(G62), .ZN(n619) );
  NAND2_X1 U689 ( .A1(G75), .A2(n641), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G88), .A2(n638), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n646), .A2(G50), .ZN(n615) );
  XOR2_X1 U693 ( .A(KEYINPUT84), .B(n615), .Z(n616) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U696 ( .A(KEYINPUT85), .B(n620), .Z(G303) );
  INV_X1 U697 ( .A(G303), .ZN(G166) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n621), .B(KEYINPUT82), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G49), .A2(n646), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G87), .A2(n622), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n637), .A2(n625), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(G288) );
  NAND2_X1 U705 ( .A1(n637), .A2(G60), .ZN(n628) );
  XOR2_X1 U706 ( .A(KEYINPUT69), .B(n628), .Z(n630) );
  NAND2_X1 U707 ( .A1(n646), .A2(G47), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U709 ( .A(KEYINPUT70), .B(n631), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G72), .A2(n641), .ZN(n632) );
  XOR2_X1 U711 ( .A(KEYINPUT68), .B(n632), .Z(n633) );
  NOR2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n638), .A2(G85), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U715 ( .A1(G61), .A2(n637), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G86), .A2(n638), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n641), .A2(G73), .ZN(n642) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U721 ( .A(KEYINPUT83), .B(n645), .Z(n648) );
  NAND2_X1 U722 ( .A1(n646), .A2(G48), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(G305) );
  XNOR2_X1 U724 ( .A(G166), .B(G299), .ZN(n651) );
  XNOR2_X1 U725 ( .A(KEYINPUT19), .B(n657), .ZN(n649) );
  XNOR2_X1 U726 ( .A(G288), .B(n649), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(G290), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n653), .B(G305), .ZN(n828) );
  XNOR2_X1 U730 ( .A(n828), .B(n654), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n655), .A2(G868), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n656), .B(KEYINPUT86), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U739 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U741 ( .A1(G220), .A2(G219), .ZN(n665) );
  XOR2_X1 U742 ( .A(KEYINPUT22), .B(n665), .Z(n666) );
  NOR2_X1 U743 ( .A1(G218), .A2(n666), .ZN(n667) );
  NAND2_X1 U744 ( .A1(G96), .A2(n667), .ZN(n825) );
  NAND2_X1 U745 ( .A1(n825), .A2(G2106), .ZN(n671) );
  NAND2_X1 U746 ( .A1(G120), .A2(G108), .ZN(n668) );
  NOR2_X1 U747 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G69), .A2(n669), .ZN(n826) );
  NAND2_X1 U749 ( .A1(n826), .A2(G567), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n827) );
  NAND2_X1 U751 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U752 ( .A1(n827), .A2(n672), .ZN(n824) );
  NAND2_X1 U753 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U754 ( .A1(G160), .A2(G40), .ZN(n701) );
  NOR2_X1 U755 ( .A1(n702), .A2(n701), .ZN(n803) );
  NAND2_X1 U756 ( .A1(G117), .A2(n866), .ZN(n674) );
  NAND2_X1 U757 ( .A1(G129), .A2(n864), .ZN(n673) );
  NAND2_X1 U758 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n512), .A2(G105), .ZN(n675) );
  XOR2_X1 U760 ( .A(KEYINPUT38), .B(n675), .Z(n676) );
  NOR2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U762 ( .A1(n860), .A2(G141), .ZN(n678) );
  NAND2_X1 U763 ( .A1(n679), .A2(n678), .ZN(n857) );
  NAND2_X1 U764 ( .A1(G1996), .A2(n857), .ZN(n687) );
  NAND2_X1 U765 ( .A1(G107), .A2(n866), .ZN(n681) );
  NAND2_X1 U766 ( .A1(G119), .A2(n864), .ZN(n680) );
  NAND2_X1 U767 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G131), .A2(n860), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G95), .A2(n512), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n684) );
  OR2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n848) );
  NAND2_X1 U772 ( .A1(G1991), .A2(n848), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U774 ( .A(KEYINPUT90), .B(n688), .Z(n962) );
  INV_X1 U775 ( .A(n962), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n803), .A2(n689), .ZN(n791) );
  XNOR2_X1 U777 ( .A(G2067), .B(KEYINPUT37), .ZN(n801) );
  NAND2_X1 U778 ( .A1(n860), .A2(G140), .ZN(n690) );
  XOR2_X1 U779 ( .A(KEYINPUT89), .B(n690), .Z(n692) );
  NAND2_X1 U780 ( .A1(n512), .A2(G104), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U782 ( .A(KEYINPUT34), .B(n693), .ZN(n698) );
  NAND2_X1 U783 ( .A1(G116), .A2(n866), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G128), .A2(n864), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U786 ( .A(KEYINPUT35), .B(n696), .Z(n697) );
  NOR2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U788 ( .A(KEYINPUT36), .B(n699), .ZN(n852) );
  NOR2_X1 U789 ( .A1(n801), .A2(n852), .ZN(n965) );
  NAND2_X1 U790 ( .A1(n803), .A2(n965), .ZN(n799) );
  NAND2_X1 U791 ( .A1(n791), .A2(n799), .ZN(n700) );
  XOR2_X1 U792 ( .A(KEYINPUT91), .B(n700), .Z(n788) );
  INV_X1 U793 ( .A(n701), .ZN(n703) );
  NAND2_X2 U794 ( .A1(n703), .A2(n702), .ZN(n752) );
  NAND2_X1 U795 ( .A1(G8), .A2(n752), .ZN(n781) );
  NOR2_X1 U796 ( .A1(G1966), .A2(n781), .ZN(n744) );
  XOR2_X1 U797 ( .A(KEYINPUT25), .B(G2078), .Z(n933) );
  NOR2_X1 U798 ( .A1(n933), .A2(n752), .ZN(n704) );
  XNOR2_X1 U799 ( .A(n704), .B(KEYINPUT95), .ZN(n706) );
  XOR2_X1 U800 ( .A(G1961), .B(KEYINPUT94), .Z(n982) );
  NAND2_X1 U801 ( .A1(n982), .A2(n752), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n737) );
  NOR2_X1 U803 ( .A1(G171), .A2(n737), .ZN(n712) );
  NOR2_X1 U804 ( .A1(G2084), .A2(n752), .ZN(n747) );
  NOR2_X1 U805 ( .A1(n747), .A2(n744), .ZN(n707) );
  XNOR2_X1 U806 ( .A(KEYINPUT100), .B(n707), .ZN(n708) );
  NAND2_X1 U807 ( .A1(n708), .A2(G8), .ZN(n709) );
  XNOR2_X1 U808 ( .A(KEYINPUT30), .B(n709), .ZN(n710) );
  NOR2_X1 U809 ( .A1(G168), .A2(n710), .ZN(n711) );
  NOR2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U811 ( .A(KEYINPUT31), .B(n713), .Z(n742) );
  INV_X1 U812 ( .A(n752), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n722), .A2(G2072), .ZN(n714) );
  XNOR2_X1 U814 ( .A(n714), .B(KEYINPUT27), .ZN(n716) );
  XOR2_X1 U815 ( .A(G1956), .B(KEYINPUT96), .Z(n991) );
  NOR2_X1 U816 ( .A1(n722), .A2(n991), .ZN(n715) );
  NOR2_X1 U817 ( .A1(n716), .A2(n715), .ZN(n731) );
  NOR2_X1 U818 ( .A1(n920), .A2(n731), .ZN(n717) );
  XOR2_X1 U819 ( .A(n717), .B(KEYINPUT28), .Z(n735) );
  NAND2_X1 U820 ( .A1(n752), .A2(G1348), .ZN(n720) );
  INV_X1 U821 ( .A(n752), .ZN(n718) );
  NAND2_X1 U822 ( .A1(n718), .A2(G2067), .ZN(n719) );
  NAND2_X1 U823 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U824 ( .A(KEYINPUT98), .B(n721), .Z(n728) );
  XOR2_X1 U825 ( .A(G1996), .B(KEYINPUT97), .Z(n934) );
  NAND2_X1 U826 ( .A1(n722), .A2(n934), .ZN(n723) );
  XNOR2_X1 U827 ( .A(KEYINPUT26), .B(n723), .ZN(n724) );
  NAND2_X1 U828 ( .A1(n724), .A2(n513), .ZN(n725) );
  NOR2_X1 U829 ( .A1(n921), .A2(n725), .ZN(n726) );
  NAND2_X1 U830 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U831 ( .A1(n728), .A2(n902), .ZN(n729) );
  AND2_X1 U832 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U833 ( .A1(n920), .A2(n731), .ZN(n732) );
  NAND2_X1 U834 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U835 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U836 ( .A(n736), .B(KEYINPUT29), .ZN(n739) );
  AND2_X1 U837 ( .A1(G171), .A2(n737), .ZN(n738) );
  NOR2_X1 U838 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U839 ( .A(n740), .B(KEYINPUT99), .ZN(n741) );
  NAND2_X1 U840 ( .A1(n742), .A2(n741), .ZN(n751) );
  INV_X1 U841 ( .A(n751), .ZN(n743) );
  NOR2_X1 U842 ( .A1(n744), .A2(n743), .ZN(n746) );
  XNOR2_X1 U843 ( .A(n746), .B(n745), .ZN(n750) );
  NAND2_X1 U844 ( .A1(G8), .A2(n747), .ZN(n748) );
  XOR2_X1 U845 ( .A(KEYINPUT93), .B(n748), .Z(n749) );
  NAND2_X1 U846 ( .A1(n750), .A2(n749), .ZN(n761) );
  NAND2_X1 U847 ( .A1(G286), .A2(n751), .ZN(n757) );
  NOR2_X1 U848 ( .A1(G1971), .A2(n781), .ZN(n754) );
  NOR2_X1 U849 ( .A1(G2090), .A2(n752), .ZN(n753) );
  NOR2_X1 U850 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U851 ( .A1(n755), .A2(G303), .ZN(n756) );
  NAND2_X1 U852 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U853 ( .A1(n758), .A2(G8), .ZN(n759) );
  XNOR2_X1 U854 ( .A(n759), .B(KEYINPUT32), .ZN(n760) );
  NAND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n776) );
  NOR2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n908) );
  NOR2_X1 U857 ( .A1(G1971), .A2(G303), .ZN(n762) );
  NOR2_X1 U858 ( .A1(n908), .A2(n762), .ZN(n764) );
  INV_X1 U859 ( .A(KEYINPUT33), .ZN(n763) );
  AND2_X1 U860 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U861 ( .A1(n776), .A2(n765), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n910) );
  INV_X1 U863 ( .A(n910), .ZN(n766) );
  NOR2_X1 U864 ( .A1(n781), .A2(n766), .ZN(n767) );
  NOR2_X1 U865 ( .A1(KEYINPUT33), .A2(n767), .ZN(n770) );
  NAND2_X1 U866 ( .A1(n908), .A2(KEYINPUT33), .ZN(n768) );
  NOR2_X1 U867 ( .A1(n768), .A2(n781), .ZN(n769) );
  NOR2_X1 U868 ( .A1(n770), .A2(n769), .ZN(n771) );
  AND2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U870 ( .A(G1981), .B(G305), .Z(n904) );
  NAND2_X1 U871 ( .A1(n773), .A2(n904), .ZN(n785) );
  NOR2_X1 U872 ( .A1(G2090), .A2(G303), .ZN(n774) );
  NAND2_X1 U873 ( .A1(G8), .A2(n774), .ZN(n775) );
  NAND2_X1 U874 ( .A1(n776), .A2(n775), .ZN(n777) );
  AND2_X1 U875 ( .A1(n777), .A2(n781), .ZN(n783) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XOR2_X1 U877 ( .A(n778), .B(KEYINPUT92), .Z(n779) );
  XNOR2_X1 U878 ( .A(KEYINPUT24), .B(n779), .ZN(n780) );
  NOR2_X1 U879 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U880 ( .A1(n783), .A2(n782), .ZN(n784) );
  AND2_X1 U881 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U882 ( .A(n786), .B(KEYINPUT102), .ZN(n787) );
  NOR2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n790) );
  XNOR2_X1 U884 ( .A(G1986), .B(G290), .ZN(n919) );
  NAND2_X1 U885 ( .A1(n919), .A2(n803), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n806) );
  INV_X1 U887 ( .A(n791), .ZN(n794) );
  NOR2_X1 U888 ( .A1(G1986), .A2(G290), .ZN(n792) );
  NOR2_X1 U889 ( .A1(G1991), .A2(n848), .ZN(n954) );
  NOR2_X1 U890 ( .A1(n792), .A2(n954), .ZN(n793) );
  NOR2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n796) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n857), .ZN(n795) );
  XOR2_X1 U893 ( .A(KEYINPUT103), .B(n795), .Z(n958) );
  NOR2_X1 U894 ( .A1(n796), .A2(n958), .ZN(n797) );
  XNOR2_X1 U895 ( .A(n797), .B(KEYINPUT39), .ZN(n798) );
  XNOR2_X1 U896 ( .A(n798), .B(KEYINPUT104), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n801), .A2(n852), .ZN(n973) );
  NAND2_X1 U899 ( .A1(n802), .A2(n973), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U902 ( .A(KEYINPUT40), .B(n807), .ZN(G329) );
  XOR2_X1 U903 ( .A(G2438), .B(KEYINPUT106), .Z(n809) );
  XNOR2_X1 U904 ( .A(G2454), .B(G2435), .ZN(n808) );
  XNOR2_X1 U905 ( .A(n809), .B(n808), .ZN(n810) );
  XOR2_X1 U906 ( .A(n810), .B(G2430), .Z(n812) );
  XNOR2_X1 U907 ( .A(G1341), .B(G1348), .ZN(n811) );
  XNOR2_X1 U908 ( .A(n812), .B(n811), .ZN(n816) );
  XOR2_X1 U909 ( .A(G2427), .B(KEYINPUT107), .Z(n814) );
  XNOR2_X1 U910 ( .A(G2443), .B(G2446), .ZN(n813) );
  XNOR2_X1 U911 ( .A(n814), .B(n813), .ZN(n815) );
  XOR2_X1 U912 ( .A(n816), .B(n815), .Z(n818) );
  XNOR2_X1 U913 ( .A(KEYINPUT105), .B(G2451), .ZN(n817) );
  XNOR2_X1 U914 ( .A(n818), .B(n817), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n819), .A2(G14), .ZN(n897) );
  XOR2_X1 U916 ( .A(KEYINPUT108), .B(n897), .Z(G401) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U919 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n822) );
  XOR2_X1 U921 ( .A(KEYINPUT109), .B(n822), .Z(n823) );
  NAND2_X1 U922 ( .A1(n824), .A2(n823), .ZN(G188) );
  XNOR2_X1 U923 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  INV_X1 U929 ( .A(n827), .ZN(G319) );
  XNOR2_X1 U930 ( .A(n921), .B(n828), .ZN(n830) );
  XNOR2_X1 U931 ( .A(G171), .B(n902), .ZN(n829) );
  XNOR2_X1 U932 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U933 ( .A(n831), .B(G286), .Z(n832) );
  NOR2_X1 U934 ( .A1(G37), .A2(n832), .ZN(G397) );
  NAND2_X1 U935 ( .A1(G136), .A2(n860), .ZN(n834) );
  NAND2_X1 U936 ( .A1(G100), .A2(n512), .ZN(n833) );
  NAND2_X1 U937 ( .A1(n834), .A2(n833), .ZN(n839) );
  NAND2_X1 U938 ( .A1(G124), .A2(n864), .ZN(n835) );
  XNOR2_X1 U939 ( .A(n835), .B(KEYINPUT44), .ZN(n837) );
  NAND2_X1 U940 ( .A1(n866), .A2(G112), .ZN(n836) );
  NAND2_X1 U941 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U942 ( .A1(n839), .A2(n838), .ZN(G162) );
  NAND2_X1 U943 ( .A1(G142), .A2(n860), .ZN(n841) );
  NAND2_X1 U944 ( .A1(G106), .A2(n512), .ZN(n840) );
  NAND2_X1 U945 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n842), .B(KEYINPUT45), .ZN(n844) );
  NAND2_X1 U947 ( .A1(G130), .A2(n864), .ZN(n843) );
  NAND2_X1 U948 ( .A1(n844), .A2(n843), .ZN(n847) );
  NAND2_X1 U949 ( .A1(G118), .A2(n866), .ZN(n845) );
  XNOR2_X1 U950 ( .A(KEYINPUT113), .B(n845), .ZN(n846) );
  NOR2_X1 U951 ( .A1(n847), .A2(n846), .ZN(n856) );
  XNOR2_X1 U952 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n848), .B(KEYINPUT46), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n854) );
  XNOR2_X1 U956 ( .A(G164), .B(G160), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n857), .B(G162), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n873) );
  NAND2_X1 U961 ( .A1(G139), .A2(n860), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G103), .A2(n512), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n871) );
  NAND2_X1 U964 ( .A1(n864), .A2(G127), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT114), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G115), .A2(n866), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n967) );
  XNOR2_X1 U970 ( .A(n956), .B(n967), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n874) );
  NOR2_X1 U972 ( .A1(G37), .A2(n874), .ZN(G395) );
  XNOR2_X1 U973 ( .A(G1991), .B(KEYINPUT41), .ZN(n884) );
  XOR2_X1 U974 ( .A(G1976), .B(G1971), .Z(n876) );
  XNOR2_X1 U975 ( .A(G1996), .B(G1986), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n880) );
  XOR2_X1 U977 ( .A(G1981), .B(G1956), .Z(n878) );
  XNOR2_X1 U978 ( .A(G1966), .B(G1961), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U980 ( .A(n880), .B(n879), .Z(n882) );
  XNOR2_X1 U981 ( .A(KEYINPUT112), .B(G2474), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(G229) );
  XOR2_X1 U984 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n886) );
  XNOR2_X1 U985 ( .A(KEYINPUT110), .B(G2678), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U987 ( .A(KEYINPUT42), .B(G2090), .Z(n888) );
  XNOR2_X1 U988 ( .A(G2067), .B(G2072), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(n890), .B(n889), .Z(n892) );
  XNOR2_X1 U991 ( .A(G2096), .B(G2100), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n894) );
  XOR2_X1 U993 ( .A(G2084), .B(G2078), .Z(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(G227) );
  NOR2_X1 U995 ( .A1(G397), .A2(G395), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n895), .B(KEYINPUT116), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G229), .A2(G227), .ZN(n898) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n898), .ZN(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n901), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1004 ( .A(KEYINPUT56), .B(G16), .Z(n929) );
  XNOR2_X1 U1005 ( .A(n902), .B(G1348), .ZN(n903) );
  XNOR2_X1 U1006 ( .A(n903), .B(KEYINPUT123), .ZN(n927) );
  XNOR2_X1 U1007 ( .A(G1966), .B(G168), .ZN(n905) );
  NAND2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1009 ( .A(n906), .B(KEYINPUT57), .ZN(n907) );
  XNOR2_X1 U1010 ( .A(KEYINPUT122), .B(n907), .ZN(n917) );
  INV_X1 U1011 ( .A(n908), .ZN(n909) );
  NAND2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1013 ( .A(n911), .B(KEYINPUT124), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(G166), .B(G1971), .ZN(n913) );
  XNOR2_X1 U1015 ( .A(G171), .B(G1961), .ZN(n912) );
  NAND2_X1 U1016 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n925) );
  XOR2_X1 U1020 ( .A(n920), .B(G1956), .Z(n923) );
  XNOR2_X1 U1021 ( .A(n921), .B(G1341), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n952) );
  XOR2_X1 U1026 ( .A(G2072), .B(G33), .Z(n930) );
  NAND2_X1 U1027 ( .A1(n930), .A2(G28), .ZN(n940) );
  XNOR2_X1 U1028 ( .A(G2067), .B(G26), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(G1991), .B(G25), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(n933), .B(G27), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G32), .B(n934), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT53), .B(n941), .Z(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT54), .B(G34), .Z(n942) );
  XNOR2_X1 U1038 ( .A(G2084), .B(n942), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G35), .B(G2090), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n947), .B(KEYINPUT55), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G29), .B(KEYINPUT121), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(G11), .A2(n950), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n981) );
  XOR2_X1 U1047 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n976) );
  XOR2_X1 U1048 ( .A(G160), .B(G2084), .Z(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n961) );
  XOR2_X1 U1051 ( .A(G2090), .B(G162), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT51), .B(n959), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1057 ( .A(KEYINPUT118), .B(n966), .Z(n972) );
  XOR2_X1 U1058 ( .A(G2072), .B(n967), .Z(n969) );
  XOR2_X1 U1059 ( .A(G164), .B(G2078), .Z(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1061 ( .A(KEYINPUT50), .B(n970), .Z(n971) );
  NOR2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(n976), .B(n975), .ZN(n977) );
  NOR2_X1 U1065 ( .A1(KEYINPUT55), .A2(n977), .ZN(n978) );
  XOR2_X1 U1066 ( .A(KEYINPUT120), .B(n978), .Z(n979) );
  NAND2_X1 U1067 ( .A1(G29), .A2(n979), .ZN(n980) );
  NAND2_X1 U1068 ( .A1(n981), .A2(n980), .ZN(n1009) );
  XNOR2_X1 U1069 ( .A(n982), .B(G5), .ZN(n1002) );
  XNOR2_X1 U1070 ( .A(G1986), .B(G24), .ZN(n987) );
  XNOR2_X1 U1071 ( .A(G1971), .B(G22), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1976), .B(G23), .ZN(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(KEYINPUT127), .B(n985), .ZN(n986) );
  NOR2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1076 ( .A(KEYINPUT58), .B(n988), .Z(n1000) );
  XNOR2_X1 U1077 ( .A(KEYINPUT59), .B(G1348), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n989), .B(G4), .ZN(n995) );
  XOR2_X1 U1079 ( .A(G1981), .B(KEYINPUT125), .Z(n990) );
  XNOR2_X1 U1080 ( .A(G6), .B(n990), .ZN(n993) );
  XOR2_X1 U1081 ( .A(n991), .B(G20), .Z(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(G19), .B(G1341), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1086 ( .A(KEYINPUT60), .B(n998), .Z(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(KEYINPUT126), .B(G1966), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G21), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(KEYINPUT61), .B(n1006), .Z(n1007) );
  NOR2_X1 U1093 ( .A1(G16), .A2(n1007), .ZN(n1008) );
  NOR2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(n1010), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1096 ( .A(G311), .ZN(G150) );
endmodule

