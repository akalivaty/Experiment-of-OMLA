//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n646, new_n647, new_n648, new_n649, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT69), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n466), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n461), .B2(new_n462), .ZN(new_n491));
  AND2_X1   g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n466), .A2(G138), .A3(new_n479), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n466), .A2(KEYINPUT4), .A3(G138), .ZN(new_n497));
  NAND2_X1  g072(.A1(G102), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(G2105), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n503), .A2(KEYINPUT70), .A3(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  XOR2_X1   g086(.A(new_n511), .B(KEYINPUT71), .Z(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n509), .A2(G88), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n506), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n514), .A2(new_n515), .A3(new_n517), .A4(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n518), .B1(new_n510), .B2(new_n512), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n517), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT72), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n528), .ZN(G166));
  NAND4_X1  g104(.A1(new_n519), .A2(new_n521), .A3(G51), .A4(G543), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n507), .A2(new_n508), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n536));
  AND2_X1   g111(.A1(KEYINPUT73), .A2(G89), .ZN(new_n537));
  NOR2_X1   g112(.A1(KEYINPUT73), .A2(G89), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n535), .A2(new_n536), .A3(new_n516), .A4(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n535), .A2(G63), .A3(new_n536), .ZN(new_n542));
  NAND3_X1  g117(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n541), .A2(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND3_X1  g122(.A1(new_n535), .A2(G64), .A3(new_n536), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT74), .B(G90), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n535), .A2(new_n536), .A3(new_n516), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n516), .A2(G52), .A3(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n551), .A2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  NAND2_X1  g133(.A1(new_n509), .A2(G56), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n518), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT75), .B(G81), .Z(new_n562));
  NAND3_X1  g137(.A1(new_n509), .A2(new_n516), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n516), .A2(G43), .A3(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND3_X1  g146(.A1(new_n523), .A2(KEYINPUT9), .A3(G53), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n516), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n509), .A2(G91), .A3(new_n516), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  NOR3_X1   g156(.A1(new_n580), .A2(new_n581), .A3(new_n518), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n535), .A2(G65), .A3(new_n536), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT76), .B1(new_n585), .B2(G651), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n579), .B1(new_n582), .B2(new_n586), .ZN(G299));
  AND2_X1   g162(.A1(new_n525), .A2(new_n528), .ZN(G303));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g164(.A1(G49), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n522), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n516), .A2(KEYINPUT77), .A3(G49), .A4(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n509), .A2(G87), .A3(new_n516), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G288));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n518), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n535), .A2(G61), .A3(new_n536), .ZN(new_n600));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n602), .A2(KEYINPUT78), .A3(G651), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n509), .A2(G86), .A3(new_n516), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n599), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n599), .A2(new_n603), .A3(KEYINPUT79), .A4(new_n606), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(G305));
  NAND2_X1  g186(.A1(new_n523), .A2(G47), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n509), .A2(G85), .A3(new_n516), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G72), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n509), .B2(G60), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n619));
  OAI21_X1  g194(.A(G651), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI211_X1 g195(.A(KEYINPUT80), .B(new_n617), .C1(new_n509), .C2(G60), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n620), .A2(KEYINPUT81), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n503), .A2(KEYINPUT70), .A3(G543), .ZN(new_n624));
  AOI21_X1  g199(.A(KEYINPUT70), .B1(new_n503), .B2(G543), .ZN(new_n625));
  OAI211_X1 g200(.A(G60), .B(new_n536), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n616), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n518), .B1(new_n627), .B2(KEYINPUT80), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n618), .A2(new_n619), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n615), .B1(new_n622), .B2(new_n630), .ZN(G290));
  NAND2_X1  g206(.A1(G301), .A2(G868), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n509), .A2(G92), .A3(new_n516), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT10), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n509), .A2(KEYINPUT10), .A3(G92), .A4(new_n516), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n516), .A2(G54), .A3(G543), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n535), .A2(G66), .A3(new_n536), .ZN(new_n639));
  NAND2_X1  g214(.A1(G79), .A2(G543), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n641), .B2(G651), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n632), .B1(new_n643), .B2(G868), .ZN(G284));
  OAI21_X1  g219(.A(new_n632), .B1(new_n643), .B2(G868), .ZN(G321));
  NAND2_X1  g220(.A1(G286), .A2(G868), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n581), .B1(new_n580), .B2(new_n518), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n585), .A2(KEYINPUT76), .A3(G651), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n578), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n646), .B1(new_n649), .B2(G868), .ZN(G297));
  OAI21_X1  g225(.A(new_n646), .B1(new_n649), .B2(G868), .ZN(G280));
  INV_X1    g226(.A(G559), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n643), .B1(new_n652), .B2(G860), .ZN(G148));
  NOR2_X1   g228(.A1(new_n566), .A2(G868), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n643), .A2(KEYINPUT82), .A3(new_n652), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n637), .A2(new_n642), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n656), .B1(new_n657), .B2(G559), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n654), .B1(new_n659), .B2(G868), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g236(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g237(.A1(new_n481), .A2(G2104), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT12), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT13), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n481), .A2(G135), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT85), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n484), .A2(G123), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n479), .A2(KEYINPUT86), .A3(G111), .ZN(new_n671));
  OAI21_X1  g246(.A(KEYINPUT86), .B1(new_n479), .B2(G111), .ZN(new_n672));
  OR2_X1    g247(.A1(G99), .A2(G2105), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(G2104), .A3(new_n673), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n669), .B(new_n670), .C1(new_n671), .C2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n667), .B(new_n677), .C1(G2100), .C2(new_n665), .ZN(G156));
  XNOR2_X1  g253(.A(G2427), .B(G2438), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2430), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT15), .B(G2435), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(KEYINPUT14), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  XOR2_X1   g260(.A(G1341), .B(G1348), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2451), .B(G2454), .Z(new_n690));
  XNOR2_X1  g265(.A(G2443), .B(G2446), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(G14), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G401));
  XOR2_X1   g271(.A(G2084), .B(G2090), .Z(new_n697));
  XNOR2_X1  g272(.A(G2067), .B(G2678), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n697), .ZN(new_n700));
  XOR2_X1   g275(.A(G2072), .B(G2078), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(KEYINPUT89), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(KEYINPUT17), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n697), .B2(new_n698), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n703), .A2(KEYINPUT17), .ZN(new_n706));
  OAI221_X1 g281(.A(new_n699), .B1(new_n698), .B2(new_n702), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n699), .A2(new_n701), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT18), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(new_n676), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G2100), .ZN(G227));
  XNOR2_X1  g287(.A(G1971), .B(G1976), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT19), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(G1961), .B(G1966), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1956), .B(G2474), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT20), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n717), .A2(new_n719), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n721), .B(new_n724), .C1(new_n714), .C2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT91), .B(G1986), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(G1991), .B(G1996), .ZN(new_n730));
  INV_X1    g305(.A(G1981), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n729), .B(new_n732), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(G229));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G32), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n484), .A2(G129), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT97), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n479), .A2(G105), .A3(G2104), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT26), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n739), .B(new_n741), .C1(new_n481), .C2(G141), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n736), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT98), .Z(new_n746));
  XOR2_X1   g321(.A(KEYINPUT27), .B(G1996), .Z(new_n747));
  AND2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n675), .A2(new_n735), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(G28), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n735), .B1(new_n751), .B2(G28), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  NOR2_X1   g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G16), .ZN(new_n758));
  NOR2_X1   g333(.A1(G168), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(G21), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n748), .A2(new_n749), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G27), .A2(G29), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G164), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2078), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n735), .A2(G33), .ZN(new_n768));
  NAND2_X1  g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  INV_X1    g344(.A(G127), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n463), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n479), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n775));
  NAND2_X1  g350(.A1(G103), .A2(G2104), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G2105), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n479), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n481), .A2(G139), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n768), .B1(new_n780), .B2(new_n735), .ZN(new_n781));
  INV_X1    g356(.A(G2084), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n735), .B1(KEYINPUT24), .B2(G34), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(KEYINPUT24), .B2(G34), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n477), .B2(G29), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n781), .A2(G2072), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n767), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n758), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n758), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(G1961), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(G1961), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n781), .B2(G2072), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n787), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n760), .A2(new_n761), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n785), .A2(new_n782), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT96), .Z(new_n797));
  NAND4_X1  g372(.A1(new_n763), .A2(new_n793), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n481), .A2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n484), .A2(G119), .ZN(new_n801));
  NOR2_X1   g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(new_n479), .B2(G107), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G25), .B(new_n804), .S(G29), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT92), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G1991), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G16), .A2(G24), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT81), .B1(new_n620), .B2(new_n621), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n628), .A2(new_n623), .A3(new_n629), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n614), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n809), .B1(new_n812), .B2(G16), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n813), .A2(G1986), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(G1986), .ZN(new_n815));
  OR3_X1    g390(.A1(new_n808), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G6), .B(G305), .S(G16), .Z(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G22), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G166), .B2(G16), .ZN(new_n821));
  INV_X1    g396(.A(G1971), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G16), .A2(G23), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT93), .Z(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G288), .B2(new_n758), .ZN(new_n826));
  INV_X1    g401(.A(G1976), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n819), .A2(new_n823), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n816), .B1(KEYINPUT34), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n832), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n735), .A2(G35), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G162), .B2(new_n735), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT101), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT29), .ZN(new_n842));
  INV_X1    g417(.A(G2090), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n758), .A2(G20), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n649), .B2(new_n758), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G1956), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n758), .A2(G19), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n566), .B2(new_n758), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(G1341), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n481), .A2(G140), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n484), .A2(G128), .ZN(new_n856));
  NOR2_X1   g431(.A1(G104), .A2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(new_n479), .B2(G116), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G29), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n735), .A2(G26), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT28), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G2067), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n758), .A2(G4), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n643), .B2(new_n758), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G1348), .ZN(new_n869));
  AOI211_X1 g444(.A(new_n866), .B(new_n869), .C1(new_n842), .C2(new_n843), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n850), .A2(KEYINPUT103), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n851), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n799), .A2(new_n838), .A3(new_n872), .ZN(G150));
  INV_X1    g448(.A(G150), .ZN(G311));
  NAND2_X1  g449(.A1(new_n559), .A2(new_n560), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G651), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n563), .A2(new_n564), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n535), .A2(G67), .A3(new_n536), .ZN(new_n878));
  NAND2_X1  g453(.A1(G80), .A2(G543), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(G651), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n535), .A2(G93), .A3(new_n536), .A4(new_n516), .ZN(new_n882));
  XOR2_X1   g457(.A(KEYINPUT104), .B(G55), .Z(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(G543), .A3(new_n516), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n876), .A2(new_n877), .A3(new_n881), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n518), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  OAI22_X1  g463(.A1(new_n561), .A2(new_n565), .B1(new_n888), .B2(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT38), .Z(new_n891));
  NOR2_X1   g466(.A1(new_n657), .A2(new_n652), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n894));
  AOI21_X1  g469(.A(G860), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n881), .A2(new_n886), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G860), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT37), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT105), .Z(G145));
  XNOR2_X1  g476(.A(new_n501), .B(new_n859), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n780), .ZN(new_n903));
  AOI22_X1  g478(.A1(G130), .A2(new_n484), .B1(new_n481), .B2(G142), .ZN(new_n904));
  OAI21_X1  g479(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  INV_X1    g481(.A(G118), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n905), .A2(new_n906), .B1(new_n907), .B2(G2105), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n906), .B2(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n664), .B(new_n910), .Z(new_n911));
  XNOR2_X1  g486(.A(new_n903), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n743), .B(new_n804), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n675), .B(new_n477), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(new_n488), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n916), .B2(new_n914), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g494(.A(new_n659), .B(new_n890), .ZN(new_n920));
  NAND2_X1  g495(.A1(G299), .A2(new_n643), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n649), .A2(new_n657), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NOR2_X1   g501(.A1(G299), .A2(new_n643), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n649), .A2(new_n657), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n922), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n920), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g511(.A1(G305), .A2(G166), .ZN(new_n937));
  NAND3_X1  g512(.A1(G303), .A2(new_n609), .A3(new_n610), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G288), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n812), .A2(new_n941), .ZN(new_n942));
  AOI211_X1 g517(.A(G288), .B(new_n614), .C1(new_n810), .C2(new_n811), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT108), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  NAND2_X1  g520(.A1(G290), .A2(G288), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n812), .A2(new_n941), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n940), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT108), .B1(new_n942), .B2(new_n943), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n939), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n925), .A2(new_n953), .A3(new_n933), .A4(new_n934), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n936), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n936), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n897), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(G868), .B2(new_n958), .ZN(G295));
  OAI21_X1  g534(.A(new_n957), .B1(G868), .B2(new_n958), .ZN(G331));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n518), .B1(new_n548), .B2(new_n549), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n541), .B(new_n545), .C1(new_n962), .C2(new_n555), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n518), .B1(new_n542), .B2(new_n543), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n534), .A2(new_n540), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n551), .B(new_n556), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  AND4_X1   g541(.A1(new_n889), .A2(new_n887), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n963), .A2(new_n966), .B1(new_n887), .B2(new_n889), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n922), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT41), .B1(new_n921), .B2(new_n922), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n963), .A2(new_n966), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n890), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n887), .A2(new_n963), .A3(new_n966), .A4(new_n889), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n974), .A2(new_n975), .B1(new_n921), .B2(new_n922), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n949), .A2(new_n978), .A3(new_n951), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n931), .B2(new_n969), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n946), .A2(new_n945), .A3(new_n947), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n939), .B1(new_n950), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n946), .A2(new_n947), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n983), .A2(KEYINPUT108), .B1(new_n937), .B2(new_n938), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G37), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n979), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n929), .A2(KEYINPUT110), .A3(new_n930), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n969), .B1(new_n929), .B2(KEYINPUT110), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n977), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(new_n949), .A3(new_n951), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n996), .A3(new_n986), .A4(new_n985), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n990), .A2(new_n991), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n987), .A2(new_n996), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n995), .A2(KEYINPUT43), .A3(new_n986), .A4(new_n985), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n961), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g580(.A(KEYINPUT111), .B(new_n1003), .C1(new_n998), .C2(new_n999), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(G397));
  XNOR2_X1  g582(.A(new_n859), .B(G2067), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(G1996), .B2(new_n743), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n472), .A2(G40), .A3(new_n476), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  INV_X1    g586(.A(new_n495), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(KEYINPUT4), .B2(new_n493), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1013), .B2(new_n499), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1009), .A2(new_n1010), .A3(new_n1016), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1016), .A2(G1996), .A3(new_n1010), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT113), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1019), .B2(new_n744), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1016), .A2(new_n1010), .ZN(new_n1021));
  INV_X1    g596(.A(new_n807), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n804), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n804), .A2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1021), .A2(G1986), .A3(G290), .ZN(new_n1027));
  INV_X1    g602(.A(G1986), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1021), .A2(new_n1028), .A3(new_n812), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(G8), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1034));
  INV_X1    g609(.A(G40), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1035), .B(new_n475), .C1(new_n471), .C2(G2105), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1384), .B1(new_n496), .B2(new_n500), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(G8), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1034), .A2(new_n1040), .B1(G1976), .B2(new_n941), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT116), .B(G86), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n509), .A2(new_n516), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n605), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT117), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1049), .A3(new_n605), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(new_n599), .A3(new_n603), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G1981), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n599), .A2(new_n603), .A3(new_n731), .A4(new_n606), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1044), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1052), .A2(KEYINPUT118), .A3(KEYINPUT49), .A4(new_n1053), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n941), .A2(G1976), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT52), .B1(G288), .B2(new_n827), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1043), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1036), .B1(new_n1037), .B2(KEYINPUT45), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1037), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1036), .A3(new_n1070), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n1067), .A2(G1971), .B1(new_n1071), .B2(G2090), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n525), .A2(G8), .A3(new_n528), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1072), .A2(G8), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1053), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G288), .A2(G1976), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1060), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1057), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1064), .A2(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1956), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1071), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1037), .A2(KEYINPUT45), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(new_n1016), .A3(new_n1036), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n572), .A2(new_n576), .A3(KEYINPUT122), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n649), .B(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1084), .A2(new_n1092), .A3(new_n1087), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1036), .B1(new_n1037), .B2(new_n1068), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n864), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n657), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1095), .B1(new_n1102), .B2(KEYINPUT123), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1071), .A2(new_n1096), .B1(new_n864), .B2(new_n1100), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n657), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1094), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n643), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1095), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1084), .A2(KEYINPUT61), .A3(new_n1092), .A4(new_n1087), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1085), .A2(new_n1036), .A3(new_n1016), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1115), .A2(G1996), .B1(new_n1100), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n566), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1120), .A3(new_n566), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n657), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1104), .A2(KEYINPUT60), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1119), .A2(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1107), .B1(new_n1114), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1063), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1060), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1043), .A2(new_n1060), .A3(KEYINPUT119), .A4(new_n1063), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1075), .B1(new_n1072), .B2(G8), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1076), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1125), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n761), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1069), .A2(new_n1070), .A3(new_n782), .A4(new_n1036), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1140));
  OAI21_X1  g715(.A(G168), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1135), .B1(new_n1141), .B2(G8), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT124), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1145));
  INV_X1    g720(.A(G8), .ZN(new_n1146));
  NOR2_X1   g721(.A1(G168), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1135), .B(G8), .C1(new_n1143), .C2(G286), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1142), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT53), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1085), .A2(new_n1016), .A3(new_n766), .A4(new_n1036), .ZN(new_n1154));
  INV_X1    g729(.A(G1961), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1153), .A2(new_n1154), .B1(new_n1071), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1067), .A2(KEYINPUT53), .A3(new_n766), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(G301), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(G301), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1152), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1160), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(KEYINPUT54), .A3(new_n1158), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1151), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1082), .B1(new_n1134), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT62), .B1(new_n1142), .B2(new_n1150), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT125), .ZN(new_n1168));
  OR3_X1    g743(.A1(new_n1142), .A2(KEYINPUT62), .A3(new_n1150), .ZN(new_n1169));
  AND4_X1   g744(.A1(new_n1130), .A2(new_n1129), .A3(new_n1132), .A4(new_n1160), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1171), .B(KEYINPUT62), .C1(new_n1142), .C2(new_n1150), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g749(.A(new_n1146), .B(G286), .C1(new_n1136), .C2(new_n1138), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .A4(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1177));
  AND3_X1   g752(.A1(new_n1176), .A2(KEYINPUT121), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT121), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1132), .A2(KEYINPUT63), .A3(new_n1175), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1064), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1032), .B1(new_n1174), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1021), .B1(new_n743), .B2(new_n1008), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1019), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1019), .A2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1184), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT47), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1188), .B(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n859), .A2(G2067), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1021), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1029), .B(KEYINPUT127), .Z(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT48), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1196), .B1(new_n1198), .B2(new_n1026), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1192), .A2(new_n1193), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1183), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g776(.A1(G227), .A2(new_n457), .ZN(new_n1203));
  AND3_X1   g777(.A1(new_n733), .A2(new_n695), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n1204), .A2(new_n918), .A3(new_n998), .ZN(G225));
  INV_X1    g779(.A(G225), .ZN(G308));
endmodule


