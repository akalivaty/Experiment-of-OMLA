

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XNOR2_X1 U324 ( .A(n343), .B(n342), .ZN(n351) );
  XNOR2_X1 U325 ( .A(n341), .B(G29GAT), .ZN(n342) );
  XNOR2_X1 U326 ( .A(n479), .B(KEYINPUT104), .ZN(n480) );
  XNOR2_X1 U327 ( .A(n357), .B(n356), .ZN(n575) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U329 ( .A(G43GAT), .B(G50GAT), .Z(n293) );
  NOR2_X1 U330 ( .A1(n581), .A2(n383), .ZN(n384) );
  XNOR2_X1 U331 ( .A(n367), .B(n292), .ZN(n370) );
  XNOR2_X1 U332 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U333 ( .A(n370), .B(n369), .ZN(n375) );
  XNOR2_X1 U334 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U335 ( .A(n481), .B(n480), .ZN(n525) );
  NAND2_X1 U336 ( .A1(n451), .A2(n464), .ZN(n570) );
  XNOR2_X1 U337 ( .A(n377), .B(n376), .ZN(n569) );
  INV_X1 U338 ( .A(G43GAT), .ZN(n484) );
  XNOR2_X1 U339 ( .A(KEYINPUT90), .B(n472), .ZN(n527) );
  XNOR2_X1 U340 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n453) );
  XNOR2_X1 U341 ( .A(n484), .B(KEYINPUT40), .ZN(n485) );
  XNOR2_X1 U342 ( .A(n454), .B(n453), .ZN(G1350GAT) );
  XNOR2_X1 U343 ( .A(n486), .B(n485), .ZN(G1330GAT) );
  XNOR2_X1 U344 ( .A(G22GAT), .B(G15GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n294), .B(KEYINPUT74), .ZN(n340) );
  XOR2_X1 U346 ( .A(G64GAT), .B(G78GAT), .Z(n296) );
  XNOR2_X1 U347 ( .A(KEYINPUT81), .B(KEYINPUT83), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n340), .B(n297), .ZN(n312) );
  XNOR2_X1 U350 ( .A(G155GAT), .B(G127GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n298), .B(G1GAT), .ZN(n391) );
  XOR2_X1 U352 ( .A(KEYINPUT82), .B(n391), .Z(n300) );
  NAND2_X1 U353 ( .A1(G231GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U355 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n302) );
  XNOR2_X1 U356 ( .A(KEYINPUT15), .B(KEYINPUT84), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U358 ( .A(n304), .B(n303), .Z(n310) );
  XOR2_X1 U359 ( .A(G8GAT), .B(KEYINPUT80), .Z(n306) );
  XNOR2_X1 U360 ( .A(G211GAT), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n325) );
  XOR2_X1 U362 ( .A(KEYINPUT75), .B(KEYINPUT13), .Z(n308) );
  XNOR2_X1 U363 ( .A(G57GAT), .B(G71GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n327) );
  XNOR2_X1 U365 ( .A(n325), .B(n327), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n584) );
  XNOR2_X1 U368 ( .A(n584), .B(KEYINPUT110), .ZN(n547) );
  XOR2_X1 U369 ( .A(G190GAT), .B(G36GAT), .Z(n364) );
  XOR2_X1 U370 ( .A(KEYINPUT91), .B(n364), .Z(n314) );
  NAND2_X1 U371 ( .A1(G226GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n317) );
  XOR2_X1 U373 ( .A(G176GAT), .B(G204GAT), .Z(n316) );
  XNOR2_X1 U374 ( .A(G92GAT), .B(G64GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n326) );
  XOR2_X1 U376 ( .A(n317), .B(n326), .Z(n323) );
  XOR2_X1 U377 ( .A(G197GAT), .B(KEYINPUT87), .Z(n319) );
  XNOR2_X1 U378 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n421) );
  XOR2_X1 U380 ( .A(G169GAT), .B(KEYINPUT19), .Z(n321) );
  XNOR2_X1 U381 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n435) );
  XNOR2_X1 U383 ( .A(n421), .B(n435), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n529) );
  XOR2_X1 U386 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n359) );
  XOR2_X1 U387 ( .A(G148GAT), .B(G120GAT), .Z(n392) );
  XOR2_X1 U388 ( .A(G106GAT), .B(G78GAT), .Z(n427) );
  XNOR2_X1 U389 ( .A(n392), .B(n427), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n327), .B(n326), .ZN(n334) );
  XOR2_X1 U391 ( .A(G85GAT), .B(G99GAT), .Z(n363) );
  XOR2_X1 U392 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n329) );
  XNOR2_X1 U393 ( .A(KEYINPUT76), .B(KEYINPUT31), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U395 ( .A(n363), .B(n330), .Z(n332) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U398 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n581) );
  XNOR2_X1 U400 ( .A(n581), .B(KEYINPUT64), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n337), .B(KEYINPUT41), .ZN(n560) );
  XOR2_X1 U402 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n339) );
  XNOR2_X1 U403 ( .A(KEYINPUT72), .B(KEYINPUT70), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n357) );
  XNOR2_X1 U405 ( .A(n340), .B(G36GAT), .ZN(n343) );
  AND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n341) );
  XOR2_X1 U407 ( .A(G169GAT), .B(G197GAT), .Z(n345) );
  XNOR2_X1 U408 ( .A(G113GAT), .B(G141GAT), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U410 ( .A(KEYINPUT73), .B(KEYINPUT71), .Z(n347) );
  XNOR2_X1 U411 ( .A(G1GAT), .B(G8GAT), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U413 ( .A(n349), .B(n348), .Z(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n352), .B(KEYINPUT30), .ZN(n355) );
  XNOR2_X1 U416 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n293), .B(n353), .ZN(n368) );
  XOR2_X1 U418 ( .A(n368), .B(KEYINPUT29), .Z(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  NOR2_X1 U420 ( .A1(n560), .A2(n575), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  NOR2_X1 U422 ( .A1(n360), .A2(n547), .ZN(n378) );
  XOR2_X1 U423 ( .A(KEYINPUT67), .B(G92GAT), .Z(n362) );
  XNOR2_X1 U424 ( .A(G162GAT), .B(KEYINPUT78), .ZN(n361) );
  XOR2_X1 U425 ( .A(n362), .B(n361), .Z(n377) );
  XOR2_X1 U426 ( .A(G106GAT), .B(G218GAT), .Z(n366) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U429 ( .A(KEYINPUT77), .B(n368), .Z(n369) );
  XOR2_X1 U430 ( .A(G29GAT), .B(G134GAT), .Z(n393) );
  XOR2_X1 U431 ( .A(KEYINPUT11), .B(KEYINPUT79), .Z(n372) );
  XNOR2_X1 U432 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n393), .B(n373), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  NAND2_X1 U436 ( .A1(n378), .A2(n569), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n379), .B(KEYINPUT112), .ZN(n380) );
  XNOR2_X1 U438 ( .A(KEYINPUT47), .B(n380), .ZN(n386) );
  XNOR2_X1 U439 ( .A(KEYINPUT36), .B(n569), .ZN(n588) );
  INV_X1 U440 ( .A(n584), .ZN(n563) );
  NOR2_X1 U441 ( .A1(n588), .A2(n563), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n381), .B(KEYINPUT45), .ZN(n382) );
  NAND2_X1 U443 ( .A1(n382), .A2(n575), .ZN(n383) );
  XOR2_X1 U444 ( .A(KEYINPUT113), .B(n384), .Z(n385) );
  NOR2_X1 U445 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U446 ( .A(KEYINPUT48), .B(n387), .ZN(n535) );
  NOR2_X1 U447 ( .A1(n529), .A2(n535), .ZN(n389) );
  XOR2_X1 U448 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n414) );
  XNOR2_X1 U450 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n390), .B(KEYINPUT85), .ZN(n440) );
  XNOR2_X1 U452 ( .A(n440), .B(n391), .ZN(n413) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U454 ( .A(KEYINPUT89), .B(G85GAT), .Z(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n401) );
  INV_X1 U456 ( .A(n401), .ZN(n399) );
  XOR2_X1 U457 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n397) );
  XNOR2_X1 U458 ( .A(KEYINPUT5), .B(KEYINPUT88), .ZN(n396) );
  XOR2_X1 U459 ( .A(n397), .B(n396), .Z(n400) );
  INV_X1 U460 ( .A(n400), .ZN(n398) );
  NAND2_X1 U461 ( .A1(n399), .A2(n398), .ZN(n403) );
  NAND2_X1 U462 ( .A1(n401), .A2(n400), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n403), .A2(n402), .ZN(n405) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n411) );
  XOR2_X1 U466 ( .A(G141GAT), .B(KEYINPUT2), .Z(n407) );
  XNOR2_X1 U467 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n422) );
  XNOR2_X1 U469 ( .A(n422), .B(KEYINPUT4), .ZN(n409) );
  INV_X1 U470 ( .A(G57GAT), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n472) );
  NAND2_X1 U472 ( .A1(n414), .A2(n527), .ZN(n415) );
  XNOR2_X1 U473 ( .A(KEYINPUT65), .B(n415), .ZN(n574) );
  XOR2_X1 U474 ( .A(G22GAT), .B(G211GAT), .Z(n417) );
  XNOR2_X1 U475 ( .A(G155GAT), .B(G148GAT), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n431) );
  XOR2_X1 U477 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n419) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U480 ( .A(n420), .B(G204GAT), .Z(n424) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n426) );
  INV_X1 U483 ( .A(KEYINPUT22), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n429) );
  XNOR2_X1 U485 ( .A(G50GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U487 ( .A(n431), .B(n430), .Z(n463) );
  NAND2_X1 U488 ( .A1(n574), .A2(n463), .ZN(n433) );
  XNOR2_X1 U489 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n451) );
  XNOR2_X1 U491 ( .A(G134GAT), .B(G190GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n434), .B(G99GAT), .ZN(n439) );
  XOR2_X1 U493 ( .A(n435), .B(G71GAT), .Z(n437) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U496 ( .A(n439), .B(n438), .Z(n442) );
  XNOR2_X1 U497 ( .A(n440), .B(G43GAT), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U499 ( .A(KEYINPUT86), .B(G176GAT), .Z(n444) );
  XNOR2_X1 U500 ( .A(G120GAT), .B(G15GAT), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U502 ( .A(KEYINPUT20), .B(KEYINPUT66), .Z(n446) );
  XNOR2_X1 U503 ( .A(G127GAT), .B(G183GAT), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U505 ( .A(n448), .B(n447), .Z(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n464) );
  INV_X1 U507 ( .A(n570), .ZN(n452) );
  NAND2_X1 U508 ( .A1(n547), .A2(n452), .ZN(n454) );
  XNOR2_X1 U509 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n483) );
  NOR2_X1 U510 ( .A1(n581), .A2(n575), .ZN(n498) );
  XNOR2_X1 U511 ( .A(KEYINPUT27), .B(n529), .ZN(n466) );
  NOR2_X1 U512 ( .A1(n527), .A2(n466), .ZN(n455) );
  XOR2_X1 U513 ( .A(n455), .B(KEYINPUT92), .Z(n536) );
  XNOR2_X1 U514 ( .A(n463), .B(KEYINPUT28), .ZN(n538) );
  INV_X1 U515 ( .A(n464), .ZN(n540) );
  NAND2_X1 U516 ( .A1(n538), .A2(n540), .ZN(n456) );
  NOR2_X1 U517 ( .A1(n536), .A2(n456), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(KEYINPUT93), .ZN(n475) );
  NOR2_X1 U519 ( .A1(n540), .A2(n529), .ZN(n459) );
  INV_X1 U520 ( .A(n463), .ZN(n458) );
  NOR2_X1 U521 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n460), .B(KEYINPUT95), .ZN(n462) );
  INV_X1 U523 ( .A(KEYINPUT25), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n462), .B(n461), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n465), .B(KEYINPUT26), .ZN(n573) );
  INV_X1 U527 ( .A(n466), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n573), .A2(n467), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT94), .ZN(n469) );
  NAND2_X1 U530 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U531 ( .A(KEYINPUT96), .B(n471), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(KEYINPUT97), .ZN(n495) );
  NOR2_X1 U535 ( .A1(n495), .A2(n584), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT103), .ZN(n478) );
  NOR2_X1 U537 ( .A1(n478), .A2(n588), .ZN(n481) );
  INV_X1 U538 ( .A(KEYINPUT37), .ZN(n479) );
  AND2_X1 U539 ( .A1(n498), .A2(n525), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n512) );
  NOR2_X1 U541 ( .A1(n512), .A2(n540), .ZN(n486) );
  NOR2_X1 U542 ( .A1(n575), .A2(n570), .ZN(n488) );
  XNOR2_X1 U543 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n487) );
  XNOR2_X1 U544 ( .A(n488), .B(n487), .ZN(G1348GAT) );
  NOR2_X1 U545 ( .A1(n560), .A2(n570), .ZN(n491) );
  XNOR2_X1 U546 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(G176GAT), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(G1349GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n493) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n500) );
  NAND2_X1 U552 ( .A1(n569), .A2(n584), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT16), .B(n494), .ZN(n496) );
  NOR2_X1 U554 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(KEYINPUT98), .ZN(n515) );
  NAND2_X1 U556 ( .A1(n498), .A2(n515), .ZN(n506) );
  NOR2_X1 U557 ( .A1(n527), .A2(n506), .ZN(n499) );
  XOR2_X1 U558 ( .A(n500), .B(n499), .Z(G1324GAT) );
  NOR2_X1 U559 ( .A1(n529), .A2(n506), .ZN(n502) );
  XNOR2_X1 U560 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1325GAT) );
  NOR2_X1 U562 ( .A1(n540), .A2(n506), .ZN(n504) );
  XNOR2_X1 U563 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(n505), .ZN(G1326GAT) );
  NOR2_X1 U566 ( .A1(n538), .A2(n506), .ZN(n507) );
  XOR2_X1 U567 ( .A(G22GAT), .B(n507), .Z(G1327GAT) );
  NOR2_X1 U568 ( .A1(n512), .A2(n527), .ZN(n509) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  OR2_X1 U571 ( .A1(n512), .A2(n529), .ZN(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT106), .B(n510), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G36GAT), .B(n511), .ZN(G1329GAT) );
  NOR2_X1 U574 ( .A1(n512), .A2(n538), .ZN(n514) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1331GAT) );
  INV_X1 U577 ( .A(n575), .ZN(n541) );
  NOR2_X1 U578 ( .A1(n541), .A2(n560), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n526), .A2(n515), .ZN(n521) );
  NOR2_X1 U580 ( .A1(n527), .A2(n521), .ZN(n517) );
  XNOR2_X1 U581 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G57GAT), .B(n518), .Z(G1332GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n521), .ZN(n519) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n519), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n540), .A2(n521), .ZN(n520) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n538), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U591 ( .A(G78GAT), .B(n524), .Z(G1335GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U593 ( .A1(n527), .A2(n532), .ZN(n528) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n528), .Z(G1336GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n532), .ZN(n530) );
  XOR2_X1 U596 ( .A(G92GAT), .B(n530), .Z(G1337GAT) );
  NOR2_X1 U597 ( .A1(n540), .A2(n532), .ZN(n531) );
  XOR2_X1 U598 ( .A(G99GAT), .B(n531), .Z(G1338GAT) );
  NOR2_X1 U599 ( .A1(n538), .A2(n532), .ZN(n533) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(n533), .Z(n534) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT114), .B(n537), .ZN(n555) );
  NAND2_X1 U604 ( .A1(n538), .A2(n555), .ZN(n539) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n541), .A2(n551), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n545) );
  INV_X1 U609 ( .A(n560), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n551), .A2(n543), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G120GAT), .B(n546), .Z(G1341GAT) );
  NAND2_X1 U613 ( .A1(n547), .A2(n551), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT50), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n553) );
  INV_X1 U617 ( .A(n569), .ZN(n550) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G134GAT), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n573), .A2(n555), .ZN(n565) );
  NOR2_X1 U622 ( .A1(n575), .A2(n565), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n559) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n560), .A2(n565), .ZN(n561) );
  XOR2_X1 U629 ( .A(n562), .B(n561), .Z(G1345GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n565), .ZN(n564) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U632 ( .A1(n569), .A2(n565), .ZN(n566) );
  XOR2_X1 U633 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n568) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(n572), .B(n571), .Z(G1351GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n587) );
  NOR2_X1 U640 ( .A1(n575), .A2(n587), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT59), .B(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U647 ( .A(n587), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

