//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n447, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n602, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(KEYINPUT3), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT67), .B(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(new_n464), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n463), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n468), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n464), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(G2105), .B1(G101), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n474), .A2(G136), .ZN(new_n486));
  INV_X1    g061(.A(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n467), .B2(new_n473), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n487), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n477), .A2(new_n478), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G138), .A4(new_n487), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n477), .A2(KEYINPUT68), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n472), .B2(G2104), .ZN(new_n500));
  AOI211_X1 g075(.A(KEYINPUT68), .B(new_n464), .C1(new_n469), .C2(new_n471), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n487), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(G126), .B(G2105), .C1(new_n500), .C2(new_n501), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n494), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n488), .B2(G126), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n496), .B1(new_n474), .B2(G138), .ZN(new_n512));
  OAI211_X1 g087(.A(KEYINPUT69), .B(new_n511), .C1(new_n512), .C2(new_n498), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(G164));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT70), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n520), .B1(new_n519), .B2(new_n524), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n523), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n516), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n531), .B(new_n533), .C1(new_n536), .C2(KEYINPUT72), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(KEYINPUT72), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n522), .A2(new_n540), .B1(new_n516), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n527), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(G81), .A2(new_n523), .B1(new_n517), .B2(G43), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n527), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G860), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT73), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(new_n517), .A2(G53), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n523), .A2(G91), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n561), .C1(new_n527), .C2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n523), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n517), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT75), .Z(G288));
  AOI22_X1  g145(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n527), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G86), .ZN(new_n574));
  INV_X1    g149(.A(G48), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n522), .A2(new_n574), .B1(new_n516), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n573), .A2(new_n576), .ZN(G305));
  INV_X1    g152(.A(G85), .ZN(new_n578));
  INV_X1    g153(.A(G47), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n522), .A2(new_n578), .B1(new_n516), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n527), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G290));
  INV_X1    g159(.A(G868), .ZN(new_n585));
  NOR2_X1   g160(.A1(G301), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n523), .A2(G92), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT10), .Z(new_n588));
  NAND2_X1  g163(.A1(new_n521), .A2(G66), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n527), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(G54), .B2(new_n517), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n588), .A2(KEYINPUT76), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT76), .B1(new_n588), .B2(new_n592), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n586), .B1(new_n596), .B2(new_n585), .ZN(G284));
  AOI21_X1  g172(.A(new_n586), .B1(new_n596), .B2(new_n585), .ZN(G321));
  NAND2_X1  g173(.A1(G299), .A2(new_n585), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n585), .B2(G168), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(new_n585), .B2(G168), .ZN(G280));
  NOR2_X1   g176(.A1(new_n595), .A2(G559), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(G860), .B2(new_n596), .ZN(G148));
  NAND2_X1  g178(.A1(new_n549), .A2(new_n585), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n602), .B2(new_n585), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n488), .A2(G123), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n487), .A2(G111), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G135), .B2(new_n474), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT77), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2096), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n487), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  XOR2_X1   g190(.A(KEYINPUT13), .B(G2100), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(G156));
  INV_X1    g193(.A(KEYINPUT14), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(new_n621), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n624), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G14), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n629), .A2(new_n630), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(G401));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT78), .ZN(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n638), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT17), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(G2072), .A2(G2078), .ZN(new_n645));
  OAI22_X1  g220(.A1(new_n639), .A2(new_n643), .B1(new_n445), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2096), .B(G2100), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT79), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n652), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n655), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n652), .A2(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT80), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(KEYINPUT80), .ZN(new_n662));
  AOI211_X1 g237(.A(new_n657), .B(new_n659), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT84), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(G166), .B2(new_n671), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n674), .A2(G1971), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(G1971), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(G23), .ZN(new_n677));
  INV_X1    g252(.A(new_n569), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(new_n671), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT33), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1976), .ZN(new_n681));
  NOR2_X1   g256(.A1(G6), .A2(G16), .ZN(new_n682));
  INV_X1    g257(.A(G305), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G16), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n675), .A2(new_n676), .A3(new_n681), .A4(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT83), .B(KEYINPUT34), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT81), .Z(new_n694));
  OR2_X1    g269(.A1(new_n487), .A2(G107), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n488), .A2(G119), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n474), .A2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(G29), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT82), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n671), .A2(G24), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n583), .B2(new_n671), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n690), .A2(new_n691), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT85), .B(KEYINPUT36), .Z(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NOR2_X1   g287(.A1(G4), .A2(G16), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n596), .B2(G16), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT86), .B(G1348), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n474), .A2(G141), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n488), .A2(G129), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT26), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(G105), .B2(new_n482), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n717), .A2(new_n718), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n692), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n692), .B2(G32), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n612), .A2(G29), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n716), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n692), .A2(G35), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G162), .B2(new_n692), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT29), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n730), .B1(G2090), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(G2090), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT90), .Z(new_n737));
  NOR2_X1   g312(.A1(G27), .A2(G29), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G164), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(new_n444), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G11), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT30), .B(G28), .Z(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n671), .A2(G19), .ZN(new_n744));
  INV_X1    g319(.A(new_n549), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n671), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1341), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  NOR2_X1   g323(.A1(G5), .A2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT88), .Z(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G301), .B2(new_n671), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n743), .B(new_n747), .C1(new_n748), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n671), .A2(G20), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT23), .Z(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G299), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n752), .B(new_n756), .C1(new_n727), .C2(new_n728), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n671), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n671), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n474), .A2(G139), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n762));
  NAND3_X1  g337(.A1(new_n487), .A2(G103), .A3(G2104), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  INV_X1    g341(.A(G127), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n479), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n764), .A2(new_n765), .B1(G2105), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n692), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n692), .B2(G33), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n760), .B1(new_n443), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G2084), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT24), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G34), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n484), .B2(G29), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n774), .B1(new_n443), .B2(new_n773), .C1(new_n775), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n751), .A2(new_n748), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT89), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n692), .A2(G26), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT28), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n474), .A2(G140), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n488), .A2(G128), .ZN(new_n788));
  OR2_X1    g363(.A1(G104), .A2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n789), .B(G2104), .C1(G116), .C2(new_n487), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n786), .B1(new_n791), .B2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2067), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n781), .A2(new_n775), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n759), .A2(G1966), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n784), .A2(new_n793), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n757), .A2(new_n782), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n735), .A2(new_n737), .A3(new_n740), .A4(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n711), .A2(new_n712), .A3(new_n798), .ZN(G311));
  INV_X1    g374(.A(G311), .ZN(G150));
  NAND2_X1  g375(.A1(new_n596), .A2(G559), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT38), .Z(new_n802));
  AOI22_X1  g377(.A1(G93), .A2(new_n523), .B1(new_n517), .B2(G55), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(new_n527), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(new_n549), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n802), .B(new_n807), .Z(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n809), .A2(new_n550), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n806), .A2(new_n550), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(G145));
  XNOR2_X1  g389(.A(new_n612), .B(G160), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(new_n492), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n512), .B2(new_n498), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n819), .A2(KEYINPUT91), .A3(new_n497), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n509), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n791), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(new_n724), .ZN(new_n823));
  INV_X1    g398(.A(new_n791), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n821), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n725), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(new_n770), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n823), .A2(new_n826), .A3(new_n771), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n474), .A2(G142), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n488), .A2(G130), .ZN(new_n832));
  OR2_X1    g407(.A1(G106), .A2(G2105), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n833), .B(G2104), .C1(G118), .C2(new_n487), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n700), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n615), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n698), .A2(KEYINPUT92), .A3(new_n699), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n840), .A2(new_n841), .A3(new_n835), .ZN(new_n845));
  OR3_X1    g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n830), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n830), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n830), .A2(new_n848), .A3(KEYINPUT94), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT94), .B1(new_n830), .B2(new_n848), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n816), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g434(.A(KEYINPUT96), .B(new_n816), .C1(new_n852), .C2(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n830), .A2(new_n845), .A3(new_n843), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n816), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n855), .B2(new_n854), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT40), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n869));
  AOI211_X1 g444(.A(new_n869), .B(new_n866), .C1(new_n859), .C2(new_n860), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(new_n870), .ZN(G395));
  NAND2_X1  g446(.A1(new_n806), .A2(new_n585), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n602), .B(new_n807), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n588), .A2(new_n592), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G299), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT97), .B(KEYINPUT41), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(KEYINPUT41), .B2(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n876), .B(G299), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n874), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(KEYINPUT99), .ZN(new_n886));
  NAND2_X1  g461(.A1(G166), .A2(new_n683), .ZN(new_n887));
  NAND2_X1  g462(.A1(G303), .A2(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n583), .B(new_n569), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT98), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(KEYINPUT98), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n892), .A2(new_n893), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n885), .A2(KEYINPUT99), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n886), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n900), .ZN(new_n903));
  OAI211_X1 g478(.A(KEYINPUT99), .B(new_n885), .C1(new_n903), .C2(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n873), .B1(new_n905), .B2(G868), .ZN(G295));
  XNOR2_X1  g481(.A(G295), .B(KEYINPUT100), .ZN(G331));
  NAND2_X1  g482(.A1(new_n897), .A2(KEYINPUT102), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n895), .B2(new_n896), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n807), .B(G301), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n911), .A2(G286), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(G286), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n912), .A2(new_n881), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n877), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n908), .B(new_n910), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n897), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n915), .A2(KEYINPUT104), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n883), .A2(new_n878), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(KEYINPUT103), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n877), .A2(KEYINPUT41), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(KEYINPUT103), .A3(new_n924), .ZN(new_n925));
  AND4_X1   g500(.A1(new_n912), .A2(new_n923), .A3(new_n913), .A4(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n915), .A2(KEYINPUT104), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n921), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n908), .A2(new_n910), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n918), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n920), .B1(KEYINPUT43), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT105), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n916), .A2(new_n935), .A3(new_n918), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n936), .A2(KEYINPUT106), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(KEYINPUT106), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n937), .A2(KEYINPUT44), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n931), .A2(new_n941), .A3(new_n932), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n940), .A3(new_n942), .ZN(G397));
  AOI21_X1  g518(.A(KEYINPUT91), .B1(new_n819), .B2(new_n497), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n817), .B(new_n498), .C1(new_n502), .C2(KEYINPUT4), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n511), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT45), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(G160), .A2(G40), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(G1996), .ZN(new_n952));
  NAND2_X1  g527(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G2067), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n791), .B(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(new_n725), .ZN(new_n957));
  OAI221_X1 g532(.A(new_n954), .B1(KEYINPUT125), .B2(KEYINPUT46), .C1(new_n951), .C2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n724), .B(G1996), .Z(new_n960));
  AND2_X1   g535(.A1(new_n960), .A2(new_n956), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT124), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n824), .A2(new_n955), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n951), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n951), .A2(G1986), .A3(G290), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n967), .A2(KEYINPUT48), .ZN(new_n968));
  INV_X1    g543(.A(new_n702), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n700), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n961), .A2(new_n962), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n951), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n967), .A2(KEYINPUT48), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n966), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n959), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT126), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT122), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n946), .A2(new_n978), .A3(new_n947), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n946), .A2(KEYINPUT108), .A3(new_n978), .A4(new_n947), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n510), .A2(new_n947), .A3(new_n513), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n949), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n981), .A2(new_n775), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n821), .B2(G1384), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n513), .A4(new_n947), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n950), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1966), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G8), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n994));
  NAND2_X1  g569(.A1(G286), .A2(G8), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT116), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT51), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n985), .B2(new_n991), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(new_n998), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n997), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT62), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n977), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n946), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n983), .A2(new_n986), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n950), .ZN(new_n1009));
  INV_X1    g584(.A(G1971), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT109), .B(G2090), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n981), .A2(new_n982), .A3(new_n984), .A4(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(KEYINPUT107), .A3(new_n1010), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G303), .A2(G8), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT55), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(G8), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n978), .B1(new_n946), .B2(new_n947), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n510), .A2(new_n978), .A3(new_n513), .A4(new_n947), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n950), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1025), .A2(new_n1014), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n1026), .B2(new_n1001), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n1001), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n678), .A2(G1976), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G305), .B(KEYINPUT49), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n573), .B2(KEYINPUT110), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1030), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1028), .A2(G8), .A3(new_n1031), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1034), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1021), .A2(new_n1027), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n748), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1007), .A2(new_n1008), .A3(new_n444), .A4(new_n950), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1048));
  AND3_X1   g623(.A1(new_n1047), .A2(KEYINPUT119), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT119), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n946), .A2(new_n947), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n949), .B1(new_n1052), .B2(new_n986), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n444), .A4(new_n988), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n987), .A2(new_n444), .A3(new_n950), .A4(new_n988), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT117), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1055), .A2(new_n1057), .A3(KEYINPUT53), .ZN(new_n1058));
  OAI21_X1  g633(.A(G171), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1044), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n999), .B(KEYINPUT51), .C1(new_n1002), .C2(new_n998), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1062), .A2(KEYINPUT122), .A3(KEYINPUT62), .A4(new_n997), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1006), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G288), .A2(G1976), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1039), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G305), .A2(G1981), .ZN(new_n1067));
  XOR2_X1   g642(.A(new_n1067), .B(KEYINPUT111), .Z(new_n1068));
  OAI21_X1  g643(.A(new_n1030), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1021), .B2(new_n1042), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT112), .B(KEYINPUT63), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1002), .A2(G168), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1044), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1017), .A2(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1019), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1002), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1021), .A3(new_n1043), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1070), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT113), .B(G1956), .Z(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1007), .A2(new_n1008), .A3(new_n950), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(G299), .B(KEYINPUT57), .Z(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1045), .A2(new_n1087), .B1(new_n955), .B2(new_n1029), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1088), .B2(new_n595), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1089), .A2(KEYINPUT114), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT114), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1045), .A2(new_n1087), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1029), .A2(new_n955), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n595), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n596), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1084), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT115), .B1(new_n1090), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT61), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT58), .B(G1341), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1009), .A2(G1996), .B1(new_n1029), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n745), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT59), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT115), .B(new_n1111), .C1(new_n1090), .C2(new_n1104), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1103), .A2(new_n1106), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1094), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1044), .A2(new_n1004), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n444), .A2(KEYINPUT53), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n949), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n950), .A2(KEYINPUT121), .ZN(new_n1119));
  AND4_X1   g694(.A1(new_n1007), .A2(new_n987), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1046), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1047), .A2(KEYINPUT119), .A3(new_n1048), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1045), .A2(KEYINPUT120), .A3(new_n748), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1122), .A2(new_n1127), .A3(G301), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1059), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1055), .A2(new_n1057), .A3(KEYINPUT53), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1127), .A2(G301), .A3(new_n1133), .A4(new_n1046), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1122), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1135));
  OAI211_X1 g710(.A(KEYINPUT54), .B(new_n1134), .C1(new_n1135), .C2(G301), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1115), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1064), .B(new_n1078), .C1(new_n1114), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n1139));
  INV_X1    g714(.A(G1986), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n583), .B(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n972), .B1(new_n971), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1138), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n976), .B1(new_n1143), .B2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g720(.A1(new_n861), .A2(new_n867), .ZN(new_n1147));
  OAI21_X1  g721(.A(G319), .B1(new_n632), .B2(new_n633), .ZN(new_n1148));
  NOR2_X1   g722(.A1(G227), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g723(.A1(new_n1149), .A2(KEYINPUT127), .ZN(new_n1150));
  AND2_X1   g724(.A1(new_n1149), .A2(KEYINPUT127), .ZN(new_n1151));
  NOR3_X1   g725(.A1(G229), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AND3_X1   g726(.A1(new_n1147), .A2(new_n931), .A3(new_n1152), .ZN(G308));
  NAND3_X1  g727(.A1(new_n1147), .A2(new_n931), .A3(new_n1152), .ZN(G225));
endmodule


