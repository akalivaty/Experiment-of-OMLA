

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742;

  INV_X1 U362 ( .A(n614), .ZN(n341) );
  INV_X1 U363 ( .A(KEYINPUT56), .ZN(n343) );
  AND2_X1 U364 ( .A1(n632), .A2(n609), .ZN(n709) );
  NAND2_X1 U365 ( .A1(n715), .A2(n607), .ZN(n608) );
  NAND2_X1 U366 ( .A1(n388), .A2(n348), .ZN(n387) );
  NOR2_X1 U367 ( .A1(n742), .A2(n616), .ZN(n561) );
  OR2_X1 U368 ( .A1(n570), .A2(n476), .ZN(n477) );
  XNOR2_X1 U369 ( .A(n566), .B(n468), .ZN(n570) );
  BUF_X1 U370 ( .A(G953), .Z(n339) );
  XNOR2_X1 U371 ( .A(n452), .B(KEYINPUT90), .ZN(n453) );
  NAND2_X1 U372 ( .A1(n451), .A2(G224), .ZN(n452) );
  INV_X2 U373 ( .A(G953), .ZN(n451) );
  XNOR2_X2 U374 ( .A(n405), .B(n404), .ZN(n566) );
  NAND2_X1 U375 ( .A1(n340), .A2(n376), .ZN(n373) );
  NAND2_X1 U376 ( .A1(n375), .A2(KEYINPUT108), .ZN(n340) );
  XNOR2_X2 U377 ( .A(n384), .B(n407), .ZN(n381) );
  XNOR2_X1 U378 ( .A(n342), .B(n341), .ZN(G57) );
  NAND2_X1 U379 ( .A1(n356), .A2(n364), .ZN(n342) );
  XNOR2_X1 U380 ( .A(n344), .B(n343), .ZN(G51) );
  NAND2_X1 U381 ( .A1(n357), .A2(n364), .ZN(n344) );
  INV_X1 U382 ( .A(G902), .ZN(n446) );
  BUF_X1 U383 ( .A(n451), .Z(n736) );
  XNOR2_X2 U384 ( .A(n385), .B(KEYINPUT74), .ZN(n525) );
  NOR2_X2 U385 ( .A1(n514), .A2(n639), .ZN(n385) );
  NAND2_X2 U386 ( .A1(n529), .A2(n511), .ZN(n513) );
  XNOR2_X2 U387 ( .A(n550), .B(n448), .ZN(n562) );
  XNOR2_X2 U388 ( .A(n547), .B(n546), .ZN(n742) );
  XNOR2_X2 U389 ( .A(n508), .B(KEYINPUT35), .ZN(n631) );
  NOR2_X2 U390 ( .A1(n507), .A2(n581), .ZN(n508) );
  XNOR2_X2 U391 ( .A(n387), .B(n386), .ZN(n602) );
  INV_X2 U392 ( .A(n526), .ZN(n645) );
  INV_X1 U393 ( .A(G137), .ZN(n430) );
  AND2_X1 U394 ( .A1(n392), .A2(n406), .ZN(n579) );
  AND2_X1 U395 ( .A1(n378), .A2(n377), .ZN(n392) );
  AND2_X1 U396 ( .A1(n427), .A2(n636), .ZN(n393) );
  XNOR2_X1 U397 ( .A(n552), .B(KEYINPUT1), .ZN(n514) );
  XNOR2_X1 U398 ( .A(n437), .B(G469), .ZN(n552) );
  NOR2_X1 U399 ( .A1(G902), .A2(n700), .ZN(n437) );
  XNOR2_X1 U400 ( .A(n445), .B(n436), .ZN(n700) );
  XNOR2_X1 U401 ( .A(n428), .B(G128), .ZN(n458) );
  XNOR2_X1 U402 ( .A(n430), .B(G131), .ZN(n407) );
  XNOR2_X1 U403 ( .A(n416), .B(n446), .ZN(n601) );
  XNOR2_X1 U404 ( .A(n395), .B(G125), .ZN(n455) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n478) );
  NAND2_X1 U406 ( .A1(n392), .A2(n545), .ZN(n355) );
  AND2_X2 U407 ( .A1(n632), .A2(n609), .ZN(n345) );
  INV_X1 U408 ( .A(G143), .ZN(n428) );
  INV_X1 U409 ( .A(G146), .ZN(n395) );
  INV_X1 U410 ( .A(KEYINPUT68), .ZN(n439) );
  XNOR2_X1 U411 ( .A(n433), .B(n432), .ZN(n460) );
  INV_X1 U412 ( .A(G104), .ZN(n432) );
  NAND2_X1 U413 ( .A1(n372), .A2(n379), .ZN(n371) );
  INV_X1 U414 ( .A(n549), .ZN(n379) );
  NAND2_X1 U415 ( .A1(n639), .A2(KEYINPUT108), .ZN(n372) );
  XNOR2_X1 U416 ( .A(n455), .B(n394), .ZN(n728) );
  XNOR2_X1 U417 ( .A(G140), .B(KEYINPUT10), .ZN(n394) );
  XNOR2_X1 U418 ( .A(n362), .B(n411), .ZN(n413) );
  XNOR2_X1 U419 ( .A(n410), .B(n363), .ZN(n362) );
  INV_X1 U420 ( .A(KEYINPUT23), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n458), .B(n429), .ZN(n488) );
  INV_X1 U422 ( .A(G134), .ZN(n429) );
  XNOR2_X1 U423 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U424 ( .A(G107), .B(KEYINPUT7), .Z(n482) );
  BUF_X1 U425 ( .A(n595), .Z(n366) );
  XNOR2_X1 U426 ( .A(G119), .B(G116), .ZN(n438) );
  XNOR2_X1 U427 ( .A(G128), .B(G137), .ZN(n410) );
  INV_X1 U428 ( .A(KEYINPUT45), .ZN(n386) );
  XNOR2_X1 U429 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n588) );
  NAND2_X1 U430 ( .A1(n645), .A2(n368), .ZN(n367) );
  NOR2_X1 U431 ( .A1(n654), .A2(n543), .ZN(n368) );
  NAND2_X1 U432 ( .A1(n654), .A2(n543), .ZN(n369) );
  XNOR2_X1 U433 ( .A(KEYINPUT93), .B(KEYINPUT15), .ZN(n416) );
  XNOR2_X1 U434 ( .A(n454), .B(n458), .ZN(n401) );
  XOR2_X1 U435 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n454) );
  XNOR2_X1 U436 ( .A(n455), .B(n457), .ZN(n399) );
  XNOR2_X1 U437 ( .A(KEYINPUT17), .B(KEYINPUT94), .ZN(n457) );
  XNOR2_X1 U438 ( .A(n459), .B(n403), .ZN(n722) );
  XNOR2_X1 U439 ( .A(n460), .B(n346), .ZN(n403) );
  INV_X1 U440 ( .A(KEYINPUT88), .ZN(n404) );
  XNOR2_X1 U441 ( .A(n361), .B(n360), .ZN(n590) );
  INV_X1 U442 ( .A(KEYINPUT106), .ZN(n360) );
  INV_X1 U443 ( .A(n515), .ZN(n427) );
  BUF_X1 U444 ( .A(n514), .Z(n638) );
  INV_X1 U445 ( .A(KEYINPUT6), .ZN(n448) );
  XNOR2_X1 U446 ( .A(G119), .B(G110), .ZN(n412) );
  XNOR2_X1 U447 ( .A(n484), .B(n483), .ZN(n486) );
  INV_X1 U448 ( .A(n366), .ZN(n406) );
  XNOR2_X1 U449 ( .A(n359), .B(n358), .ZN(G60) );
  INV_X1 U450 ( .A(KEYINPUT60), .ZN(n358) );
  XOR2_X1 U451 ( .A(KEYINPUT16), .B(G122), .Z(n346) );
  XOR2_X1 U452 ( .A(n456), .B(G146), .Z(n347) );
  INV_X1 U453 ( .A(n550), .ZN(n526) );
  AND2_X1 U454 ( .A1(n539), .A2(n618), .ZN(n348) );
  AND2_X1 U455 ( .A1(n370), .A2(n369), .ZN(n349) );
  AND2_X1 U456 ( .A1(n393), .A2(n380), .ZN(n350) );
  INV_X1 U457 ( .A(KEYINPUT108), .ZN(n380) );
  XOR2_X1 U458 ( .A(n629), .B(n628), .Z(n351) );
  XOR2_X1 U459 ( .A(n624), .B(n623), .Z(n352) );
  XOR2_X1 U460 ( .A(n610), .B(n611), .Z(n353) );
  AND2_X1 U461 ( .A1(n613), .A2(n339), .ZN(n714) );
  INV_X1 U462 ( .A(n714), .ZN(n364) );
  XNOR2_X2 U463 ( .A(n354), .B(KEYINPUT86), .ZN(n731) );
  NAND2_X2 U464 ( .A1(n605), .A2(n603), .ZN(n354) );
  NOR2_X1 U465 ( .A1(n373), .A2(n371), .ZN(n378) );
  XNOR2_X2 U466 ( .A(n355), .B(KEYINPUT39), .ZN(n597) );
  AND2_X1 U467 ( .A1(n578), .A2(n577), .ZN(n587) );
  NAND2_X1 U468 ( .A1(n597), .A2(n689), .ZN(n547) );
  XNOR2_X1 U469 ( .A(n612), .B(n353), .ZN(n356) );
  XNOR2_X1 U470 ( .A(n625), .B(n352), .ZN(n357) );
  NAND2_X1 U471 ( .A1(n365), .A2(n364), .ZN(n359) );
  NAND2_X1 U472 ( .A1(n565), .A2(n689), .ZN(n361) );
  OR2_X1 U473 ( .A1(n550), .A2(KEYINPUT30), .ZN(n370) );
  NOR2_X2 U474 ( .A1(n580), .A2(n581), .ZN(n688) );
  INV_X1 U475 ( .A(n393), .ZN(n639) );
  AND2_X1 U476 ( .A1(n631), .A2(n617), .ZN(n391) );
  XNOR2_X1 U477 ( .A(n630), .B(n351), .ZN(n365) );
  NAND2_X1 U478 ( .A1(n349), .A2(n367), .ZN(n377) );
  NAND2_X1 U479 ( .A1(n553), .A2(n393), .ZN(n383) );
  INV_X1 U480 ( .A(n553), .ZN(n375) );
  NAND2_X1 U481 ( .A1(n350), .A2(n553), .ZN(n376) );
  XNOR2_X2 U482 ( .A(n381), .B(n488), .ZN(n729) );
  XNOR2_X2 U483 ( .A(n382), .B(KEYINPUT64), .ZN(n384) );
  XNOR2_X2 U484 ( .A(KEYINPUT4), .B(KEYINPUT66), .ZN(n382) );
  NOR2_X1 U485 ( .A1(n645), .A2(n383), .ZN(n530) );
  XNOR2_X2 U486 ( .A(n523), .B(n522), .ZN(n619) );
  XNOR2_X1 U487 ( .A(n384), .B(n399), .ZN(n398) );
  NAND2_X1 U488 ( .A1(n525), .A2(n562), .ZN(n450) );
  XNOR2_X1 U489 ( .A(n389), .B(n524), .ZN(n388) );
  NAND2_X1 U490 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U491 ( .A(n619), .ZN(n390) );
  NAND2_X1 U492 ( .A1(n396), .A2(n521), .ZN(n523) );
  NAND2_X1 U493 ( .A1(n396), .A2(n537), .ZN(n538) );
  NAND2_X1 U494 ( .A1(n396), .A2(n517), .ZN(n617) );
  XNOR2_X2 U495 ( .A(n513), .B(n512), .ZN(n396) );
  XNOR2_X1 U496 ( .A(n397), .B(n722), .ZN(n624) );
  XNOR2_X1 U497 ( .A(n400), .B(n398), .ZN(n397) );
  XNOR2_X1 U498 ( .A(n402), .B(n401), .ZN(n400) );
  XNOR2_X1 U499 ( .A(n453), .B(n456), .ZN(n402) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n459) );
  NOR2_X2 U501 ( .A1(n595), .A2(n654), .ZN(n405) );
  XNOR2_X2 U502 ( .A(n465), .B(n464), .ZN(n595) );
  AND2_X1 U503 ( .A1(G221), .A2(n480), .ZN(n408) );
  AND2_X1 U504 ( .A1(n603), .A2(KEYINPUT2), .ZN(n604) );
  NAND2_X1 U505 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U506 ( .A(n443), .B(KEYINPUT5), .ZN(n444) );
  INV_X1 U507 ( .A(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n610) );
  INV_X1 U509 ( .A(KEYINPUT9), .ZN(n481) );
  INV_X1 U510 ( .A(KEYINPUT30), .ZN(n543) );
  NAND2_X1 U511 ( .A1(G234), .A2(n451), .ZN(n409) );
  XOR2_X1 U512 ( .A(KEYINPUT8), .B(n409), .Z(n480) );
  XNOR2_X1 U513 ( .A(n728), .B(n408), .ZN(n415) );
  XOR2_X1 U514 ( .A(KEYINPUT24), .B(KEYINPUT96), .Z(n411) );
  XNOR2_X1 U515 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U516 ( .A(n415), .B(n414), .ZN(n710) );
  NOR2_X1 U517 ( .A1(n710), .A2(G902), .ZN(n421) );
  NAND2_X1 U518 ( .A1(G234), .A2(n601), .ZN(n417) );
  XNOR2_X1 U519 ( .A(KEYINPUT20), .B(n417), .ZN(n422) );
  NAND2_X1 U520 ( .A1(G217), .A2(n422), .ZN(n419) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n418) );
  XNOR2_X1 U522 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X2 U523 ( .A(n421), .B(n420), .ZN(n515) );
  NAND2_X1 U524 ( .A1(G221), .A2(n422), .ZN(n426) );
  XOR2_X1 U525 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n424) );
  INV_X1 U526 ( .A(KEYINPUT97), .ZN(n423) );
  XNOR2_X1 U527 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U528 ( .A(n426), .B(n425), .ZN(n636) );
  INV_X1 U529 ( .A(n636), .ZN(n510) );
  INV_X1 U530 ( .A(KEYINPUT65), .ZN(n431) );
  XNOR2_X1 U531 ( .A(n431), .B(G101), .ZN(n456) );
  XNOR2_X2 U532 ( .A(n729), .B(n347), .ZN(n445) );
  XNOR2_X1 U533 ( .A(G110), .B(G107), .ZN(n433) );
  NAND2_X1 U534 ( .A1(G227), .A2(n736), .ZN(n434) );
  XNOR2_X1 U535 ( .A(n434), .B(G140), .ZN(n435) );
  XNOR2_X1 U536 ( .A(n460), .B(n435), .ZN(n436) );
  XNOR2_X1 U537 ( .A(n438), .B(KEYINPUT3), .ZN(n441) );
  XNOR2_X1 U538 ( .A(n439), .B(G113), .ZN(n440) );
  NOR2_X1 U539 ( .A1(G953), .A2(G237), .ZN(n496) );
  NAND2_X1 U540 ( .A1(n496), .A2(G210), .ZN(n442) );
  XNOR2_X1 U541 ( .A(n459), .B(n442), .ZN(n443) );
  NAND2_X1 U542 ( .A1(n610), .A2(n446), .ZN(n447) );
  XNOR2_X2 U543 ( .A(n447), .B(G472), .ZN(n550) );
  XNOR2_X1 U544 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n449) );
  XNOR2_X1 U545 ( .A(n450), .B(n449), .ZN(n651) );
  NAND2_X1 U546 ( .A1(n624), .A2(n601), .ZN(n465) );
  NOR2_X1 U547 ( .A1(G902), .A2(G237), .ZN(n462) );
  INV_X1 U548 ( .A(KEYINPUT75), .ZN(n461) );
  XNOR2_X1 U549 ( .A(n462), .B(n461), .ZN(n467) );
  INV_X1 U550 ( .A(n467), .ZN(n463) );
  NAND2_X1 U551 ( .A1(n463), .A2(G210), .ZN(n464) );
  INV_X1 U552 ( .A(G214), .ZN(n466) );
  OR2_X1 U553 ( .A1(n467), .A2(n466), .ZN(n591) );
  INV_X1 U554 ( .A(n591), .ZN(n654) );
  XNOR2_X1 U555 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n468) );
  NAND2_X1 U556 ( .A1(G234), .A2(G237), .ZN(n469) );
  XNOR2_X1 U557 ( .A(n469), .B(KEYINPUT14), .ZN(n470) );
  XNOR2_X1 U558 ( .A(KEYINPUT72), .B(n470), .ZN(n473) );
  AND2_X1 U559 ( .A1(n473), .A2(n339), .ZN(n471) );
  NAND2_X1 U560 ( .A1(G902), .A2(n471), .ZN(n540) );
  NOR2_X1 U561 ( .A1(G898), .A2(n540), .ZN(n472) );
  XNOR2_X1 U562 ( .A(n472), .B(KEYINPUT95), .ZN(n475) );
  AND2_X1 U563 ( .A1(n473), .A2(G952), .ZN(n667) );
  AND2_X1 U564 ( .A1(n667), .A2(n736), .ZN(n542) );
  INV_X1 U565 ( .A(n542), .ZN(n474) );
  AND2_X1 U566 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X2 U567 ( .A(n477), .B(KEYINPUT0), .ZN(n527) );
  NOR2_X1 U568 ( .A1(n651), .A2(n527), .ZN(n479) );
  XNOR2_X1 U569 ( .A(n479), .B(n478), .ZN(n507) );
  NAND2_X1 U570 ( .A1(G217), .A2(n480), .ZN(n484) );
  XNOR2_X1 U571 ( .A(G116), .B(G122), .ZN(n485) );
  XNOR2_X1 U572 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U573 ( .A(n488), .B(n487), .ZN(n707) );
  NOR2_X1 U574 ( .A1(G902), .A2(n707), .ZN(n490) );
  XNOR2_X1 U575 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U576 ( .A(n490), .B(n489), .ZN(n492) );
  INV_X1 U577 ( .A(G478), .ZN(n491) );
  XNOR2_X1 U578 ( .A(n492), .B(n491), .ZN(n533) );
  INV_X1 U579 ( .A(n533), .ZN(n506) );
  XNOR2_X1 U580 ( .A(KEYINPUT13), .B(G475), .ZN(n505) );
  XOR2_X1 U581 ( .A(KEYINPUT11), .B(G104), .Z(n494) );
  XNOR2_X1 U582 ( .A(G131), .B(G143), .ZN(n493) );
  XNOR2_X1 U583 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U584 ( .A(n728), .B(n495), .ZN(n503) );
  XOR2_X1 U585 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n498) );
  NAND2_X1 U586 ( .A1(G214), .A2(n496), .ZN(n497) );
  XNOR2_X1 U587 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U588 ( .A(n499), .B(KEYINPUT100), .Z(n501) );
  XNOR2_X1 U589 ( .A(G113), .B(G122), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U591 ( .A(n503), .B(n502), .ZN(n629) );
  NOR2_X1 U592 ( .A1(G902), .A2(n629), .ZN(n504) );
  XNOR2_X1 U593 ( .A(n505), .B(n504), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n506), .A2(n532), .ZN(n581) );
  INV_X1 U595 ( .A(n527), .ZN(n529) );
  INV_X1 U596 ( .A(n532), .ZN(n509) );
  NAND2_X1 U597 ( .A1(n533), .A2(n509), .ZN(n657) );
  NOR2_X1 U598 ( .A1(n657), .A2(n510), .ZN(n511) );
  XNOR2_X1 U599 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n512) );
  INV_X1 U600 ( .A(n638), .ZN(n518) );
  NAND2_X1 U601 ( .A1(n526), .A2(n515), .ZN(n516) );
  NOR2_X1 U602 ( .A1(n518), .A2(n516), .ZN(n517) );
  NAND2_X1 U603 ( .A1(n518), .A2(n515), .ZN(n519) );
  NOR2_X1 U604 ( .A1(n562), .A2(n519), .ZN(n520) );
  XOR2_X1 U605 ( .A(KEYINPUT81), .B(n520), .Z(n521) );
  XOR2_X1 U606 ( .A(KEYINPUT80), .B(KEYINPUT32), .Z(n522) );
  NAND2_X1 U607 ( .A1(n525), .A2(n645), .ZN(n647) );
  NOR2_X1 U608 ( .A1(n647), .A2(n527), .ZN(n528) );
  XNOR2_X1 U609 ( .A(n528), .B(KEYINPUT31), .ZN(n695) );
  NAND2_X1 U610 ( .A1(n529), .A2(n530), .ZN(n680) );
  NAND2_X1 U611 ( .A1(n695), .A2(n680), .ZN(n535) );
  NAND2_X1 U612 ( .A1(n532), .A2(n533), .ZN(n531) );
  XNOR2_X2 U613 ( .A(KEYINPUT103), .B(n531), .ZN(n689) );
  OR2_X1 U614 ( .A1(n533), .A2(n532), .ZN(n696) );
  INV_X1 U615 ( .A(n696), .ZN(n684) );
  NOR2_X1 U616 ( .A1(n689), .A2(n684), .ZN(n653) );
  INV_X1 U617 ( .A(n653), .ZN(n534) );
  NAND2_X1 U618 ( .A1(n535), .A2(n534), .ZN(n539) );
  INV_X1 U619 ( .A(n515), .ZN(n635) );
  NAND2_X1 U620 ( .A1(n638), .A2(n635), .ZN(n536) );
  NOR2_X1 U621 ( .A1(n562), .A2(n536), .ZN(n537) );
  XNOR2_X1 U622 ( .A(n538), .B(KEYINPUT104), .ZN(n618) );
  NOR2_X1 U623 ( .A1(G900), .A2(n540), .ZN(n541) );
  NOR2_X1 U624 ( .A1(n542), .A2(n541), .ZN(n549) );
  XNOR2_X1 U625 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n544) );
  XNOR2_X1 U626 ( .A(n595), .B(n544), .ZN(n655) );
  INV_X1 U627 ( .A(n655), .ZN(n545) );
  INV_X1 U628 ( .A(KEYINPUT40), .ZN(n546) );
  NAND2_X1 U629 ( .A1(n636), .A2(n515), .ZN(n548) );
  NOR2_X1 U630 ( .A1(n549), .A2(n548), .ZN(n563) );
  AND2_X1 U631 ( .A1(n563), .A2(n645), .ZN(n551) );
  XNOR2_X1 U632 ( .A(n551), .B(KEYINPUT28), .ZN(n554) );
  INV_X1 U633 ( .A(n552), .ZN(n553) );
  AND2_X1 U634 ( .A1(n554), .A2(n553), .ZN(n572) );
  INV_X1 U635 ( .A(n657), .ZN(n556) );
  OR2_X1 U636 ( .A1(n655), .A2(n654), .ZN(n652) );
  INV_X1 U637 ( .A(n652), .ZN(n555) );
  NAND2_X1 U638 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U639 ( .A(n557), .B(KEYINPUT41), .ZN(n669) );
  NAND2_X1 U640 ( .A1(n572), .A2(n669), .ZN(n560) );
  INV_X1 U641 ( .A(KEYINPUT110), .ZN(n558) );
  XNOR2_X1 U642 ( .A(n558), .B(KEYINPUT42), .ZN(n559) );
  XNOR2_X1 U643 ( .A(n560), .B(n559), .ZN(n616) );
  XNOR2_X1 U644 ( .A(n561), .B(KEYINPUT46), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n564), .B(KEYINPUT105), .ZN(n565) );
  INV_X1 U646 ( .A(n566), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n590), .A2(n567), .ZN(n568) );
  XNOR2_X1 U648 ( .A(n568), .B(KEYINPUT36), .ZN(n569) );
  NOR2_X2 U649 ( .A1(n569), .A2(n638), .ZN(n698) );
  INV_X1 U650 ( .A(n570), .ZN(n571) );
  NAND2_X1 U651 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U652 ( .A(n573), .B(KEYINPUT47), .ZN(n575) );
  INV_X1 U653 ( .A(n573), .ZN(n690) );
  NAND2_X1 U654 ( .A1(n690), .A2(n653), .ZN(n574) );
  AND2_X1 U655 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U656 ( .A1(n698), .A2(n576), .ZN(n577) );
  XNOR2_X1 U657 ( .A(n579), .B(KEYINPUT109), .ZN(n580) );
  XNOR2_X1 U658 ( .A(n688), .B(KEYINPUT85), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n653), .A2(KEYINPUT47), .ZN(n582) );
  XNOR2_X1 U660 ( .A(KEYINPUT84), .B(n582), .ZN(n583) );
  AND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT82), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X2 U664 ( .A(n589), .B(n588), .ZN(n605) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U666 ( .A(KEYINPUT107), .B(n592), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n593), .A2(n638), .ZN(n594) );
  XNOR2_X1 U668 ( .A(n594), .B(KEYINPUT43), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n596), .A2(n366), .ZN(n620) );
  NAND2_X1 U670 ( .A1(n597), .A2(n684), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT111), .ZN(n741) );
  INV_X1 U672 ( .A(n741), .ZN(n599) );
  AND2_X1 U673 ( .A1(n620), .A2(n599), .ZN(n603) );
  NOR2_X1 U674 ( .A1(n602), .A2(n731), .ZN(n600) );
  NOR2_X1 U675 ( .A1(n600), .A2(KEYINPUT2), .ZN(n633) );
  NOR2_X2 U676 ( .A1(n633), .A2(n601), .ZN(n609) );
  INV_X1 U677 ( .A(n602), .ZN(n715) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT87), .ZN(n607) );
  XNOR2_X2 U680 ( .A(n608), .B(KEYINPUT76), .ZN(n632) );
  NAND2_X1 U681 ( .A1(n709), .A2(G472), .ZN(n612) );
  XNOR2_X1 U682 ( .A(KEYINPUT91), .B(KEYINPUT62), .ZN(n611) );
  INV_X1 U683 ( .A(G952), .ZN(n613) );
  INV_X1 U684 ( .A(KEYINPUT63), .ZN(n614) );
  XOR2_X1 U685 ( .A(G137), .B(n616), .Z(G39) );
  XNOR2_X1 U686 ( .A(n617), .B(G110), .ZN(G12) );
  XNOR2_X1 U687 ( .A(n618), .B(G101), .ZN(G3) );
  XOR2_X1 U688 ( .A(n619), .B(G119), .Z(G21) );
  XNOR2_X1 U689 ( .A(n620), .B(G140), .ZN(G42) );
  NAND2_X1 U690 ( .A1(n709), .A2(G210), .ZN(n625) );
  XOR2_X1 U691 ( .A(KEYINPUT83), .B(KEYINPUT89), .Z(n622) );
  XNOR2_X1 U692 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n621) );
  XOR2_X1 U693 ( .A(n622), .B(n621), .Z(n623) );
  NAND2_X1 U694 ( .A1(n345), .A2(G475), .ZN(n630) );
  XNOR2_X1 U695 ( .A(KEYINPUT92), .B(KEYINPUT120), .ZN(n627) );
  XOR2_X1 U696 ( .A(n627), .B(KEYINPUT59), .Z(n628) );
  XNOR2_X1 U697 ( .A(n631), .B(G122), .ZN(G24) );
  INV_X1 U698 ( .A(n632), .ZN(n634) );
  NOR2_X1 U699 ( .A1(n634), .A2(n633), .ZN(n676) );
  NOR2_X1 U700 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U701 ( .A(KEYINPUT49), .B(n637), .ZN(n643) );
  NAND2_X1 U702 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U703 ( .A(n640), .B(KEYINPUT114), .ZN(n641) );
  XNOR2_X1 U704 ( .A(KEYINPUT50), .B(n641), .ZN(n642) );
  NAND2_X1 U705 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U706 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U707 ( .A(n646), .B(KEYINPUT115), .ZN(n648) );
  NAND2_X1 U708 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U709 ( .A(KEYINPUT51), .B(n649), .Z(n650) );
  NAND2_X1 U710 ( .A1(n650), .A2(n669), .ZN(n664) );
  BUF_X1 U711 ( .A(n651), .Z(n671) );
  INV_X1 U712 ( .A(n671), .ZN(n662) );
  OR2_X1 U713 ( .A1(n653), .A2(n652), .ZN(n659) );
  AND2_X1 U714 ( .A1(n655), .A2(n654), .ZN(n656) );
  OR2_X1 U715 ( .A1(n657), .A2(n656), .ZN(n658) );
  AND2_X1 U716 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U717 ( .A(KEYINPUT116), .B(n660), .Z(n661) );
  NAND2_X1 U718 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U719 ( .A1(n664), .A2(n663), .ZN(n666) );
  XOR2_X1 U720 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n665) );
  XNOR2_X1 U721 ( .A(n666), .B(n665), .ZN(n668) );
  NAND2_X1 U722 ( .A1(n668), .A2(n667), .ZN(n674) );
  INV_X1 U723 ( .A(n669), .ZN(n670) );
  NOR2_X1 U724 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U725 ( .A1(n672), .A2(n339), .ZN(n673) );
  NAND2_X1 U726 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U727 ( .A1(n676), .A2(n675), .ZN(n678) );
  XNOR2_X1 U728 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n677) );
  XNOR2_X1 U729 ( .A(n678), .B(n677), .ZN(G75) );
  INV_X1 U730 ( .A(n689), .ZN(n692) );
  NOR2_X1 U731 ( .A1(n692), .A2(n680), .ZN(n679) );
  XOR2_X1 U732 ( .A(G104), .B(n679), .Z(G6) );
  NOR2_X1 U733 ( .A1(n696), .A2(n680), .ZN(n682) );
  XNOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n681) );
  XNOR2_X1 U735 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U736 ( .A(G107), .B(n683), .ZN(G9) );
  XOR2_X1 U737 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n686) );
  NAND2_X1 U738 ( .A1(n690), .A2(n684), .ZN(n685) );
  XNOR2_X1 U739 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U740 ( .A(G128), .B(n687), .ZN(G30) );
  XOR2_X1 U741 ( .A(n688), .B(G143), .Z(G45) );
  NAND2_X1 U742 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U743 ( .A(n691), .B(G146), .ZN(G48) );
  NOR2_X1 U744 ( .A1(n692), .A2(n695), .ZN(n694) );
  XNOR2_X1 U745 ( .A(G113), .B(KEYINPUT113), .ZN(n693) );
  XNOR2_X1 U746 ( .A(n694), .B(n693), .ZN(G15) );
  NOR2_X1 U747 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U748 ( .A(G116), .B(n697), .Z(G18) );
  XNOR2_X1 U749 ( .A(n698), .B(G125), .ZN(n699) );
  XNOR2_X1 U750 ( .A(n699), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  XNOR2_X1 U752 ( .A(n700), .B(KEYINPUT119), .ZN(n701) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U754 ( .A1(n345), .A2(G469), .ZN(n703) );
  XOR2_X1 U755 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U756 ( .A1(n714), .A2(n705), .ZN(G54) );
  NAND2_X1 U757 ( .A1(n345), .A2(G478), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U759 ( .A1(n714), .A2(n708), .ZN(G63) );
  NAND2_X1 U760 ( .A1(n345), .A2(G217), .ZN(n712) );
  XOR2_X1 U761 ( .A(n710), .B(KEYINPUT121), .Z(n711) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U763 ( .A1(n714), .A2(n713), .ZN(G66) );
  NAND2_X1 U764 ( .A1(n715), .A2(n736), .ZN(n720) );
  NAND2_X1 U765 ( .A1(n339), .A2(G224), .ZN(n716) );
  XNOR2_X1 U766 ( .A(KEYINPUT61), .B(n716), .ZN(n717) );
  NAND2_X1 U767 ( .A1(n717), .A2(G898), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(KEYINPUT122), .ZN(n719) );
  NAND2_X1 U769 ( .A1(n720), .A2(n719), .ZN(n727) );
  XNOR2_X1 U770 ( .A(G101), .B(KEYINPUT123), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n724) );
  NOR2_X1 U772 ( .A1(G898), .A2(n736), .ZN(n723) );
  NOR2_X1 U773 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U774 ( .A(KEYINPUT124), .B(n725), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(G69) );
  XNOR2_X1 U776 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U777 ( .A(n730), .B(KEYINPUT125), .ZN(n734) );
  BUF_X1 U778 ( .A(n731), .Z(n732) );
  XOR2_X1 U779 ( .A(n734), .B(n732), .Z(n733) );
  NAND2_X1 U780 ( .A1(n733), .A2(n736), .ZN(n739) );
  XOR2_X1 U781 ( .A(G227), .B(n734), .Z(n735) );
  NOR2_X1 U782 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U783 ( .A1(G900), .A2(n737), .ZN(n738) );
  NAND2_X1 U784 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U785 ( .A(KEYINPUT126), .B(n740), .Z(G72) );
  XOR2_X1 U786 ( .A(G134), .B(n741), .Z(G36) );
  XOR2_X1 U787 ( .A(n742), .B(G131), .Z(G33) );
endmodule

