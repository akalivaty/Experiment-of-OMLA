//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G190gat), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  OR3_X1    g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT27), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT27), .B1(new_n206), .B2(new_n207), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n205), .B1(new_n211), .B2(new_n203), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  NOR3_X1   g014(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n213), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT69), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n222), .B(new_n213), .C1(new_n218), .C2(new_n219), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n212), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n213), .A2(new_n228), .ZN(new_n229));
  AOI211_X1 g028(.A(new_n227), .B(new_n229), .C1(new_n207), .C2(new_n209), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n214), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n226), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT25), .B1(new_n236), .B2(KEYINPUT64), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n239));
  OAI221_X1 g038(.A(new_n238), .B1(G183gat), .B2(G190gat), .C1(new_n239), .C2(new_n228), .ZN(new_n240));
  OAI211_X1 g039(.A(KEYINPUT25), .B(new_n214), .C1(new_n231), .C2(KEYINPUT23), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n237), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n232), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n235), .B(KEYINPUT66), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n228), .B1(new_n213), .B2(KEYINPUT65), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(new_n207), .B2(new_n209), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n241), .B1(new_n248), .B2(new_n238), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n232), .B1(new_n249), .B2(new_n237), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT66), .B1(new_n250), .B2(new_n235), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n225), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G127gat), .B(G134gat), .Z(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT70), .B1(new_n255), .B2(G113gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n257));
  INV_X1    g056(.A(G113gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(G120gat), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n256), .B(new_n259), .C1(new_n258), .C2(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G120gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n253), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n235), .B1(new_n243), .B2(new_n244), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n245), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n264), .A3(new_n225), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n266), .A2(G227gat), .A3(new_n271), .A4(G233gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT32), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT33), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G15gat), .B(G43gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G71gat), .B(G99gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n278), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n272), .B(KEYINPUT32), .C1(new_n274), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n271), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n224), .B1(new_n269), .B2(new_n245), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n264), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n288), .A2(KEYINPUT34), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(KEYINPUT34), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n266), .A2(new_n271), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n292), .A2(new_n288), .A3(KEYINPUT34), .A4(new_n283), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n282), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n293), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(new_n279), .A3(new_n281), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT36), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(KEYINPUT72), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n304), .B2(new_n299), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT83), .B(G50gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n308), .A3(new_n312), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G141gat), .B(G148gat), .Z(new_n319));
  INV_X1    g118(.A(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G162gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT2), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G155gat), .B(G162gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n324), .A3(new_n322), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n318), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(G228gat), .B2(G233gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n328), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n326), .A2(KEYINPUT77), .A3(new_n328), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n316), .A2(KEYINPUT84), .A3(new_n317), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n314), .B1(new_n312), .B2(new_n308), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT84), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT29), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT3), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT85), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n341), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n327), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n336), .A4(new_n335), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT3), .B1(new_n318), .B2(new_n330), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n326), .B2(new_n328), .ZN(new_n350));
  OAI211_X1 g149(.A(G228gat), .B(G233gat), .C1(new_n350), .C2(new_n331), .ZN(new_n351));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G22gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n348), .B2(new_n351), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n356), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(new_n351), .ZN(new_n360));
  INV_X1    g159(.A(new_n352), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n359), .B1(new_n362), .B2(new_n353), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n307), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n356), .B1(new_n354), .B2(new_n357), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n359), .A3(new_n353), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n306), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT5), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n264), .A2(new_n333), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n261), .A2(new_n326), .A3(new_n263), .A4(new_n328), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(KEYINPUT78), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n264), .A2(new_n374), .A3(new_n333), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n370), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n264), .A2(new_n333), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(new_n264), .A3(new_n329), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n380), .B2(KEYINPUT4), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n326), .A2(KEYINPUT77), .A3(new_n328), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT77), .B1(new_n326), .B2(new_n328), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n265), .B(KEYINPUT4), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n377), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(new_n370), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OAI22_X1  g186(.A1(new_n376), .A2(new_n377), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT79), .B1(new_n378), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n391), .A3(KEYINPUT4), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n265), .B(new_n389), .C1(new_n382), .C2(new_n383), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT5), .B1(new_n394), .B2(new_n380), .ZN(new_n395));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396));
  INV_X1    g195(.A(G85gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n388), .A2(new_n395), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n401), .B1(new_n388), .B2(new_n395), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT80), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n408), .B(new_n401), .C1(new_n388), .C2(new_n395), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n402), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n407), .A2(KEYINPUT81), .A3(new_n404), .A4(new_n409), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n405), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n318), .ZN(new_n415));
  INV_X1    g214(.A(new_n267), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT73), .B1(new_n416), .B2(new_n224), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n225), .A2(new_n418), .A3(new_n267), .ZN(new_n419));
  INV_X1    g218(.A(G226gat), .ZN(new_n420));
  INV_X1    g219(.A(G233gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(KEYINPUT29), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n285), .A2(new_n422), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n415), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n417), .A2(new_n419), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n422), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n252), .A2(new_n423), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n415), .A3(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G64gat), .B(G92gat), .Z(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n434), .B(new_n435), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n427), .A2(new_n431), .A3(KEYINPUT30), .A4(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n422), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n417), .B2(new_n419), .ZN(new_n440));
  INV_X1    g239(.A(new_n423), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n285), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n440), .A2(new_n442), .A3(new_n318), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n436), .B1(new_n443), .B2(new_n426), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT76), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT76), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n438), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n431), .A3(new_n437), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n446), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n369), .B1(new_n414), .B2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n424), .A2(new_n425), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n415), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n429), .A2(new_n318), .A3(new_n430), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n427), .A2(new_n431), .A3(new_n455), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n436), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n405), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n403), .A2(new_n407), .A3(new_n404), .A4(new_n409), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n449), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n436), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n455), .B1(new_n427), .B2(new_n431), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n454), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT87), .B(new_n454), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n444), .A3(new_n438), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n377), .B1(new_n394), .B2(new_n380), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n373), .A2(new_n375), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(KEYINPUT39), .C1(new_n385), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n400), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(KEYINPUT40), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT40), .B1(new_n476), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n402), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n472), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n368), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n453), .B1(new_n471), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n305), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n414), .A2(new_n452), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n295), .A2(new_n368), .A3(new_n297), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n295), .A2(new_n368), .A3(KEYINPUT88), .A4(new_n297), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n302), .B1(new_n295), .B2(new_n297), .ZN(new_n492));
  INV_X1    g291(.A(new_n303), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(new_n369), .ZN(new_n494));
  AOI211_X1 g293(.A(KEYINPUT35), .B(new_n472), .C1(new_n462), .C2(new_n463), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n491), .A2(KEYINPUT35), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n485), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT16), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OR2_X1    g299(.A1(G15gat), .A2(G22gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(G15gat), .A2(G22gat), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT91), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n500), .B1(new_n503), .B2(G1gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n498), .A2(new_n505), .A3(G1gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(G8gat), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT92), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n498), .A2(new_n505), .ZN(new_n510));
  INV_X1    g309(.A(G1gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G8gat), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n506), .A4(new_n500), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT93), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n510), .A2(new_n511), .B1(new_n499), .B2(new_n498), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n513), .A4(new_n506), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT90), .B(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(G29gat), .A2(G36gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT14), .ZN(new_n525));
  OAI211_X1 g324(.A(KEYINPUT15), .B(new_n520), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n525), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n522), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n530), .A3(KEYINPUT17), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n509), .A2(new_n519), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n506), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(G8gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n508), .A2(KEYINPUT92), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n519), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n531), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT94), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n535), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n535), .A2(new_n541), .A3(KEYINPUT18), .A4(new_n544), .ZN(new_n548));
  INV_X1    g347(.A(new_n531), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n509), .A2(new_n549), .A3(new_n519), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n543), .B(KEYINPUT13), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n556));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G169gat), .B(G197gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT12), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n555), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n547), .A2(new_n548), .A3(new_n554), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n561), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n547), .A2(new_n561), .A3(new_n548), .A4(new_n554), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT95), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571));
  INV_X1    g370(.A(G71gat), .ZN(new_n572));
  INV_X1    g371(.A(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G57gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(G64gat), .ZN(new_n576));
  INV_X1    g375(.A(G64gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(G57gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n574), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n576), .B2(new_n578), .ZN(new_n581));
  AND2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G57gat), .B(G64gat), .Z(new_n587));
  OAI211_X1 g386(.A(new_n587), .B(new_n574), .C1(new_n580), .C2(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n540), .B1(KEYINPUT21), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(new_n207), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G211gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n595), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n592), .B(new_n599), .Z(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT8), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT7), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n397), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n602), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G99gat), .B(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n601), .B1(new_n397), .B2(new_n606), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n533), .B(new_n534), .C1(new_n612), .C2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n612), .A2(new_n617), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n531), .A2(new_n619), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT97), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n627), .A2(new_n631), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n600), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n636), .A2(KEYINPUT98), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n619), .A2(new_n589), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n586), .B(new_n588), .C1(new_n612), .C2(new_n617), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n640), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT100), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n647), .A3(new_n643), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n648), .A2(KEYINPUT99), .B1(new_n642), .B2(KEYINPUT10), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n641), .A2(new_n650), .A3(new_n647), .A4(new_n643), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n640), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n646), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n646), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n648), .A2(KEYINPUT99), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n642), .A2(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n651), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n639), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT101), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n663), .A3(new_n639), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n657), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n656), .B1(new_n665), .B2(new_n655), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n637), .A2(new_n638), .A3(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n497), .A2(new_n570), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n412), .A2(new_n413), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT102), .B1(new_n669), .B2(new_n405), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n414), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g474(.A1(new_n668), .A2(new_n472), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT42), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(G8gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT103), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(G1325gat));
  INV_X1    g481(.A(new_n304), .ZN(new_n683));
  AOI21_X1  g482(.A(G15gat), .B1(new_n668), .B2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n305), .A2(G15gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n684), .B1(new_n668), .B2(new_n685), .ZN(G1326gat));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n369), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n494), .A2(new_n495), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n299), .B1(new_n492), .B2(new_n493), .ZN(new_n693));
  INV_X1    g492(.A(new_n300), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n695), .B(new_n453), .C1(new_n471), .C2(new_n483), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n634), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n570), .ZN(new_n698));
  INV_X1    g497(.A(new_n600), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .A4(new_n666), .ZN(new_n700));
  INV_X1    g499(.A(new_n673), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n700), .A2(G29gat), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT45), .Z(new_n703));
  INV_X1    g502(.A(new_n562), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n704), .A3(new_n666), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n697), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n634), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n485), .B2(new_n496), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n708), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n705), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n701), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n703), .A2(new_n717), .ZN(G1328gat));
  INV_X1    g517(.A(new_n472), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n700), .A2(new_n719), .A3(new_n521), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT46), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n521), .B1(new_n716), .B2(new_n719), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n683), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n700), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT47), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n724), .B1(new_n715), .B2(new_n305), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n729), .A2(new_n730), .A3(new_n726), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n726), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1330gat));
  NAND3_X1  g532(.A1(new_n715), .A2(G50gat), .A3(new_n369), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n700), .A2(new_n368), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(G50gat), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g536(.A1(new_n637), .A2(new_n562), .A3(new_n638), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n497), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n701), .A2(new_n666), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  INV_X1    g541(.A(new_n666), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n719), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  OAI21_X1  g548(.A(G71gat), .B1(new_n744), .B2(new_n695), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n683), .A2(new_n572), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n744), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g552(.A1(new_n744), .A2(new_n368), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n573), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n704), .A2(new_n600), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n666), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n711), .B2(new_n714), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n701), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n712), .B(new_n756), .C1(new_n485), .C2(new_n496), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n697), .A2(KEYINPUT106), .A3(KEYINPUT51), .A4(new_n756), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n397), .A3(new_n740), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n762), .A2(new_n771), .ZN(G1336gat));
  NOR3_X1   g571(.A1(new_n719), .A2(G92gat), .A3(new_n666), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  INV_X1    g574(.A(new_n710), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n708), .B1(new_n713), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n692), .A2(new_n696), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n709), .B1(new_n778), .B2(new_n712), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n472), .B(new_n758), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n774), .A2(new_n775), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n774), .A2(KEYINPUT108), .A3(new_n775), .A4(new_n781), .ZN(new_n785));
  INV_X1    g584(.A(new_n781), .ZN(new_n786));
  INV_X1    g585(.A(new_n773), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n769), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n764), .A2(KEYINPUT107), .A3(new_n765), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n787), .B1(new_n791), .B2(new_n768), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT52), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n784), .A2(new_n785), .A3(new_n793), .ZN(G1337gat));
  NAND3_X1  g593(.A1(new_n760), .A2(KEYINPUT109), .A3(new_n305), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G99gat), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT109), .B1(new_n760), .B2(new_n305), .ZN(new_n797));
  INV_X1    g596(.A(new_n770), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n304), .A2(G99gat), .A3(new_n666), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n796), .A2(new_n797), .B1(new_n798), .B2(new_n799), .ZN(G1338gat));
  OAI211_X1 g599(.A(new_n369), .B(new_n758), .C1(new_n777), .C2(new_n779), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT53), .B1(new_n801), .B2(G106gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n368), .A2(G106gat), .A3(new_n666), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n801), .A2(KEYINPUT110), .A3(G106gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n791), .B2(new_n768), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT110), .B1(new_n801), .B2(G106gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(G1339gat));
  NOR2_X1   g610(.A1(new_n738), .A2(new_n743), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n660), .A2(new_n639), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n813), .A2(new_n652), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI211_X1 g615(.A(KEYINPUT101), .B(new_n640), .C1(new_n649), .C2(new_n651), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n663), .B1(new_n660), .B2(new_n639), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n819), .A2(new_n820), .A3(new_n655), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n819), .B2(new_n655), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT55), .B(new_n816), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n656), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT54), .B1(new_n662), .B2(new_n664), .ZN(new_n826));
  INV_X1    g625(.A(new_n655), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT111), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n819), .A2(new_n820), .A3(new_n655), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT55), .B1(new_n830), .B2(new_n816), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n825), .A2(new_n831), .A3(new_n562), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n533), .A2(new_n534), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n540), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n549), .B1(new_n509), .B2(new_n519), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT112), .B(new_n543), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n541), .A2(new_n550), .A3(new_n552), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n535), .A2(new_n541), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT112), .B1(new_n839), .B2(new_n543), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n560), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n567), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n743), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n567), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT113), .B1(new_n845), .B2(new_n666), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n634), .B1(new_n832), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n825), .A2(new_n831), .A3(new_n634), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n842), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n600), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(KEYINPUT114), .A3(new_n850), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n812), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n701), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n489), .A2(new_n490), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n719), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n258), .B1(new_n859), .B2(new_n562), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(new_n704), .A3(new_n824), .A4(new_n823), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n844), .A2(new_n846), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n712), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR4_X1   g665(.A1(new_n825), .A2(new_n831), .A3(new_n634), .A4(new_n845), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n852), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n854), .A2(new_n699), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n812), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n701), .A2(new_n472), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n871), .A2(new_n494), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(G113gat), .A3(new_n698), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n860), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT115), .ZN(G1340gat));
  INV_X1    g675(.A(new_n859), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n255), .A3(new_n743), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n873), .A2(new_n743), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n255), .B2(new_n879), .ZN(G1341gat));
  AOI21_X1  g679(.A(G127gat), .B1(new_n877), .B2(new_n600), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n600), .A2(G127gat), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n873), .B2(new_n882), .ZN(G1342gat));
  NAND2_X1  g682(.A1(new_n873), .A2(new_n712), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(G134gat), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n859), .A2(G134gat), .A3(new_n634), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n886), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(G1343gat));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n845), .A2(new_n666), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n815), .B1(new_n828), .B2(new_n829), .ZN(new_n895));
  XNOR2_X1  g694(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n823), .B(new_n824), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n570), .B1(new_n898), .B2(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n861), .A2(new_n896), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n824), .A4(new_n823), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n894), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n850), .B1(new_n903), .B2(new_n712), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n812), .B1(new_n904), .B2(new_n699), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT57), .B1(new_n905), .B2(new_n368), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n871), .A2(new_n907), .A3(new_n369), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n872), .B2(new_n695), .ZN(new_n910));
  NOR4_X1   g709(.A1(new_n701), .A2(new_n305), .A3(KEYINPUT117), .A4(new_n472), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n906), .A2(new_n908), .A3(new_n704), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G141gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n695), .A2(new_n369), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n719), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n916), .B2(new_n915), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n570), .A2(G141gat), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n918), .A2(new_n673), .A3(new_n871), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n893), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n893), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n908), .A3(new_n698), .A4(new_n912), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(G141gat), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT121), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(G141gat), .ZN(new_n926));
  INV_X1    g725(.A(new_n922), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n918), .A2(new_n673), .A3(new_n871), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n913), .A2(G141gat), .B1(new_n930), .B2(new_n919), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n928), .B(new_n929), .C1(new_n893), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n925), .A2(new_n932), .ZN(G1344gat));
  INV_X1    g732(.A(G148gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n934), .A3(new_n743), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT57), .B1(new_n855), .B2(new_n368), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n903), .A2(new_n712), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n845), .B1(new_n849), .B2(KEYINPUT122), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(KEYINPUT122), .B2(new_n849), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n600), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n667), .A2(new_n698), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n907), .B(new_n369), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n743), .A3(new_n912), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n936), .B1(new_n945), .B2(G148gat), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n906), .A2(new_n908), .A3(new_n912), .ZN(new_n947));
  AOI211_X1 g746(.A(KEYINPUT59), .B(new_n934), .C1(new_n947), .C2(new_n743), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n935), .B1(new_n946), .B2(new_n948), .ZN(G1345gat));
  AOI21_X1  g748(.A(G155gat), .B1(new_n930), .B2(new_n600), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n699), .A2(new_n320), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n947), .B2(new_n951), .ZN(G1346gat));
  NAND3_X1  g751(.A1(new_n930), .A2(new_n321), .A3(new_n712), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n947), .A2(new_n712), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n321), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n673), .A2(new_n719), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n871), .A2(new_n494), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n871), .A2(KEYINPUT125), .A3(new_n494), .A4(new_n956), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n698), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G169gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n673), .B1(new_n869), .B2(new_n870), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n719), .B1(new_n964), .B2(KEYINPUT123), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n966), .B1(new_n855), .B2(new_n673), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n562), .A2(G169gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n857), .A3(new_n969), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(G1348gat));
  AND2_X1   g772(.A1(new_n968), .A2(new_n857), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n743), .ZN(new_n975));
  INV_X1    g774(.A(G176gat), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n666), .A2(new_n976), .ZN(new_n977));
  AOI22_X1  g776(.A1(new_n975), .A2(new_n976), .B1(new_n961), .B2(new_n977), .ZN(G1349gat));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT60), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n959), .A2(new_n600), .A3(new_n960), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G183gat), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n600), .A2(new_n202), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n967), .A3(new_n857), .A4(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n979), .A2(new_n980), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  AND4_X1   g786(.A1(new_n981), .A2(new_n983), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n986), .B1(new_n982), .B2(G183gat), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n981), .B1(new_n989), .B2(new_n985), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n988), .A2(new_n990), .ZN(G1350gat));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n209), .A3(new_n712), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n959), .A2(new_n712), .A3(new_n960), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n993), .B1(new_n994), .B2(G190gat), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n994), .A2(new_n993), .A3(G190gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G1351gat));
  INV_X1    g796(.A(new_n915), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n968), .A2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(G197gat), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n999), .A2(new_n1000), .A3(new_n704), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n956), .A2(new_n695), .ZN(new_n1002));
  INV_X1    g801(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n937), .A2(new_n943), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g803(.A(G197gat), .B1(new_n1004), .B2(new_n570), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1001), .A2(new_n1005), .ZN(G1352gat));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n666), .A2(G204gat), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n965), .A2(new_n967), .A3(new_n998), .A4(new_n1008), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n1009), .A2(KEYINPUT127), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1009), .A2(KEYINPUT127), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n944), .A2(new_n743), .A3(new_n1003), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(G204gat), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n968), .A2(new_n1015), .A3(new_n998), .A4(new_n1008), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1009), .A2(KEYINPUT127), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n1016), .A2(KEYINPUT62), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1012), .A2(new_n1014), .A3(new_n1018), .ZN(G1353gat));
  NAND3_X1  g818(.A1(new_n999), .A2(new_n310), .A3(new_n600), .ZN(new_n1020));
  NAND4_X1  g819(.A1(new_n937), .A2(new_n943), .A3(new_n600), .A4(new_n1003), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1021), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g822(.A(KEYINPUT63), .B1(new_n1021), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(G1354gat));
  NOR3_X1   g824(.A1(new_n1004), .A2(new_n311), .A3(new_n634), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n999), .A2(new_n712), .ZN(new_n1027));
  AOI21_X1  g826(.A(new_n1026), .B1(new_n1027), .B2(new_n311), .ZN(G1355gat));
endmodule


