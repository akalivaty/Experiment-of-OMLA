//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT79), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT79), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n206), .A3(G141gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n203), .A2(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT80), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT80), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(KEYINPUT2), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n210), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n203), .A2(G141gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n212), .B1(new_n223), .B2(new_n208), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n220), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT3), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n220), .B1(new_n207), .B2(new_n209), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n228), .A2(new_n218), .B1(new_n220), .B2(new_n224), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(G127gat), .B(G134gat), .Z(new_n233));
  INV_X1    g032(.A(G113gat), .ZN(new_n234));
  INV_X1    g033(.A(G120gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G113gat), .A2(G120gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n233), .A2(new_n238), .A3(KEYINPUT1), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240));
  AND2_X1   g039(.A1(G113gat), .A2(G120gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(G113gat), .A2(G120gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(KEYINPUT67), .A3(new_n237), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n233), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT68), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n249), .A3(new_n233), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n239), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT81), .B1(new_n232), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n239), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n246), .A2(new_n249), .A3(new_n233), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n249), .B1(new_n246), .B2(new_n233), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n227), .A4(new_n231), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n251), .A2(new_n260), .A3(new_n229), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n253), .B(new_n229), .C1(new_n254), .C2(new_n255), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n202), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT94), .B(KEYINPUT39), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT0), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G85gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT39), .ZN(new_n274));
  INV_X1    g073(.A(new_n202), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n226), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n262), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n256), .A2(KEYINPUT83), .A3(new_n226), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n265), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT40), .ZN(new_n282));
  OR3_X1    g081(.A1(new_n273), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n273), .B2(new_n281), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT82), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n262), .B2(KEYINPUT4), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n251), .A2(KEYINPUT82), .A3(new_n260), .A4(new_n229), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n263), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n259), .A2(new_n288), .A3(new_n202), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n278), .A2(new_n275), .A3(new_n279), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(KEYINPUT5), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n275), .B1(new_n252), .B2(new_n258), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT5), .B1(new_n261), .B2(new_n263), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n272), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n283), .A2(new_n284), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  INV_X1    g103(.A(G190gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G169gat), .ZN(new_n307));
  INV_X1    g106(.A(G176gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT65), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n306), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI211_X1 g118(.A(KEYINPUT66), .B(new_n306), .C1(new_n313), .C2(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n304), .A2(KEYINPUT27), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT27), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G183gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n323), .A3(new_n305), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT28), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT27), .B(G183gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(new_n305), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n319), .A2(new_n320), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n333), .A2(KEYINPUT64), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(KEYINPUT64), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n305), .A2(G183gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n304), .A2(G190gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT24), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT24), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n306), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n336), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT23), .ZN(new_n343));
  INV_X1    g142(.A(new_n315), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT25), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n344), .B1(KEYINPUT23), .B2(new_n331), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n336), .A2(new_n339), .A3(new_n348), .A4(new_n341), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n342), .A2(new_n347), .B1(new_n349), .B2(new_n345), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n303), .B1(new_n330), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n313), .A2(new_n316), .ZN(new_n354));
  INV_X1    g153(.A(new_n306), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT66), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n317), .A2(new_n318), .ZN(new_n358));
  INV_X1    g157(.A(new_n329), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n347), .A2(new_n339), .A3(new_n341), .A4(new_n336), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n349), .A2(new_n345), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n353), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n351), .B1(new_n364), .B2(new_n303), .ZN(new_n365));
  INV_X1    g164(.A(G211gat), .ZN(new_n366));
  INV_X1    g165(.A(G218gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G211gat), .A2(G218gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT74), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n372), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT22), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT73), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT73), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n369), .A2(new_n378), .A3(new_n375), .ZN(new_n379));
  XNOR2_X1  g178(.A(G197gat), .B(G204gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n380), .A2(new_n379), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n383), .A2(new_n371), .A3(new_n373), .A4(new_n377), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n384), .A3(KEYINPUT75), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT75), .B1(new_n382), .B2(new_n384), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n365), .A2(KEYINPUT77), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT77), .B1(new_n365), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n386), .A2(new_n387), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n360), .B2(new_n363), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n351), .B(new_n392), .C1(new_n393), .C2(new_n303), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT78), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n320), .A2(new_n329), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n396), .A2(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n302), .B1(new_n397), .B2(KEYINPUT29), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n351), .A4(new_n392), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n301), .B1(new_n391), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n302), .B1(new_n360), .B2(new_n363), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n352), .B1(new_n330), .B2(new_n350), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n404), .B1(new_n405), .B2(new_n302), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n406), .B2(new_n392), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n365), .A2(KEYINPUT77), .A3(new_n388), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n407), .A2(new_n408), .B1(new_n395), .B2(new_n400), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n300), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n412), .A3(new_n300), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n411), .A2(KEYINPUT93), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT93), .B1(new_n411), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n297), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G78gat), .B(G106gat), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT87), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT31), .B(G50gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G22gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(G228gat), .A2(G233gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n231), .A2(new_n352), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n382), .A2(new_n384), .A3(new_n352), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n229), .B1(new_n425), .B2(new_n230), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT88), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n392), .A2(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n426), .A2(new_n427), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n422), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n382), .A2(new_n384), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n230), .B1(new_n431), .B2(KEYINPUT29), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n226), .ZN(new_n433));
  INV_X1    g232(.A(new_n422), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n433), .B(new_n434), .C1(new_n392), .C2(new_n424), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n421), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n430), .A2(new_n421), .A3(new_n435), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(KEYINPUT89), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(KEYINPUT89), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n420), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n430), .A2(new_n435), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT90), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT90), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n430), .A2(new_n444), .A3(new_n435), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(G22gat), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n430), .A2(KEYINPUT91), .A3(new_n421), .A4(new_n435), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n447), .A2(new_n420), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT91), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n437), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n441), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n295), .A2(KEYINPUT6), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n271), .B1(new_n292), .B2(new_n293), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n259), .A2(new_n288), .A3(new_n202), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n454), .B(new_n455), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n455), .B1(new_n291), .B2(new_n454), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n453), .B1(new_n462), .B2(new_n296), .ZN(new_n463));
  XOR2_X1   g262(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n464));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n365), .B2(new_n392), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n398), .A2(new_n351), .A3(new_n388), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n407), .A2(new_n408), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n395), .A2(new_n400), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n301), .B(new_n468), .C1(new_n471), .C2(KEYINPUT37), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT96), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n300), .B1(new_n469), .B2(new_n470), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n300), .A2(new_n465), .ZN(new_n476));
  OAI211_X1 g275(.A(KEYINPUT96), .B(new_n468), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n475), .A2(new_n476), .B1(new_n465), .B2(new_n409), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n479), .A2(new_n464), .B1(new_n300), .B2(new_n409), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n416), .A2(new_n452), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G227gat), .ZN(new_n483));
  INV_X1    g282(.A(G233gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n251), .A2(KEYINPUT69), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT69), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n256), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n360), .A2(new_n363), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n397), .A2(new_n487), .A3(new_n256), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n485), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g293(.A(KEYINPUT34), .B(new_n485), .C1(new_n490), .C2(new_n491), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n485), .A3(new_n491), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT32), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G15gat), .B(G43gat), .Z(new_n501));
  XNOR2_X1  g300(.A(G71gat), .B(G99gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n503), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n497), .B(KEYINPUT32), .C1(new_n499), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n504), .B2(new_n506), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n496), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT71), .B(new_n496), .C1(new_n508), .C2(new_n510), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n507), .A2(new_n496), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n513), .A2(KEYINPUT36), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n494), .A2(new_n495), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n504), .B2(new_n506), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n411), .A2(new_n413), .ZN(new_n525));
  INV_X1    g324(.A(new_n461), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n458), .A2(new_n459), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n295), .A2(new_n528), .ZN(new_n529));
  AOI211_X1 g328(.A(KEYINPUT85), .B(new_n272), .C1(new_n291), .C2(new_n294), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n526), .B(new_n527), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n453), .B1(new_n531), .B2(KEYINPUT86), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n462), .B(new_n533), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n525), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n452), .A2(KEYINPUT92), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n537));
  OR3_X1    g336(.A1(new_n537), .A2(new_n440), .A3(KEYINPUT92), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n482), .B(new_n524), .C1(new_n535), .C2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n520), .B1(new_n537), .B2(new_n440), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(new_n463), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n414), .A2(new_n415), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT35), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AND4_X1   g344(.A1(new_n514), .A2(new_n452), .A3(new_n516), .A4(new_n513), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n535), .A3(KEYINPUT35), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G43gat), .B(G50gat), .Z(new_n549));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT97), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(KEYINPUT15), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT98), .B(KEYINPUT15), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n549), .A2(new_n555), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NOR3_X1   g357(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT99), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n554), .B(new_n556), .C1(new_n558), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G29gat), .A2(G36gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n558), .B2(new_n559), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n551), .A2(KEYINPUT15), .A3(new_n563), .A4(new_n553), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT17), .ZN(new_n567));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT16), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(G1gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(G1gat), .B2(new_n568), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G8gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n565), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n567), .A2(new_n574), .B1(new_n565), .B2(new_n572), .ZN(new_n575));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n577), .A2(KEYINPUT18), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(KEYINPUT18), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n565), .B(new_n572), .Z(new_n580));
  XOR2_X1   g379(.A(new_n576), .B(KEYINPUT13), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G197gat), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT11), .B(G169gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT12), .Z(new_n589));
  OR2_X1    g388(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT100), .ZN(new_n593));
  XOR2_X1   g392(.A(G134gat), .B(G162gat), .Z(new_n594));
  AOI21_X1  g393(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT102), .Z(new_n597));
  NAND3_X1  g396(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(G85gat), .ZN(new_n600));
  INV_X1    g399(.A(G92gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(KEYINPUT8), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT103), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G99gat), .B(G106gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n598), .B1(new_n609), .B2(new_n566), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT104), .ZN(new_n611));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT105), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n565), .A2(new_n573), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n567), .A2(new_n615), .A3(new_n609), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT106), .Z(new_n618));
  AOI21_X1  g417(.A(new_n614), .B1(new_n611), .B2(new_n616), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT107), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n597), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT101), .A2(G57gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G64gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(G71gat), .A2(G78gat), .ZN(new_n626));
  OR2_X1    g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT9), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n631));
  AND2_X1   g430(.A1(G57gat), .A2(G64gat), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n626), .B(new_n627), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n609), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT108), .B1(new_n609), .B2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT108), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n609), .A2(new_n638), .A3(new_n634), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT10), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n623), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n623), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n637), .A2(new_n644), .A3(new_n639), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n643), .A2(new_n645), .A3(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT21), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n634), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(G127gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n572), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n655), .B2(new_n634), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G155gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(G183gat), .B(G211gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n663), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n617), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n596), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n620), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n622), .A2(new_n654), .A3(new_n668), .A4(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n548), .A2(new_n593), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT109), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n592), .B(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT35), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n678), .B(new_n525), .C1(new_n532), .C2(new_n534), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n544), .B1(new_n679), .B2(new_n546), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n677), .B1(new_n680), .B2(new_n540), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n673), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n532), .A2(new_n534), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  INV_X1    g487(.A(new_n543), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AND3_X1   g489(.A1(new_n684), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(G8gat), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n692), .B1(new_n684), .B2(new_n689), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT42), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(KEYINPUT42), .B2(new_n691), .ZN(G1325gat));
  INV_X1    g494(.A(G15gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n684), .A2(new_n696), .A3(new_n520), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n524), .B1(new_n675), .B2(new_n683), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n698), .B2(new_n696), .ZN(G1326gat));
  INV_X1    g498(.A(new_n539), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT110), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n684), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n702), .B2(new_n704), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(new_n671), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n621), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n668), .A3(new_n653), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n685), .A2(G29gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n681), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n622), .A2(KEYINPUT113), .A3(new_n671), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n621), .B2(new_n709), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n548), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n710), .B1(new_n680), .B2(new_n540), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n718), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n653), .B(KEYINPUT111), .Z(new_n724));
  INV_X1    g523(.A(new_n668), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n592), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT112), .Z(new_n727));
  NAND3_X1  g526(.A1(new_n723), .A2(new_n686), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G29gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1328gat));
  AND2_X1   g531(.A1(new_n681), .A2(new_n711), .ZN(new_n733));
  INV_X1    g532(.A(G36gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n689), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT46), .Z(new_n736));
  AND2_X1   g535(.A1(new_n723), .A2(new_n727), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n689), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n739), .B2(new_n734), .ZN(G1329gat));
  INV_X1    g539(.A(G43gat), .ZN(new_n741));
  INV_X1    g540(.A(new_n524), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n742), .A3(new_n727), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n723), .A2(KEYINPUT115), .A3(new_n742), .A4(new_n727), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n733), .A2(new_n741), .A3(new_n520), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(G43gat), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(new_n748), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n747), .A2(new_n749), .B1(new_n751), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g551(.A(G50gat), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n733), .A2(new_n753), .A3(new_n700), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n700), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(G50gat), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n452), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n753), .B1(new_n737), .B2(new_n759), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n756), .A2(KEYINPUT48), .B1(new_n758), .B2(new_n760), .ZN(G1331gat));
  INV_X1    g560(.A(new_n592), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n621), .A2(new_n709), .A3(new_n725), .ZN(new_n763));
  INV_X1    g562(.A(new_n724), .ZN(new_n764));
  AND4_X1   g563(.A1(new_n548), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n686), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT116), .B(G57gat), .Z(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1332gat));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n689), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT49), .B(G64gat), .Z(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(G1333gat));
  NAND2_X1  g571(.A1(new_n765), .A2(new_n742), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n521), .A2(G71gat), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n773), .A2(G71gat), .B1(new_n765), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n765), .A2(new_n700), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g577(.A1(new_n592), .A2(new_n654), .A3(new_n668), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n723), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n686), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G85gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n592), .A2(new_n668), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT51), .B1(new_n722), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT117), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n622), .A2(new_n671), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n548), .A2(new_n787), .A3(new_n783), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n786), .B1(new_n790), .B2(new_n785), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n686), .A2(new_n600), .A3(new_n653), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n782), .B1(new_n791), .B2(new_n792), .ZN(G1336gat));
  NOR3_X1   g592(.A1(new_n724), .A2(G92gat), .A3(new_n543), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n723), .A2(new_n689), .A3(new_n779), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(new_n601), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n790), .A2(new_n794), .B1(new_n798), .B2(G92gat), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n796), .A2(new_n800), .B1(new_n797), .B2(new_n801), .ZN(G1337gat));
  NAND2_X1  g601(.A1(new_n780), .A2(new_n742), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G99gat), .ZN(new_n804));
  OR3_X1    g603(.A1(new_n654), .A2(new_n521), .A3(G99gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n791), .B2(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n724), .A2(G106gat), .A3(new_n452), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n786), .B(new_n807), .C1(new_n790), .C2(new_n785), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n723), .A2(new_n759), .A3(new_n779), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT53), .B1(new_n809), .B2(G106gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n718), .B1(new_n548), .B2(new_n787), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n719), .B1(new_n680), .B2(new_n540), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n700), .B(new_n779), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n788), .A2(new_n789), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n807), .B1(new_n816), .B2(new_n784), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n818), .B2(KEYINPUT53), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n820), .B(new_n821), .C1(new_n815), .C2(new_n817), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n811), .B1(new_n819), .B2(new_n822), .ZN(G1339gat));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n672), .B2(new_n592), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n763), .A2(KEYINPUT119), .A3(new_n762), .A4(new_n654), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n715), .A2(new_n717), .ZN(new_n828));
  INV_X1    g627(.A(new_n643), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n649), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n640), .A2(new_n623), .A3(new_n642), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(KEYINPUT54), .A3(new_n643), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n652), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n833), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n592), .A3(new_n838), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n575), .A2(new_n576), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n840), .A2(KEYINPUT120), .B1(new_n580), .B2(new_n582), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(KEYINPUT120), .B2(new_n840), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n588), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n590), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n654), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n844), .B(KEYINPUT121), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n838), .A2(new_n652), .A3(new_n834), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n715), .A3(new_n717), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n827), .B1(new_n852), .B2(new_n725), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n685), .A2(new_n689), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n700), .A2(new_n521), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(new_n234), .A3(new_n677), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n853), .A2(new_n685), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n859), .A2(new_n543), .A3(new_n546), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n592), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n858), .B1(new_n861), .B2(new_n234), .ZN(G1340gat));
  NOR3_X1   g661(.A1(new_n857), .A2(new_n235), .A3(new_n724), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n653), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n235), .ZN(G1341gat));
  NOR2_X1   g664(.A1(new_n725), .A2(new_n659), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OR3_X1    g666(.A1(new_n857), .A2(KEYINPUT122), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT122), .B1(new_n857), .B2(new_n867), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(G127gat), .B1(new_n860), .B2(new_n668), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n710), .A2(new_n689), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n873), .A3(new_n546), .A4(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n857), .B2(new_n710), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G1343gat));
  AOI21_X1  g678(.A(new_n845), .B1(new_n593), .B2(new_n850), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n851), .B1(new_n880), .B2(new_n787), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n827), .B1(new_n881), .B2(new_n725), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT57), .B1(new_n882), .B2(new_n539), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n668), .B1(new_n848), .B2(new_n851), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n884), .B(new_n759), .C1(new_n885), .C2(new_n827), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n855), .A2(new_n524), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n883), .A2(new_n593), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G141gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n742), .A2(new_n452), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n686), .B(new_n890), .C1(new_n885), .C2(new_n827), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n689), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n677), .A2(G141gat), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT58), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n883), .A2(new_n592), .A3(new_n886), .A4(new_n887), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n896), .A2(G141gat), .B1(new_n892), .B2(new_n893), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n204), .A2(new_n206), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n654), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT57), .B1(new_n853), .B2(new_n452), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n835), .A2(new_n838), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n846), .B1(new_n677), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n710), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT123), .B1(new_n906), .B2(new_n710), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n787), .A2(new_n850), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n911), .A3(new_n849), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n668), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n593), .A2(new_n672), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n884), .B(new_n700), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n905), .A2(new_n915), .A3(new_n653), .A4(new_n887), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n903), .A2(new_n203), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n654), .A2(new_n900), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n916), .A2(new_n917), .B1(new_n892), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n901), .B2(new_n725), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n892), .A2(new_n215), .A3(new_n668), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n901), .B2(new_n828), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n874), .A2(new_n216), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n891), .B2(new_n925), .ZN(G1347gat));
  AND2_X1   g725(.A1(new_n546), .A2(new_n689), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n854), .A2(new_n685), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n307), .B1(new_n928), .B2(new_n762), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n686), .A2(new_n543), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n677), .A2(new_n307), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n854), .A2(new_n856), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n929), .A2(KEYINPUT124), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1348gat));
  NAND3_X1  g736(.A1(new_n854), .A2(new_n856), .A3(new_n930), .ZN(new_n938));
  OAI21_X1  g737(.A(G176gat), .B1(new_n938), .B2(new_n724), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n653), .A2(new_n308), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n928), .B2(new_n940), .ZN(G1349gat));
  OAI21_X1  g740(.A(G183gat), .B1(new_n938), .B2(new_n725), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n853), .A2(new_n686), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n943), .A2(new_n326), .A3(new_n668), .A4(new_n927), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT60), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n942), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1350gat));
  NAND4_X1  g748(.A1(new_n854), .A2(new_n787), .A3(new_n856), .A4(new_n930), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n951), .A3(G190gat), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n950), .B2(G190gat), .ZN(new_n954));
  INV_X1    g753(.A(new_n828), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n305), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n953), .A2(new_n954), .B1(new_n928), .B2(new_n956), .ZN(G1351gat));
  NAND2_X1  g756(.A1(new_n890), .A2(new_n689), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n943), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n592), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n905), .A2(new_n915), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n930), .A2(new_n524), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT126), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n593), .A2(G197gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n962), .B1(new_n967), .B2(new_n968), .ZN(G1352gat));
  NAND4_X1  g768(.A1(new_n905), .A2(new_n915), .A3(new_n764), .A4(new_n965), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n654), .A2(G204gat), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n943), .A2(new_n959), .A3(new_n960), .A4(new_n971), .ZN(new_n972));
  AOI22_X1  g771(.A1(new_n970), .A2(G204gat), .B1(new_n972), .B2(KEYINPUT62), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  INV_X1    g773(.A(new_n972), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n972), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n961), .A2(new_n366), .A3(new_n668), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n905), .A2(new_n915), .A3(new_n668), .A4(new_n965), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  OAI21_X1  g783(.A(G218gat), .B1(new_n966), .B2(new_n710), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n961), .A2(new_n367), .A3(new_n955), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


