

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  INV_X1 U322 ( .A(KEYINPUT90), .ZN(n446) );
  XNOR2_X1 U323 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n416) );
  XNOR2_X1 U324 ( .A(n477), .B(KEYINPUT37), .ZN(n478) );
  XNOR2_X1 U325 ( .A(n346), .B(n345), .ZN(n351) );
  INV_X1 U326 ( .A(KEYINPUT54), .ZN(n430) );
  XNOR2_X1 U327 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n407) );
  XNOR2_X1 U328 ( .A(n430), .B(KEYINPUT120), .ZN(n431) );
  XNOR2_X1 U329 ( .A(n408), .B(n407), .ZN(n415) );
  XNOR2_X1 U330 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U331 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U332 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U333 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U334 ( .A(n454), .B(KEYINPUT121), .ZN(n455) );
  XNOR2_X1 U335 ( .A(n452), .B(n423), .ZN(n350) );
  XNOR2_X1 U336 ( .A(n351), .B(n350), .ZN(n411) );
  XNOR2_X1 U337 ( .A(n479), .B(n478), .ZN(n519) );
  XOR2_X1 U338 ( .A(n411), .B(n352), .Z(n565) );
  INV_X1 U339 ( .A(G43GAT), .ZN(n481) );
  XNOR2_X1 U340 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U341 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U342 ( .A(n484), .B(n483), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT67), .B(KEYINPUT85), .Z(n291) );
  XNOR2_X1 U344 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n290) );
  XNOR2_X1 U345 ( .A(n291), .B(n290), .ZN(n307) );
  XOR2_X1 U346 ( .A(KEYINPUT88), .B(G190GAT), .Z(n293) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G99GAT), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U349 ( .A(n294), .B(G176GAT), .Z(n296) );
  XOR2_X1 U350 ( .A(G134GAT), .B(KEYINPUT0), .Z(n324) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(n324), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G127GAT), .Z(n371) );
  XOR2_X1 U354 ( .A(n371), .B(KEYINPUT20), .Z(n298) );
  NAND2_X1 U355 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U356 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U357 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U358 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n302) );
  XNOR2_X1 U359 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U361 ( .A(G169GAT), .B(n303), .Z(n426) );
  XOR2_X1 U362 ( .A(G120GAT), .B(G71GAT), .Z(n329) );
  XNOR2_X1 U363 ( .A(n426), .B(n329), .ZN(n304) );
  XNOR2_X1 U364 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U365 ( .A(n307), .B(n306), .Z(n472) );
  XOR2_X1 U366 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n309) );
  XNOR2_X1 U367 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n328) );
  XOR2_X1 U369 ( .A(G85GAT), .B(G162GAT), .Z(n311) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U372 ( .A(KEYINPUT1), .B(G155GAT), .Z(n313) );
  XNOR2_X1 U373 ( .A(G127GAT), .B(G148GAT), .ZN(n312) );
  XNOR2_X1 U374 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U375 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U376 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n317) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U379 ( .A(KEYINPUT92), .B(n318), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n323) );
  XOR2_X1 U381 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n322) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(KEYINPUT91), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n451) );
  XOR2_X1 U384 ( .A(n323), .B(n451), .Z(n326) );
  XOR2_X1 U385 ( .A(G113GAT), .B(G1GAT), .Z(n355) );
  XNOR2_X1 U386 ( .A(n355), .B(n324), .ZN(n325) );
  XNOR2_X1 U387 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U388 ( .A(n328), .B(n327), .Z(n520) );
  XOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT13), .Z(n383) );
  XNOR2_X1 U390 ( .A(n329), .B(n383), .ZN(n331) );
  XOR2_X1 U391 ( .A(KEYINPUT33), .B(G92GAT), .Z(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U393 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n333) );
  XNOR2_X1 U394 ( .A(KEYINPUT77), .B(KEYINPUT74), .ZN(n332) );
  XOR2_X1 U395 ( .A(n333), .B(n332), .Z(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n339) );
  INV_X1 U397 ( .A(n339), .ZN(n337) );
  NAND2_X1 U398 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  INV_X1 U399 ( .A(n338), .ZN(n336) );
  NAND2_X1 U400 ( .A1(n337), .A2(n336), .ZN(n341) );
  NAND2_X1 U401 ( .A1(n339), .A2(n338), .ZN(n340) );
  NAND2_X1 U402 ( .A1(n341), .A2(n340), .ZN(n346) );
  XNOR2_X1 U403 ( .A(G99GAT), .B(G106GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n342), .B(G85GAT), .ZN(n392) );
  XNOR2_X1 U405 ( .A(n392), .B(KEYINPUT31), .ZN(n344) );
  INV_X1 U406 ( .A(KEYINPUT73), .ZN(n343) );
  XOR2_X1 U407 ( .A(G78GAT), .B(KEYINPUT75), .Z(n347) );
  XNOR2_X1 U408 ( .A(G148GAT), .B(n347), .ZN(n452) );
  XOR2_X1 U409 ( .A(KEYINPUT76), .B(G64GAT), .Z(n349) );
  XNOR2_X1 U410 ( .A(G176GAT), .B(G204GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n423) );
  XNOR2_X1 U412 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n352) );
  INV_X1 U413 ( .A(n565), .ZN(n551) );
  XOR2_X1 U414 ( .A(G29GAT), .B(G43GAT), .Z(n354) );
  XNOR2_X1 U415 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n401) );
  XOR2_X1 U417 ( .A(n401), .B(n355), .Z(n357) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U420 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n359) );
  XNOR2_X1 U421 ( .A(KEYINPUT70), .B(KEYINPUT30), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U423 ( .A(n361), .B(n360), .Z(n369) );
  XOR2_X1 U424 ( .A(G15GAT), .B(G50GAT), .Z(n363) );
  XNOR2_X1 U425 ( .A(G169GAT), .B(G36GAT), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U427 ( .A(G8GAT), .B(G22GAT), .Z(n365) );
  XNOR2_X1 U428 ( .A(G197GAT), .B(G141GAT), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n573) );
  NOR2_X1 U432 ( .A1(n551), .A2(n573), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n370), .B(KEYINPUT46), .ZN(n390) );
  XOR2_X1 U434 ( .A(n371), .B(KEYINPUT83), .Z(n373) );
  NAND2_X1 U435 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U437 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n375) );
  XNOR2_X1 U438 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U441 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n379) );
  XNOR2_X1 U442 ( .A(G1GAT), .B(KEYINPUT81), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U444 ( .A(G8GAT), .B(n380), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n387) );
  XOR2_X1 U446 ( .A(G22GAT), .B(G155GAT), .Z(n439) );
  XOR2_X1 U447 ( .A(n383), .B(n439), .Z(n385) );
  XNOR2_X1 U448 ( .A(G78GAT), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U450 ( .A(n387), .B(n386), .Z(n389) );
  XNOR2_X1 U451 ( .A(G183GAT), .B(G71GAT), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n568) );
  NOR2_X1 U453 ( .A1(n390), .A2(n568), .ZN(n406) );
  XOR2_X1 U454 ( .A(G50GAT), .B(G162GAT), .Z(n438) );
  XNOR2_X1 U455 ( .A(n438), .B(KEYINPUT68), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n391), .B(KEYINPUT11), .ZN(n405) );
  XOR2_X1 U457 ( .A(n392), .B(KEYINPUT10), .Z(n394) );
  NAND2_X1 U458 ( .A1(G232GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U460 ( .A(KEYINPUT78), .B(KEYINPUT69), .Z(n396) );
  XNOR2_X1 U461 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U463 ( .A(n398), .B(n397), .Z(n403) );
  XOR2_X1 U464 ( .A(G92GAT), .B(G218GAT), .Z(n400) );
  XNOR2_X1 U465 ( .A(G36GAT), .B(G190GAT), .ZN(n399) );
  XNOR2_X1 U466 ( .A(n400), .B(n399), .ZN(n420) );
  XNOR2_X1 U467 ( .A(n401), .B(n420), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n557) );
  NAND2_X1 U470 ( .A1(n406), .A2(n557), .ZN(n408) );
  XNOR2_X1 U471 ( .A(KEYINPUT79), .B(n557), .ZN(n541) );
  INV_X1 U472 ( .A(n541), .ZN(n485) );
  XNOR2_X1 U473 ( .A(KEYINPUT36), .B(n485), .ZN(n585) );
  INV_X1 U474 ( .A(n568), .ZN(n582) );
  NOR2_X1 U475 ( .A1(n585), .A2(n582), .ZN(n409) );
  XNOR2_X1 U476 ( .A(KEYINPUT45), .B(n409), .ZN(n410) );
  NAND2_X1 U477 ( .A1(n410), .A2(n573), .ZN(n413) );
  INV_X1 U478 ( .A(n411), .ZN(n412) );
  NOR2_X1 U479 ( .A1(n413), .A2(n412), .ZN(n414) );
  NOR2_X1 U480 ( .A1(n415), .A2(n414), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n532) );
  XOR2_X1 U482 ( .A(G8GAT), .B(KEYINPUT95), .Z(n419) );
  NAND2_X1 U483 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U485 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U486 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n422), .B(G211GAT), .ZN(n445) );
  XNOR2_X1 U488 ( .A(n445), .B(n423), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n428) );
  INV_X1 U490 ( .A(n426), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n524) );
  XNOR2_X1 U492 ( .A(n524), .B(KEYINPUT119), .ZN(n429) );
  NOR2_X1 U493 ( .A1(n532), .A2(n429), .ZN(n432) );
  NOR2_X1 U494 ( .A1(n520), .A2(n433), .ZN(n434) );
  XNOR2_X1 U495 ( .A(n434), .B(KEYINPUT66), .ZN(n572) );
  XOR2_X1 U496 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n436) );
  XNOR2_X1 U497 ( .A(KEYINPUT23), .B(G204GAT), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n442) );
  XOR2_X1 U499 ( .A(G106GAT), .B(G218GAT), .Z(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U502 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U503 ( .A1(G228GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n445), .B(KEYINPUT22), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n471) );
  AND2_X1 U508 ( .A1(n572), .A2(n471), .ZN(n456) );
  INV_X1 U509 ( .A(KEYINPUT55), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U511 ( .A1(n472), .A2(n457), .ZN(n569) );
  NAND2_X1 U512 ( .A1(n569), .A2(n541), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  INV_X1 U514 ( .A(n573), .ZN(n560) );
  NAND2_X1 U515 ( .A1(n560), .A2(n411), .ZN(n490) );
  INV_X1 U516 ( .A(n472), .ZN(n533) );
  NAND2_X1 U517 ( .A1(n533), .A2(n524), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n460), .A2(n471), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT98), .ZN(n462) );
  XNOR2_X1 U520 ( .A(KEYINPUT25), .B(n462), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n524), .B(KEYINPUT27), .ZN(n469) );
  NOR2_X1 U522 ( .A1(n533), .A2(n471), .ZN(n464) );
  XNOR2_X1 U523 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n463) );
  XOR2_X1 U524 ( .A(n464), .B(n463), .Z(n571) );
  AND2_X1 U525 ( .A1(n469), .A2(n571), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n467), .A2(n520), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT99), .ZN(n474) );
  NAND2_X1 U529 ( .A1(n469), .A2(n520), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT96), .ZN(n545) );
  XOR2_X1 U531 ( .A(KEYINPUT28), .B(n471), .Z(n527) );
  NOR2_X1 U532 ( .A1(n545), .A2(n527), .ZN(n534) );
  NAND2_X1 U533 ( .A1(n534), .A2(n472), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n488) );
  NAND2_X1 U535 ( .A1(n582), .A2(n488), .ZN(n475) );
  XOR2_X1 U536 ( .A(KEYINPUT105), .B(n475), .Z(n476) );
  NOR2_X1 U537 ( .A1(n585), .A2(n476), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n477) );
  NOR2_X1 U539 ( .A1(n490), .A2(n519), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT38), .ZN(n506) );
  NAND2_X1 U541 ( .A1(n506), .A2(n533), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n482) );
  XOR2_X1 U543 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n487) );
  NAND2_X1 U544 ( .A1(n568), .A2(n485), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n489) );
  NAND2_X1 U546 ( .A1(n489), .A2(n488), .ZN(n509) );
  NOR2_X1 U547 ( .A1(n509), .A2(n490), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n491), .B(KEYINPUT100), .ZN(n501) );
  NAND2_X1 U549 ( .A1(n501), .A2(n520), .ZN(n495) );
  XOR2_X1 U550 ( .A(KEYINPUT102), .B(KEYINPUT34), .Z(n493) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(G1324GAT) );
  XOR2_X1 U554 ( .A(G8GAT), .B(KEYINPUT103), .Z(n497) );
  NAND2_X1 U555 ( .A1(n524), .A2(n501), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n499) );
  NAND2_X1 U558 ( .A1(n501), .A2(n533), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G15GAT), .B(n500), .ZN(G1326GAT) );
  NAND2_X1 U561 ( .A1(n501), .A2(n527), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  NAND2_X1 U564 ( .A1(n520), .A2(n506), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NAND2_X1 U566 ( .A1(n506), .A2(n524), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U568 ( .A1(n506), .A2(n527), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  NOR2_X1 U571 ( .A1(n551), .A2(n560), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(KEYINPUT109), .ZN(n518) );
  NOR2_X1 U573 ( .A1(n518), .A2(n509), .ZN(n514) );
  NAND2_X1 U574 ( .A1(n520), .A2(n514), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n524), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n533), .A2(n514), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U581 ( .A1(n514), .A2(n527), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(n517), .ZN(G1335GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n522) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n528), .A2(n520), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n528), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n533), .A2(n528), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n530) );
  NAND2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n532), .A2(n535), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n560), .A2(n542), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U602 ( .A1(n542), .A2(n565), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n542), .A2(n568), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U610 ( .A1(n532), .A2(n545), .ZN(n546) );
  NAND2_X1 U611 ( .A1(n546), .A2(n571), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n573), .A2(n556), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n551), .A2(n556), .ZN(n552) );
  XOR2_X1 U619 ( .A(n553), .B(n552), .Z(G1345GAT) );
  NOR2_X1 U620 ( .A1(n582), .A2(n556), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT118), .B(n558), .Z(n559) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n569), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n563) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT122), .B(n564), .Z(n567) );
  NAND2_X1 U632 ( .A1(n569), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n584) );
  NOR2_X1 U637 ( .A1(n573), .A2(n584), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT59), .B(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n411), .A2(n584), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

