//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n614, new_n615, new_n616, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919;
  XNOR2_X1  g000(.A(KEYINPUT67), .B(G197gat), .ZN(new_n202));
  INV_X1    g001(.A(G204gat), .ZN(new_n203));
  AND2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n202), .A2(new_n203), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n204), .A2(new_n205), .B1(KEYINPUT22), .B2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G211gat), .B(G218gat), .Z(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT29), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT68), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G155gat), .B(G162gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n211), .B1(new_n212), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n211), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n226), .B2(KEYINPUT29), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n225), .B1(new_n227), .B2(new_n221), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT71), .ZN(new_n229));
  OAI211_X1 g028(.A(G228gat), .B(G233gat), .C1(new_n225), .C2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n228), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G22gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G78gat), .B(G106gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT31), .ZN(new_n235));
  INV_X1    g034(.A(G50gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n231), .B(G22gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n237), .A2(KEYINPUT72), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n231), .A2(new_n232), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT72), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT73), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n233), .A2(new_n237), .B1(KEYINPUT72), .B2(new_n242), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n246), .A2(KEYINPUT73), .A3(new_n241), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT5), .ZN(new_n248));
  INV_X1    g047(.A(G120gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G113gat), .ZN(new_n250));
  INV_X1    g049(.A(G113gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G120gat), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT1), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G127gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G134gat), .ZN(new_n255));
  INV_X1    g054(.A(G127gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n253), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G134gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(KEYINPUT3), .B2(new_n221), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n224), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n259), .ZN(new_n263));
  OR3_X1    g062(.A1(new_n263), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n263), .B2(new_n221), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G225gat), .A2(G233gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n248), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n263), .B(new_n222), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(new_n268), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n224), .A2(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n274), .B2(new_n248), .ZN(new_n275));
  XNOR2_X1  g074(.A(G1gat), .B(G29gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT0), .ZN(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G85gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n279), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT6), .B1(new_n275), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n283), .B2(new_n275), .ZN(new_n285));
  INV_X1    g084(.A(new_n275), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(KEYINPUT6), .A3(new_n282), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT24), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(G183gat), .A3(G190gat), .ZN(new_n297));
  INV_X1    g096(.A(G183gat), .ZN(new_n298));
  INV_X1    g097(.A(G190gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT24), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n295), .B(new_n302), .C1(new_n294), .C2(new_n293), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n302), .B2(KEYINPUT64), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n303), .A2(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n299), .ZN(new_n310));
  XOR2_X1   g109(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n290), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(KEYINPUT26), .B2(new_n293), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n293), .A2(KEYINPUT26), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n314), .A2(new_n315), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(G226gat), .A3(G233gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n306), .A2(new_n307), .B1(new_n316), .B2(new_n312), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(KEYINPUT29), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n322), .A3(new_n211), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n211), .B1(new_n319), .B2(new_n322), .ZN(new_n325));
  XNOR2_X1  g124(.A(G8gat), .B(G36gat), .ZN(new_n326));
  INV_X1    g125(.A(G64gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G92gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  OR4_X1    g129(.A1(KEYINPUT30), .A2(new_n324), .A3(new_n325), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n325), .ZN(new_n332));
  INV_X1    g131(.A(new_n330), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n323), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n324), .B2(new_n325), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT30), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OAI22_X1  g137(.A1(new_n245), .A2(new_n247), .B1(new_n289), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n263), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n260), .ZN(new_n341));
  INV_X1    g140(.A(G227gat), .ZN(new_n342));
  INV_X1    g141(.A(G233gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT34), .ZN(new_n345));
  XNOR2_X1  g144(.A(G15gat), .B(G43gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(G71gat), .ZN(new_n347));
  INV_X1    g146(.A(G99gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  AOI211_X1 g148(.A(new_n342), .B(new_n343), .C1(new_n340), .C2(new_n341), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(KEYINPUT33), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n340), .A2(new_n341), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n342), .A2(new_n343), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n359), .B2(new_n349), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n345), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n345), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n351), .A2(new_n355), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(new_n359), .A3(new_n349), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT36), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT66), .B1(new_n356), .B2(new_n360), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n361), .A3(new_n365), .ZN(new_n370));
  OAI211_X1 g169(.A(KEYINPUT66), .B(new_n345), .C1(new_n356), .C2(new_n360), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n368), .B1(new_n372), .B2(new_n367), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n282), .B(KEYINPUT74), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n270), .B(new_n374), .C1(new_n274), .C2(new_n248), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n284), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT75), .B(KEYINPUT38), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n332), .A2(KEYINPUT37), .A3(new_n323), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT37), .B1(new_n332), .B2(new_n323), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n330), .B(new_n378), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n275), .A2(new_n283), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT6), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n376), .A2(new_n381), .A3(new_n383), .A4(new_n334), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n284), .A2(new_n375), .B1(new_n382), .B2(KEYINPUT6), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n387), .A2(KEYINPUT76), .A3(new_n334), .A4(new_n381), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n330), .B1(new_n379), .B2(new_n380), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n377), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n273), .A2(KEYINPUT39), .A3(new_n268), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n374), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n271), .A2(new_n268), .ZN(new_n394));
  OAI211_X1 g193(.A(KEYINPUT39), .B(new_n394), .C1(new_n273), .C2(new_n268), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(KEYINPUT40), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n331), .A2(new_n336), .A3(new_n375), .A4(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT40), .B1(new_n393), .B2(new_n395), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n244), .A2(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n391), .A2(new_n400), .A3(KEYINPUT77), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT77), .B1(new_n391), .B2(new_n400), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n339), .B(new_n373), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n370), .A2(new_n371), .B1(new_n246), .B2(new_n241), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n289), .A2(new_n338), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT35), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT35), .B1(new_n246), .B2(new_n241), .ZN(new_n408));
  INV_X1    g207(.A(new_n366), .ZN(new_n409));
  INV_X1    g208(.A(new_n387), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n408), .A2(new_n337), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n403), .A2(KEYINPUT78), .A3(new_n412), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G229gat), .A2(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n419));
  INV_X1    g218(.A(G29gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(KEYINPUT79), .A2(G29gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(G36gat), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(G29gat), .A2(G36gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n421), .A2(KEYINPUT80), .A3(G36gat), .A4(new_n422), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G43gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n236), .ZN(new_n432));
  NOR2_X1   g231(.A1(G43gat), .A2(G50gat), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT15), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n432), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT82), .B(G50gat), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(G43gat), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT81), .B(KEYINPUT15), .Z(new_n438));
  OAI21_X1  g237(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT17), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n445));
  INV_X1    g244(.A(G15gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n232), .ZN(new_n447));
  INV_X1    g246(.A(G1gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(G15gat), .A2(G22gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n447), .A2(new_n449), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n448), .A2(KEYINPUT16), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G8gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n450), .B2(KEYINPUT83), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n453), .B(new_n455), .Z(new_n456));
  INV_X1    g255(.A(KEYINPUT17), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n457), .A3(new_n442), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n444), .A2(new_n445), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n440), .A2(new_n457), .A3(new_n442), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n440), .B2(new_n442), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n453), .B(new_n455), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n443), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT84), .B1(new_n464), .B2(new_n462), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n418), .B(new_n459), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT18), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G113gat), .B(G141gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G197gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT11), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(new_n291), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT12), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n473), .B(G169gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT12), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n456), .A2(new_n443), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n462), .A2(new_n442), .A3(new_n440), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n418), .B(KEYINPUT13), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n445), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n444), .A2(new_n458), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n462), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n489), .A2(KEYINPUT18), .A3(new_n418), .A4(new_n459), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n468), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n479), .B1(new_n468), .B2(new_n469), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n468), .A2(new_n490), .A3(new_n486), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n417), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G99gat), .B(G106gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT7), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(G85gat), .A3(G92gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504));
  INV_X1    g303(.A(G85gat), .ZN(new_n505));
  AOI22_X1  g304(.A1(KEYINPUT8), .A2(new_n504), .B1(new_n505), .B2(new_n329), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n498), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n506), .A3(new_n498), .ZN(new_n509));
  NAND2_X1  g308(.A1(G71gat), .A2(G78gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT9), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n327), .A2(G57gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n327), .A2(G57gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n512), .B(KEYINPUT86), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G71gat), .B(G78gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G57gat), .B(G64gat), .Z(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT86), .A3(new_n516), .A4(new_n512), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n508), .A2(new_n509), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n522));
  INV_X1    g321(.A(new_n498), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n503), .A2(new_n524), .A3(new_n506), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n503), .B2(new_n506), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n522), .B(new_n523), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n503), .A2(new_n506), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT93), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n503), .A2(new_n506), .A3(new_n524), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n498), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n509), .A2(KEYINPUT94), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n518), .A2(new_n520), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT10), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538));
  INV_X1    g337(.A(new_n509), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(new_n507), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n508), .A2(KEYINPUT90), .A3(new_n509), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(KEYINPUT10), .A3(new_n534), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n518), .A2(new_n520), .ZN(new_n546));
  AOI211_X1 g345(.A(new_n536), .B(new_n546), .C1(new_n540), .C2(new_n541), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT95), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n537), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n535), .A2(new_n550), .ZN(new_n552));
  XNOR2_X1  g351(.A(G120gat), .B(G148gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(new_n292), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(new_n203), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n551), .B2(new_n552), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n534), .A2(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n462), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n456), .B1(KEYINPUT21), .B2(new_n534), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n534), .A2(KEYINPUT21), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G183gat), .B(G211gat), .Z(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n570), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G162gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT89), .B(G134gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n488), .A2(new_n542), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT91), .Z(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n464), .A2(new_n542), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n585), .B(new_n586), .C1(new_n488), .C2(new_n542), .ZN(new_n588));
  INV_X1    g387(.A(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI211_X1 g389(.A(KEYINPUT92), .B(new_n581), .C1(new_n587), .C2(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n587), .A2(KEYINPUT92), .A3(new_n590), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT92), .B1(new_n587), .B2(new_n590), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n594), .B2(new_n581), .ZN(new_n595));
  NOR4_X1   g394(.A1(new_n497), .A2(new_n560), .A3(new_n577), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n289), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g397(.A1(new_n417), .A2(new_n496), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n577), .A2(new_n595), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n559), .A3(new_n338), .A4(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT42), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n603), .A2(new_n605), .B1(G8gat), .B2(new_n601), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(new_n607), .ZN(G1325gat));
  AOI21_X1  g409(.A(G15gat), .B1(new_n596), .B2(new_n409), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n373), .A2(new_n446), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n596), .B2(new_n612), .ZN(G1326gat));
  OR2_X1    g412(.A1(new_n245), .A2(new_n247), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT43), .B(G22gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(G1327gat));
  INV_X1    g416(.A(new_n595), .ZN(new_n618));
  NOR4_X1   g417(.A1(new_n497), .A2(new_n560), .A3(new_n576), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n421), .A2(new_n422), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n289), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n621), .A2(KEYINPUT45), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(KEYINPUT45), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT44), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n415), .A2(new_n416), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n407), .A2(new_n627), .A3(new_n411), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT35), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n404), .B2(new_n405), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n631), .A2(new_n629), .A3(new_n337), .A4(new_n410), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n366), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT96), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n403), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n595), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n624), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n576), .A2(new_n560), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n626), .A2(new_n638), .A3(new_n496), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(new_n288), .ZN(new_n641));
  OAI22_X1  g440(.A1(new_n622), .A2(new_n623), .B1(new_n620), .B2(new_n641), .ZN(G1328gat));
  NAND3_X1  g441(.A1(new_n599), .A2(new_n595), .A3(new_n639), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n643), .A2(G36gat), .A3(new_n337), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT46), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(G36gat), .B1(new_n640), .B2(new_n337), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(G1329gat));
  NAND3_X1  g448(.A1(new_n619), .A2(new_n431), .A3(new_n409), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT47), .ZN(new_n651));
  OAI21_X1  g450(.A(G43gat), .B1(new_n640), .B2(new_n373), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n650), .B2(new_n652), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(G1330gat));
  OAI21_X1  g454(.A(new_n436), .B1(new_n640), .B2(new_n631), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n619), .A2(new_n614), .ZN(new_n657));
  OAI211_X1 g456(.A(KEYINPUT48), .B(new_n656), .C1(new_n657), .C2(new_n436), .ZN(new_n658));
  INV_X1    g457(.A(new_n614), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n643), .A2(new_n659), .A3(new_n436), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n640), .A2(new_n659), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n436), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n658), .B1(new_n662), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g462(.A(new_n496), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n600), .A2(new_n560), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT97), .Z(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n635), .B2(new_n403), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n289), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g468(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n337), .B(KEYINPUT98), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT99), .Z(new_n673));
  NOR2_X1   g472(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1333gat));
  INV_X1    g474(.A(new_n373), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n667), .A2(G71gat), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT100), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n667), .A2(new_n409), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(G71gat), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g480(.A1(new_n667), .A2(new_n614), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT101), .B(G78gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1335gat));
  NOR2_X1   g483(.A1(new_n576), .A2(new_n496), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n626), .A2(new_n638), .A3(new_n560), .A4(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G85gat), .B1(new_n686), .B2(new_n288), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n637), .A2(new_n496), .A3(new_n576), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT51), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n505), .A3(new_n560), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n690), .B2(new_n288), .ZN(G1336gat));
  NAND3_X1  g490(.A1(new_n671), .A2(new_n329), .A3(new_n560), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT102), .Z(new_n693));
  AND2_X1   g492(.A1(new_n688), .A2(KEYINPUT51), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n688), .A2(KEYINPUT51), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n671), .ZN(new_n697));
  OAI21_X1  g496(.A(G92gat), .B1(new_n686), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT52), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G92gat), .B1(new_n686), .B2(new_n337), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n700), .B(KEYINPUT103), .C1(new_n702), .C2(new_n699), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n699), .B1(new_n696), .B2(new_n701), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(G1337gat));
  OAI21_X1  g507(.A(G99gat), .B1(new_n686), .B2(new_n373), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n689), .A2(new_n348), .A3(new_n409), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(new_n559), .ZN(G1338gat));
  AND3_X1   g510(.A1(new_n626), .A2(new_n638), .A3(new_n685), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n712), .A2(KEYINPUT105), .A3(new_n560), .A4(new_n244), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n686), .B2(new_n631), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(G106gat), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n559), .A2(G106gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n689), .A2(new_n244), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT104), .B(KEYINPUT53), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n721));
  OAI21_X1  g520(.A(G106gat), .B1(new_n686), .B2(new_n659), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT53), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n716), .A2(new_n718), .A3(new_n725), .A4(new_n719), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n721), .A2(new_n724), .A3(new_n726), .ZN(G1339gat));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n600), .A2(new_n559), .A3(new_n664), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n418), .B1(new_n489), .B2(new_n459), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n474), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n494), .B2(new_n480), .ZN(new_n735));
  INV_X1    g534(.A(new_n550), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n535), .A2(new_n536), .B1(new_n547), .B2(KEYINPUT95), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n545), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT54), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n556), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n537), .A2(new_n736), .A3(new_n545), .A4(new_n548), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n551), .A2(KEYINPUT54), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT55), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n735), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(KEYINPUT54), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n738), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n549), .A2(new_n739), .A3(new_n550), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n555), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n557), .B1(new_n749), .B2(KEYINPUT55), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n595), .A2(new_n744), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n559), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n743), .B1(new_n492), .B2(new_n495), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n750), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n751), .B(KEYINPUT108), .C1(new_n754), .C2(new_n595), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n577), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n735), .A2(new_n559), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n493), .A2(new_n494), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n493), .A2(new_n494), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n557), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n758), .B2(new_n759), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n757), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n618), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT108), .B1(new_n767), .B2(new_n751), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n728), .B(new_n729), .C1(new_n756), .C2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n496), .A2(new_n750), .A3(new_n760), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n595), .B1(new_n772), .B2(new_n757), .ZN(new_n773));
  INV_X1    g572(.A(new_n751), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(new_n577), .A3(new_n755), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n728), .B1(new_n776), .B2(new_n729), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n779), .A2(new_n288), .A3(new_n671), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n781), .A2(new_n366), .A3(new_n614), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n664), .ZN(new_n784));
  INV_X1    g583(.A(new_n404), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n251), .A3(new_n496), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1340gat));
  OAI21_X1  g587(.A(G120gat), .B1(new_n783), .B2(new_n559), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n560), .A2(new_n249), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT110), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1341gat));
  NAND2_X1  g592(.A1(new_n786), .A2(new_n576), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT111), .Z(new_n795));
  NOR2_X1   g594(.A1(new_n577), .A2(new_n256), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n795), .A2(new_n256), .B1(new_n782), .B2(new_n796), .ZN(G1342gat));
  NOR4_X1   g596(.A1(new_n779), .A2(new_n288), .A3(new_n338), .A4(new_n618), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n258), .A3(new_n404), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT56), .Z(new_n800));
  OAI21_X1  g599(.A(G134gat), .B1(new_n783), .B2(new_n618), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1343gat));
  XOR2_X1   g601(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n803));
  NAND2_X1  g602(.A1(new_n758), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n496), .A2(new_n750), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(new_n757), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n751), .B1(new_n806), .B2(new_n595), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n577), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n809), .A2(new_n729), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT57), .B1(new_n811), .B2(new_n659), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n778), .A2(new_n813), .A3(new_n244), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n373), .A2(new_n289), .A3(new_n697), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT112), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n812), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n496), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G141gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n676), .A2(new_n631), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT116), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n780), .A2(new_n822), .ZN(new_n823));
  OR3_X1    g622(.A1(new_n823), .A2(G141gat), .A3(new_n664), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n818), .A2(new_n825), .A3(G141gat), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n820), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT58), .B1(new_n818), .B2(G141gat), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n829), .A2(KEYINPUT117), .A3(new_n824), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT117), .B1(new_n829), .B2(new_n824), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n827), .A2(new_n828), .B1(new_n830), .B2(new_n831), .ZN(G1344gat));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833));
  INV_X1    g632(.A(G148gat), .ZN(new_n834));
  AOI211_X1 g633(.A(KEYINPUT59), .B(new_n834), .C1(new_n817), .C2(new_n560), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n778), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n244), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n808), .A2(new_n729), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n614), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n813), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n729), .B1(new_n756), .B2(new_n768), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT109), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(KEYINPUT57), .A3(new_n244), .A4(new_n769), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n836), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n560), .A3(new_n816), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G148gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT59), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n835), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n823), .A2(G148gat), .A3(new_n559), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n833), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n855), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT120), .B1(new_n849), .B2(KEYINPUT59), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n851), .B(new_n859), .C1(new_n848), .C2(G148gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT121), .B(new_n857), .C1(new_n861), .C2(new_n835), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n856), .A2(new_n862), .ZN(G1345gat));
  OAI21_X1  g662(.A(new_n213), .B1(new_n823), .B2(new_n577), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n817), .A2(G155gat), .A3(new_n576), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(G1346gat));
  NAND3_X1  g665(.A1(new_n798), .A2(new_n214), .A3(new_n822), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n817), .A2(new_n595), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n214), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n778), .A2(new_n288), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(new_n785), .A3(new_n697), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n291), .A3(new_n496), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT122), .Z(new_n873));
  NAND2_X1  g672(.A1(new_n288), .A2(new_n338), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n366), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT123), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n778), .A2(new_n659), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n664), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n878), .ZN(G1348gat));
  NOR3_X1   g678(.A1(new_n877), .A2(new_n292), .A3(new_n559), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n871), .A2(new_n560), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n292), .ZN(G1349gat));
  NOR2_X1   g681(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n877), .A2(new_n577), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT124), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G183gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n309), .A3(new_n576), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n888), .B(new_n889), .Z(G1350gat));
  OAI21_X1  g689(.A(G190gat), .B1(new_n877), .B2(new_n618), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT61), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n871), .A2(new_n299), .A3(new_n595), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1351gat));
  NAND2_X1  g693(.A1(new_n821), .A2(new_n671), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT126), .ZN(new_n897));
  INV_X1    g696(.A(new_n870), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(KEYINPUT126), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(G197gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n496), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n676), .A2(new_n874), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n847), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(new_n496), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n902), .B1(new_n905), .B2(new_n901), .ZN(G1352gat));
  NAND3_X1  g705(.A1(new_n900), .A2(new_n203), .A3(new_n560), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(KEYINPUT62), .Z(new_n908));
  AND3_X1   g707(.A1(new_n847), .A2(new_n560), .A3(new_n903), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n203), .B2(new_n909), .ZN(G1353gat));
  AOI21_X1  g709(.A(new_n206), .B1(new_n904), .B2(new_n576), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(KEYINPUT63), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(KEYINPUT63), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n206), .A3(new_n576), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1354gat));
  AOI21_X1  g716(.A(G218gat), .B1(new_n900), .B2(new_n595), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n618), .A2(new_n207), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n904), .B2(new_n919), .ZN(G1355gat));
endmodule


