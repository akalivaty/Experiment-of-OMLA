//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n570, new_n571, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n459), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(new_n469), .ZN(G160));
  OAI21_X1  g045(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G112), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(G124), .A3(G2105), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT68), .ZN(new_n476));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI211_X1 g054(.A(new_n473), .B(new_n476), .C1(G136), .C2(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n459), .B2(G114), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G102), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n459), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n482), .A2(new_n484), .A3(G2104), .A4(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n474), .A2(new_n492), .A3(G138), .A4(new_n459), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n504), .A2(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  INV_X1    g088(.A(new_n509), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(new_n515), .B1(new_n497), .B2(new_n498), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n496), .B1(new_n514), .B2(new_n515), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n502), .B1(new_n513), .B2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n499), .A2(G63), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT71), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n516), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n519), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n507), .A2(new_n506), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n501), .B1(new_n534), .B2(KEYINPUT72), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n535), .B1(KEYINPUT72), .B2(new_n534), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n516), .A2(G90), .B1(new_n519), .B2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AOI22_X1  g114(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n501), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT73), .B(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n504), .A2(new_n542), .B1(new_n510), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  OR3_X1    g121(.A1(new_n541), .A2(new_n544), .A3(KEYINPUT74), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(new_n501), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n532), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n560), .A2(KEYINPUT76), .A3(G651), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n504), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n519), .A2(new_n565), .A3(G53), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n564), .A2(new_n566), .B1(G91), .B2(new_n516), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  NOR2_X1   g144(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n518), .B1(new_n517), .B2(new_n520), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n570), .A2(new_n571), .B1(new_n501), .B2(new_n500), .ZN(G303));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n497), .A2(new_n573), .A3(new_n498), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n519), .A2(G49), .B1(new_n574), .B2(G651), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT77), .B1(new_n516), .B2(G87), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT77), .A4(G87), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n575), .B1(new_n576), .B2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n497), .B2(new_n498), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n516), .A2(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n519), .A2(G48), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n516), .A2(G85), .B1(new_n519), .B2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n501), .B2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n519), .A2(G54), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n499), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n501), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n516), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G284));
  XOR2_X1   g176(.A(G284), .B(KEYINPUT80), .Z(G321));
  MUX2_X1   g177(.A(G299), .B(G286), .S(G868), .Z(G297));
  XOR2_X1   g178(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n600), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n600), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n474), .A2(new_n466), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n479), .A2(G135), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n459), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n474), .A2(G2105), .ZN(new_n619));
  OAI221_X1 g194(.A(new_n615), .B1(new_n616), .B2(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT82), .B(G2096), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n614), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT84), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2427), .B(G2430), .Z(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n630), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(G14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT85), .Z(G401));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n645), .B2(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT86), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n643), .A2(new_n644), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n648), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n656), .A2(new_n660), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT87), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(KEYINPUT87), .ZN(new_n666));
  AOI211_X1 g241(.A(new_n661), .B(new_n663), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1991), .B(G1996), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1981), .B(G1986), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n669), .B(new_n673), .ZN(G229));
  MUX2_X1   g249(.A(G6), .B(G305), .S(G16), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT32), .ZN(new_n676));
  INV_X1    g251(.A(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G22), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G166), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G1971), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n679), .A2(G23), .ZN(new_n687));
  OAI211_X1 g262(.A(G49), .B(G543), .C1(new_n508), .C2(new_n509), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n507), .A2(new_n506), .A3(G74), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n501), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT77), .ZN(new_n691));
  INV_X1    g266(.A(G87), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n510), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n690), .B1(new_n693), .B2(new_n577), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n687), .B1(new_n694), .B2(new_n679), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n678), .A2(new_n685), .A3(new_n686), .A4(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n479), .A2(G131), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n459), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G119), .ZN(new_n704));
  OAI221_X1 g279(.A(new_n701), .B1(new_n702), .B2(new_n703), .C1(new_n704), .C2(new_n619), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n705), .S(G29), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G24), .B(G290), .S(G16), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT89), .B(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT91), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n709), .B(new_n712), .C1(new_n713), .C2(KEYINPUT36), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n699), .A2(new_n700), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(KEYINPUT36), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n679), .A2(G19), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n548), .B2(new_n679), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1341), .ZN(new_n721));
  NOR2_X1   g296(.A1(G4), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n600), .B2(G16), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n721), .B1(G1348), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G35), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT95), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT29), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n724), .B1(G2090), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n723), .A2(G1348), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n729), .B2(G2090), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n725), .A2(G32), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n474), .A2(G129), .A3(G2105), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  AND3_X1   g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n733), .B1(new_n738), .B2(new_n725), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n679), .A2(G21), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G168), .B2(new_n679), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n741), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n725), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n725), .ZN(new_n748));
  INV_X1    g323(.A(G2078), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT30), .B(G28), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n751), .A2(new_n725), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n620), .B2(new_n725), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n725), .B1(new_n756), .B2(G34), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n756), .B2(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G160), .B2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n755), .B1(G2084), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n750), .B(new_n760), .C1(G2084), .C2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n479), .A2(G140), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n459), .A2(G116), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n764));
  INV_X1    g339(.A(G128), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n762), .B1(new_n763), .B2(new_n764), .C1(new_n765), .C2(new_n619), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n725), .A2(G26), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT28), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n744), .A2(G1966), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n746), .A2(new_n761), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n474), .A2(G127), .ZN(new_n774));
  AND2_X1   g349(.A1(G115), .A2(G2104), .ZN(new_n775));
  OAI21_X1  g350(.A(G2105), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n479), .A2(G139), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT93), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G29), .ZN(new_n782));
  NOR2_X1   g357(.A1(G29), .A2(G33), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT92), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G2072), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(G5), .A2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT94), .Z(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G301), .B2(new_n679), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n787), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n788), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n785), .B2(new_n786), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n732), .A2(new_n773), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n679), .A2(G20), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G299), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT98), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT97), .B(G1956), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n730), .A2(new_n795), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n717), .A2(new_n718), .A3(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  AOI22_X1  g380(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n501), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT100), .B(G55), .Z(new_n808));
  INV_X1    g383(.A(G93), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n504), .A2(new_n808), .B1(new_n510), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  NAND3_X1  g389(.A1(new_n546), .A2(new_n547), .A3(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n545), .A2(new_n811), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT101), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n599), .A2(new_n605), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT102), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(G860), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n828), .A2(KEYINPUT103), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT103), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n814), .B1(new_n830), .B2(new_n831), .ZN(G145));
  INV_X1    g407(.A(KEYINPUT105), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n489), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n491), .A2(new_n493), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n487), .A2(KEYINPUT105), .A3(new_n488), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n766), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(new_n738), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n738), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n781), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT106), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT107), .ZN(new_n844));
  INV_X1    g419(.A(G130), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n459), .A2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n619), .A2(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n479), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n612), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n705), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n850), .A2(new_n705), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n844), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n855), .A2(KEYINPUT107), .A3(new_n851), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n841), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n780), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n841), .A2(new_n861), .A3(new_n781), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n843), .A2(new_n858), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G162), .B(new_n620), .ZN(new_n864));
  XNOR2_X1  g439(.A(G160), .B(KEYINPUT104), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n843), .A2(new_n860), .A3(new_n862), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n855), .A3(new_n851), .ZN(new_n869));
  AOI21_X1  g444(.A(G37), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n863), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n857), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT108), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT108), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n868), .A2(new_n874), .A3(new_n857), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n871), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n870), .B1(new_n876), .B2(new_n866), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g453(.A(new_n821), .B(new_n607), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n599), .A2(G299), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n596), .A2(new_n562), .A3(new_n567), .A4(new_n598), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n881), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n879), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n889));
  XNOR2_X1  g464(.A(G166), .B(new_n694), .ZN(new_n890));
  XNOR2_X1  g465(.A(G290), .B(G305), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n884), .A2(new_n887), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n889), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n893), .B1(new_n889), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(G868), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(G868), .B2(new_n811), .ZN(G295));
  OAI21_X1  g474(.A(new_n898), .B1(G868), .B2(new_n811), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n901));
  NAND2_X1  g476(.A1(G171), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n536), .B2(new_n537), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(G168), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(G301), .A2(KEYINPUT109), .ZN(new_n906));
  OAI21_X1  g481(.A(G286), .B1(new_n906), .B2(new_n903), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n818), .A2(new_n820), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(new_n883), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n907), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT110), .B1(new_n821), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n905), .A2(new_n907), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n818), .A4(new_n820), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n886), .A2(new_n885), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n821), .A2(new_n910), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n908), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n892), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n915), .A2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n893), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n915), .A2(KEYINPUT111), .A3(new_n918), .A4(new_n892), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n908), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n914), .A2(new_n911), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n930), .A2(new_n916), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n917), .A2(new_n883), .A3(new_n908), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n893), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n919), .B2(new_n920), .ZN(new_n934));
  AND4_X1   g509(.A1(KEYINPUT43), .A2(new_n933), .A3(new_n934), .A4(new_n925), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n928), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n933), .A2(new_n934), .A3(new_n927), .A4(new_n925), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(G397));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n492), .B1(new_n479), .B2(G138), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n836), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT105), .B1(new_n487), .B2(new_n488), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n464), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(G40), .A3(new_n467), .A4(new_n468), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n766), .B(G2067), .Z(new_n954));
  XNOR2_X1  g529(.A(new_n738), .B(G1996), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n705), .B(new_n707), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(G1986), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT117), .ZN(new_n961));
  NAND3_X1  g536(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n963));
  INV_X1    g538(.A(G8), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(G166), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n837), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n967));
  INV_X1    g542(.A(G40), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n464), .A2(new_n469), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n487), .A2(new_n488), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n835), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n682), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n948), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G2090), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n952), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n973), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n964), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n973), .A2(new_n980), .A3(KEYINPUT115), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n966), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(G1976), .B(new_n575), .C1(new_n576), .C2(new_n578), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT113), .B1(new_n694), .B2(G1976), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n837), .A2(new_n943), .A3(new_n969), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G8), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT114), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n986), .A2(new_n987), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n694), .A2(KEYINPUT113), .A3(G1976), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n997), .A3(G8), .A4(new_n991), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(KEYINPUT52), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n835), .A2(new_n970), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n943), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n952), .B1(new_n1001), .B2(new_n949), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT45), .B(new_n943), .C1(new_n946), .C2(new_n947), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1971), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n943), .B(new_n974), .C1(new_n946), .C2(new_n947), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1006));
  AND4_X1   g581(.A1(new_n977), .A2(new_n1005), .A3(new_n969), .A4(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(G8), .B(new_n966), .C1(new_n1004), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n996), .A2(G8), .A3(new_n991), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G48), .ZN(new_n1012));
  INV_X1    g587(.A(G86), .ZN(new_n1013));
  OAI22_X1  g588(.A1(new_n504), .A2(new_n1012), .B1(new_n510), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n580), .B(KEYINPUT78), .ZN(new_n1015));
  OAI21_X1  g590(.A(G61), .B1(new_n507), .B2(new_n506), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n501), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(G1981), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n585), .A2(new_n586), .A3(new_n677), .A4(new_n587), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(KEYINPUT49), .A3(new_n1019), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1022), .A2(G8), .A3(new_n991), .A4(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1011), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n999), .A2(new_n1008), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n985), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n969), .B1(new_n1001), .B2(new_n949), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n837), .B2(new_n943), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1028), .B(new_n742), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1005), .A2(new_n1006), .A3(new_n1032), .A4(new_n969), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n952), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n950), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1028), .B1(new_n1036), .B2(new_n742), .ZN(new_n1037));
  OAI211_X1 g612(.A(G8), .B(G168), .C1(new_n1034), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n961), .B1(new_n1027), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n969), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n974), .B1(new_n837), .B2(new_n943), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1041), .A2(new_n1042), .A3(G2090), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n982), .B1(new_n1043), .B2(new_n1004), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(new_n984), .A3(G8), .ZN(new_n1045));
  INV_X1    g620(.A(new_n966), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n999), .A2(new_n1008), .A3(new_n1025), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n1039), .A4(new_n961), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT118), .B1(new_n1040), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(new_n1048), .A3(new_n1039), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT117), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1050), .A4(new_n1049), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1050), .B1(new_n1057), .B2(new_n1046), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1048), .A2(new_n1039), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1052), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1348), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n837), .A2(new_n943), .A3(new_n974), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n969), .B1(new_n971), .B2(new_n978), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n991), .A2(G2067), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(new_n599), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n562), .A2(new_n567), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n562), .B2(new_n567), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1002), .A2(new_n1003), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1072), .B(new_n1074), .C1(new_n1075), .C2(G1956), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1067), .A2(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1002), .A2(new_n1003), .A3(new_n1073), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1956), .B1(new_n976), .B2(new_n979), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1066), .A2(KEYINPUT60), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1064), .A2(KEYINPUT60), .A3(new_n1065), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n600), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n599), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1066), .A2(KEYINPUT120), .A3(KEYINPUT60), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1083), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT58), .B(G1341), .Z(new_n1092));
  NAND2_X1  g667(.A1(new_n991), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n949), .B1(G164), .B2(G1384), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1003), .A2(new_n1094), .A3(new_n969), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1095), .B2(G1996), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n548), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT59), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1099), .A3(new_n548), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1081), .A2(KEYINPUT61), .A3(new_n1076), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1081), .A2(new_n1103), .A3(new_n1076), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1078), .B(KEYINPUT119), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1101), .B(new_n1102), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1082), .B1(new_n1091), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1003), .A2(new_n1094), .A3(new_n749), .A4(new_n969), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n788), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n952), .A2(new_n1113), .A3(G2078), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n950), .B(new_n1117), .C1(new_n949), .C2(new_n1001), .ZN(new_n1118));
  AOI21_X1  g693(.A(G301), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n950), .A2(new_n1003), .A3(new_n1117), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1114), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1111), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1111), .B1(new_n1121), .B2(G171), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1114), .A2(new_n1118), .A3(new_n1115), .A4(G301), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT124), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1121), .A2(G171), .ZN(new_n1127));
  AND4_X1   g702(.A1(KEYINPUT124), .A2(new_n1127), .A3(KEYINPUT54), .A4(new_n1125), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1027), .B(new_n1123), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(new_n964), .A3(G168), .ZN(new_n1131));
  OAI21_X1  g706(.A(G8), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT123), .B(G8), .C1(new_n1034), .C2(new_n1037), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G168), .A2(new_n964), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(KEYINPUT51), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1136), .B(KEYINPUT122), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT51), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1131), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1129), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1144), .B(new_n1082), .C1(new_n1091), .C2(new_n1108), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1110), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1024), .A2(new_n1009), .A3(new_n694), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n992), .B1(new_n1147), .B2(new_n1019), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n999), .A2(new_n1025), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1008), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1060), .A2(new_n1146), .A3(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1027), .A2(new_n1119), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1142), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1137), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1157), .A2(new_n1135), .B1(new_n1140), .B2(KEYINPUT51), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1158), .A2(KEYINPUT62), .A3(new_n1131), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT125), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1142), .A2(new_n1154), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT62), .B1(new_n1158), .B2(new_n1131), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1153), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n960), .B1(new_n1152), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n953), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1167), .A2(G1996), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT46), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n954), .A2(new_n738), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n953), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT47), .ZN(new_n1175));
  OR3_X1    g750(.A1(new_n1167), .A2(G1986), .A3(G290), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT48), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n958), .A2(new_n953), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n705), .A2(new_n708), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n956), .B2(new_n1167), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n766), .A2(G2067), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT126), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1183), .A2(KEYINPUT126), .A3(new_n1184), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n953), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1181), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1175), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1166), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g765(.A(G319), .ZN(new_n1192));
  INV_X1    g766(.A(new_n640), .ZN(new_n1193));
  NOR4_X1   g767(.A1(G229), .A2(new_n1192), .A3(new_n1193), .A4(G227), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n939), .A2(new_n877), .A3(new_n1194), .ZN(G225));
  INV_X1    g769(.A(G225), .ZN(G308));
endmodule


