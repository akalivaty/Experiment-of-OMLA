//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n522, new_n523, new_n524, new_n525, new_n526, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n535, new_n537,
    new_n538, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n460), .A2(G137), .A3(new_n459), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n459), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n463), .A2(new_n467), .ZN(G160));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G136), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  MUX2_X1   g049(.A(G100), .B(G112), .S(G2105), .Z(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  NAND2_X1  g053(.A1(G114), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G102), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n459), .C1(new_n483), .C2(new_n484), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n460), .A2(new_n489), .A3(G138), .A4(new_n459), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(G164));
  INV_X1    g066(.A(G651), .ZN(new_n492));
  OR2_X1    g067(.A1(KEYINPUT5), .A2(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT5), .A2(G543), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G62), .ZN(new_n496));
  NAND2_X1  g071(.A1(G75), .A2(G543), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(new_n499), .A3(G88), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(G50), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n498), .A2(new_n502), .ZN(G166));
  NAND3_X1  g078(.A1(new_n495), .A2(G63), .A3(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT7), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n499), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G51), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT67), .B(G89), .Z(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n508), .A2(new_n511), .A3(new_n519), .ZN(G286));
  INV_X1    g095(.A(G286), .ZN(G168));
  AOI22_X1  g096(.A1(new_n495), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n492), .ZN(new_n523));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  INV_X1    g099(.A(G90), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n509), .A2(new_n524), .B1(new_n516), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G171));
  AOI22_X1  g102(.A1(new_n495), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n492), .ZN(new_n529));
  INV_X1    g104(.A(G43), .ZN(new_n530));
  INV_X1    g105(.A(G81), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n509), .A2(new_n530), .B1(new_n516), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G860), .ZN(G153));
  AND3_X1   g109(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G36), .ZN(G176));
  NAND2_X1  g111(.A1(G1), .A2(G3), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT8), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(G188));
  INV_X1    g114(.A(G65), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n493), .A2(new_n541), .A3(new_n494), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT70), .B1(new_n513), .B2(new_n512), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(G78), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(G651), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n516), .A2(KEYINPUT69), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n495), .A2(new_n499), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(G91), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n499), .A2(G53), .A3(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n499), .A2(new_n555), .A3(G53), .A4(G543), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n554), .B1(new_n553), .B2(new_n556), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n547), .B(new_n551), .C1(new_n557), .C2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  NAND2_X1  g135(.A1(new_n496), .A2(new_n497), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n562), .A2(new_n563), .A3(new_n500), .A4(new_n501), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT71), .B1(new_n498), .B2(new_n502), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(G303));
  NOR2_X1   g141(.A1(new_n513), .A2(new_n512), .ZN(new_n567));
  INV_X1    g142(.A(G74), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n492), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n510), .B2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n548), .A2(G87), .A3(new_n550), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(G288));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n493), .B2(new_n494), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(KEYINPUT72), .ZN(new_n575));
  OAI211_X1 g150(.A(KEYINPUT72), .B(G61), .C1(new_n513), .C2(new_n512), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n548), .A2(G86), .A3(new_n550), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n510), .A2(G48), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n517), .A2(G85), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n510), .A2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n495), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n492), .C2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n548), .A2(G92), .A3(new_n550), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n590), .A2(new_n591), .B1(G54), .B2(new_n510), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n542), .A2(new_n543), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n492), .B1(new_n594), .B2(KEYINPUT73), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(KEYINPUT73), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G321));
  MUX2_X1   g176(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g177(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n599), .B1(new_n604), .B2(G860), .ZN(G148));
  INV_X1    g180(.A(new_n533), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n599), .A2(new_n604), .ZN(new_n607));
  MUX2_X1   g182(.A(new_n606), .B(new_n607), .S(G868), .Z(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n471), .A2(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(KEYINPUT13), .B1(KEYINPUT76), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT13), .B2(new_n613), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n616), .A2(KEYINPUT76), .A3(new_n614), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(KEYINPUT76), .B2(new_n614), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n471), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n473), .A2(G123), .ZN(new_n620));
  MUX2_X1   g195(.A(G99), .B(G111), .S(G2105), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G2104), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT77), .B(G2096), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n617), .A2(new_n618), .A3(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT81), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT78), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(KEYINPUT14), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT80), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT16), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n635), .A2(new_n639), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n641), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n641), .B2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n631), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n650), .A2(new_n646), .A3(new_n630), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n651), .A3(G14), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n654), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(new_n656), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n660), .B2(new_n661), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n654), .A2(new_n656), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n655), .B1(new_n665), .B2(KEYINPUT17), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n659), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n667), .A2(G2096), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(G2096), .ZN(new_n669));
  OR3_X1    g244(.A1(new_n668), .A2(new_n669), .A3(new_n614), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n614), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT83), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(G229));
  NOR2_X1   g266(.A1(G6), .A2(G16), .ZN(new_n692));
  INV_X1    g267(.A(G305), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(G16), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT32), .B(G1981), .Z(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G23), .ZN(new_n698));
  INV_X1    g273(.A(G288), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT84), .B(G16), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G22), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1971), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n696), .A2(new_n702), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n704), .A2(G24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G290), .B2(new_n703), .ZN(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n715));
  OAI22_X1  g290(.A1(new_n713), .A2(new_n714), .B1(KEYINPUT85), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G25), .A2(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n471), .A2(G131), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n473), .A2(G119), .ZN(new_n719));
  MUX2_X1   g294(.A(G95), .B(G107), .S(G2105), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G2104), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n717), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  AOI211_X1 g301(.A(new_n716), .B(new_n726), .C1(new_n714), .C2(new_n713), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n710), .A2(new_n711), .A3(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n715), .A2(KEYINPUT85), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G21), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G168), .B2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT88), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT89), .Z(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G33), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n465), .A2(G103), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT25), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n471), .A2(G139), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n459), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(new_n737), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2072), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n471), .A2(G140), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n460), .A2(G128), .A3(G2105), .ZN(new_n749));
  NAND2_X1  g324(.A1(G116), .A2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G104), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G2104), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n748), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n737), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n704), .A2(G19), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n533), .B2(new_n704), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1341), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n747), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT86), .B(KEYINPUT24), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G34), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(new_n737), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G160), .B2(new_n737), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT91), .ZN(new_n771));
  NAND2_X1  g346(.A1(G162), .A2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G29), .B2(G35), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(G2090), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G27), .A2(G29), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G164), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2078), .ZN(new_n780));
  INV_X1    g355(.A(G2090), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n780), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n623), .A2(new_n737), .ZN(new_n783));
  OR2_X1    g358(.A1(KEYINPUT30), .A2(G28), .ZN(new_n784));
  NAND2_X1  g359(.A1(KEYINPUT30), .A2(G28), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT31), .B(G11), .Z(new_n787));
  NOR3_X1   g362(.A1(new_n783), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n697), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G171), .B2(new_n697), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n788), .B1(new_n790), .B2(G1961), .C1(new_n768), .C2(new_n769), .ZN(new_n791));
  NOR2_X1   g366(.A1(G29), .A2(G32), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT26), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n460), .A2(G141), .A3(new_n459), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n460), .A2(G129), .A3(G2105), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n465), .A2(G105), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n792), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT87), .Z(new_n802));
  XOR2_X1   g377(.A(KEYINPUT27), .B(G1996), .Z(new_n803));
  AOI21_X1  g378(.A(new_n791), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n763), .A2(new_n777), .A3(new_n782), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n703), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT23), .ZN(new_n807));
  INV_X1    g382(.A(G299), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n697), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1956), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n790), .A2(G1961), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT90), .ZN(new_n812));
  OAI221_X1 g387(.A(new_n812), .B1(new_n802), .B2(new_n803), .C1(new_n733), .C2(new_n734), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n736), .A2(new_n805), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n728), .A2(new_n729), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n697), .A2(G4), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n599), .B2(new_n697), .ZN(new_n817));
  INV_X1    g392(.A(G1348), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n730), .A2(new_n814), .A3(new_n815), .A4(new_n819), .ZN(G150));
  INV_X1    g395(.A(G150), .ZN(G311));
  AOI22_X1  g396(.A1(new_n495), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n492), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n509), .A2(new_n824), .B1(new_n516), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n533), .A2(new_n827), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n529), .A2(new_n532), .B1(new_n823), .B2(new_n826), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT38), .Z(new_n831));
  INV_X1    g406(.A(new_n599), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n604), .ZN(new_n833));
  INV_X1    g408(.A(new_n831), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(G559), .A3(new_n599), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(G860), .B1(new_n836), .B2(KEYINPUT39), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n833), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT93), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n827), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT94), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT95), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n843), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n853));
  INV_X1    g428(.A(new_n745), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n754), .B(KEYINPUT98), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n488), .A2(new_n490), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n486), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT97), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n800), .A2(new_n856), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n856), .A3(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n799), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n855), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n855), .B1(new_n862), .B2(new_n860), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT99), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n862), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n754), .B(KEYINPUT98), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n870), .A3(new_n863), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n854), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n864), .B2(new_n865), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(KEYINPUT100), .A3(new_n863), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n874), .B1(new_n878), .B2(new_n854), .ZN(new_n879));
  AOI211_X1 g454(.A(KEYINPUT101), .B(new_n745), .C1(new_n876), .C2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI22_X1  g456(.A1(G130), .A2(new_n473), .B1(new_n471), .B2(G142), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n883), .A2(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(KEYINPUT102), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n884), .B(new_n885), .C1(G118), .C2(new_n459), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n722), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n612), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  XOR2_X1   g467(.A(G160), .B(KEYINPUT96), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n477), .B(new_n623), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n873), .B(new_n889), .C1(new_n879), .C2(new_n880), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n891), .A2(new_n892), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT103), .B1(new_n881), .B2(new_n890), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n895), .B1(new_n900), .B2(new_n896), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n853), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n895), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n878), .A2(new_n854), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT101), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n878), .A2(new_n874), .A3(new_n854), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n872), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n892), .B1(new_n907), .B2(new_n889), .ZN(new_n908));
  INV_X1    g483(.A(new_n896), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n898), .A4(new_n897), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n902), .A2(new_n911), .ZN(G395));
  NOR2_X1   g487(.A1(new_n844), .A2(G868), .ZN(new_n913));
  INV_X1    g488(.A(new_n830), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n607), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n808), .A2(new_n592), .A3(new_n596), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n808), .B1(new_n596), .B2(new_n592), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n597), .A2(G299), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n917), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n918), .A2(new_n919), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n926), .B2(new_n915), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n693), .A2(G166), .ZN(new_n928));
  OAI21_X1  g503(.A(G305), .B1(new_n498), .B2(new_n502), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(G290), .A2(G288), .ZN(new_n931));
  NAND2_X1  g506(.A1(G290), .A2(G288), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n928), .A2(new_n931), .A3(new_n932), .A4(new_n929), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT42), .B1(new_n934), .B2(new_n936), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n927), .A2(new_n943), .ZN(new_n944));
  OAI221_X1 g519(.A(new_n924), .B1(new_n926), .B2(new_n915), .C1(new_n942), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n913), .B1(new_n946), .B2(G868), .ZN(G295));
  AOI21_X1  g522(.A(new_n913), .B1(new_n946), .B2(G868), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  OAI21_X1  g524(.A(G286), .B1(new_n523), .B2(new_n526), .ZN(new_n950));
  NAND4_X1  g525(.A1(G171), .A2(new_n508), .A3(new_n511), .A4(new_n519), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n830), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(KEYINPUT106), .A3(new_n830), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n914), .A2(new_n950), .A3(new_n951), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n920), .A2(new_n958), .A3(new_n922), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n925), .A2(new_n953), .A3(new_n957), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n939), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n898), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n926), .A2(new_n958), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n953), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n920), .A2(new_n922), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n939), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n949), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n959), .A2(new_n960), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n940), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(new_n961), .A3(KEYINPUT43), .A4(new_n898), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n969), .A2(new_n961), .A3(new_n949), .A4(new_n898), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n973), .A2(KEYINPUT44), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n962), .B2(new_n966), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT107), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND4_X1   g551(.A1(KEYINPUT107), .A2(new_n975), .A3(KEYINPUT44), .A4(new_n973), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n861), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n463), .A2(new_n467), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n754), .B(G2067), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT108), .ZN(new_n986));
  INV_X1    g561(.A(G1996), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n799), .B(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n723), .A2(new_n725), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n723), .A2(new_n725), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(G290), .B(G1986), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n984), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n576), .A2(new_n577), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT72), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n567), .B2(new_n573), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n492), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G48), .ZN(new_n1001));
  INV_X1    g576(.A(G86), .ZN(new_n1002));
  OAI22_X1  g577(.A1(new_n509), .A2(new_n1001), .B1(new_n516), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G1981), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n579), .A2(new_n1005), .A3(new_n580), .A4(new_n581), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT49), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n982), .A2(new_n979), .A3(new_n861), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(new_n1006), .A3(KEYINPUT49), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n996), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1008), .A2(G8), .ZN(new_n1016));
  AND4_X1   g591(.A1(new_n996), .A2(new_n1015), .A3(new_n1016), .A4(new_n1011), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n699), .B2(G1976), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G288), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n1009), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1016), .A2(new_n1022), .A3(new_n1024), .A4(new_n1020), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n995), .B1(new_n1018), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(KEYINPUT110), .B2(KEYINPUT55), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n564), .A2(new_n565), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n564), .A2(new_n565), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(G164), .B2(G1384), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n982), .A3(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT109), .B(G1971), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n861), .A2(KEYINPUT50), .A3(new_n979), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(G164), .B2(G1384), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n982), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1044), .B1(new_n1049), .B2(G2090), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1038), .B1(new_n1050), .B2(G8), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n861), .A2(new_n1046), .A3(new_n979), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n982), .A3(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1055), .A2(G2090), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1052), .B1(new_n1056), .B2(new_n1044), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1051), .B1(new_n1057), .B2(new_n1038), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1015), .A2(new_n1016), .A3(new_n1011), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT112), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1010), .A2(new_n996), .A3(new_n1011), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1062), .A2(KEYINPUT115), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1029), .A2(new_n1058), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G160), .A2(G40), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT53), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n980), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n482), .A2(new_n485), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1040), .B(G1384), .C1(new_n856), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1039), .A2(new_n1041), .A3(new_n1066), .A4(new_n982), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1068), .A2(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n861), .A2(new_n1046), .A3(new_n979), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1384), .B1(new_n856), .B2(new_n1069), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n982), .B1(new_n1076), .B2(new_n1046), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1961), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1053), .A2(new_n1054), .A3(new_n1080), .A4(new_n982), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1074), .A2(G301), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT54), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1082), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n979), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1065), .B1(new_n1086), .B2(new_n1040), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(KEYINPUT53), .A3(new_n1066), .A4(new_n1039), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(G171), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT125), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(G171), .C1(new_n1085), .C2(new_n1090), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1084), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1068), .A2(new_n1039), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1097), .A2(G301), .A3(new_n1082), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G286), .A2(G8), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  NAND3_X1  g679(.A1(G286), .A2(KEYINPUT122), .A3(G8), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n980), .A2(new_n1065), .A3(new_n1070), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1107), .A2(G1966), .B1(new_n1055), .B2(G2084), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1108), .B2(G8), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1966), .B1(new_n1087), .B2(new_n1071), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1055), .A2(G2084), .ZN(new_n1111));
  OAI21_X1  g686(.A(G8), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT124), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1103), .A2(new_n1115), .A3(new_n1105), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT123), .B(KEYINPUT51), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1109), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1100), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1095), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT117), .B(G1956), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1049), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n513), .A2(new_n512), .A3(KEYINPUT70), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n541), .B1(new_n493), .B2(new_n494), .ZN(new_n1129));
  OAI21_X1  g704(.A(G65), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n492), .B1(new_n1130), .B2(new_n545), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n548), .A2(G91), .A3(new_n550), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1127), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n547), .A2(KEYINPUT118), .A3(new_n551), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT57), .B1(new_n553), .B2(new_n556), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1135), .A2(new_n1136), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1039), .A2(new_n1041), .A3(new_n982), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1126), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1078), .A2(new_n818), .A3(new_n1081), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1008), .A2(G2067), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n597), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1137), .B1(new_n1126), .B2(new_n1139), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1140), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT120), .B(new_n1140), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1065), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1125), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1139), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n547), .A2(KEYINPUT118), .A3(new_n551), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT118), .B1(new_n547), .B2(new_n551), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1136), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1149), .B1(new_n1144), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT58), .B(G1341), .Z(new_n1160));
  NAND2_X1  g735(.A1(new_n1008), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1042), .B2(G1996), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n533), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1165), .A3(new_n533), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1168));
  INV_X1    g743(.A(new_n597), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(KEYINPUT60), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n597), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1171), .A2(new_n1141), .A3(new_n1142), .A4(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1159), .A2(new_n1167), .A3(new_n1170), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n1152), .A2(new_n1157), .A3(KEYINPUT121), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1149), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1147), .B(new_n1148), .C1(new_n1175), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1124), .A2(new_n1180), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1122), .A2(KEYINPUT62), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1122), .A2(KEYINPUT62), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n1099), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1064), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1112), .A2(G286), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1029), .A2(new_n1058), .A3(new_n1063), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1062), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1190), .A2(G286), .A3(new_n1112), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1057), .B1(KEYINPUT116), .B2(new_n1038), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1056), .A2(new_n1044), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(G8), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1038), .A2(KEYINPUT116), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1188), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1191), .A2(new_n1192), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1189), .A2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1190), .A2(new_n1194), .A3(new_n1037), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n699), .A2(new_n1023), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT113), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1062), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(KEYINPUT114), .B1(new_n1202), .B2(new_n1006), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1203), .A2(new_n1009), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1202), .A2(KEYINPUT114), .A3(new_n1006), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1198), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n994), .B1(new_n1185), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n992), .A2(KEYINPUT126), .A3(new_n984), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n983), .A2(G1986), .A3(G290), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT48), .Z(new_n1211));
  NAND2_X1  g786(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(KEYINPUT126), .B1(new_n992), .B2(new_n984), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n986), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n984), .B1(new_n1215), .B2(new_n799), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT46), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1217), .B1(new_n984), .B2(new_n987), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n983), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1216), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT47), .Z(new_n1221));
  INV_X1    g796(.A(new_n989), .ZN(new_n1222));
  OAI22_X1  g797(.A1(new_n1222), .A2(new_n990), .B1(G2067), .B2(new_n754), .ZN(new_n1223));
  AOI211_X1 g798(.A(new_n1214), .B(new_n1221), .C1(new_n984), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1208), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g800(.A1(new_n899), .A2(new_n901), .ZN(new_n1227));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n1228));
  NAND2_X1  g802(.A1(new_n672), .A2(G319), .ZN(new_n1229));
  OAI21_X1  g803(.A(new_n1228), .B1(G401), .B2(new_n1229), .ZN(new_n1230));
  NAND4_X1  g804(.A1(new_n652), .A2(new_n672), .A3(KEYINPUT127), .A4(G319), .ZN(new_n1231));
  AOI21_X1  g805(.A(G229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n1232), .A2(new_n967), .A3(new_n970), .ZN(new_n1233));
  NOR2_X1   g807(.A1(new_n1227), .A2(new_n1233), .ZN(G308));
  OR2_X1    g808(.A1(new_n1227), .A2(new_n1233), .ZN(G225));
endmodule


