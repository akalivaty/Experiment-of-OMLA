//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1332, new_n1333,
    new_n1334, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1388, new_n1389,
    new_n1390;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n210), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n213), .B1(new_n216), .B2(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n202), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n238), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G223), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G222), .A3(new_n251), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n250), .A2(G77), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n214), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT66), .B1(new_n258), .B2(new_n214), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT66), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n263), .A2(new_n264), .A3(G1), .A4(G13), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n267));
  XOR2_X1   g0067(.A(KEYINPUT67), .B(G226), .Z(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n267), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n262), .A2(new_n270), .A3(G274), .A4(new_n265), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(G200), .B1(new_n261), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n214), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  INV_X1    g0079(.A(G58), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT8), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n246), .A2(G20), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n276), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n275), .B1(new_n207), .B2(G20), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(G50), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n286), .A2(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n260), .A2(G190), .A3(new_n271), .A4(new_n269), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n273), .A2(new_n294), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT71), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT72), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT10), .B1(new_n298), .B2(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(KEYINPUT72), .B(KEYINPUT10), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n284), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n305), .A2(new_n202), .B1(new_n208), .B2(G68), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n208), .A2(G33), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n275), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n289), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT12), .ZN(new_n315));
  INV_X1    g0115(.A(new_n287), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n240), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n287), .A2(KEYINPUT12), .A3(G68), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n314), .A2(new_n240), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n310), .A2(new_n311), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n313), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n262), .A2(G238), .A3(new_n265), .A4(new_n267), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G226), .A2(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(G232), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(G1698), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n254), .B1(G33), .B2(G97), .ZN(new_n327));
  INV_X1    g0127(.A(new_n259), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n271), .B(new_n323), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT13), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT14), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(G169), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n329), .A2(KEYINPUT13), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(KEYINPUT13), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(G179), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n331), .B1(new_n330), .B2(G169), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n322), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(G200), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n321), .C1(new_n340), .C2(new_n330), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G20), .A2(G77), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT15), .B(G87), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n344), .B1(new_n277), .B2(new_n305), .C1(new_n307), .C2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n346), .A2(new_n275), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n316), .A2(new_n308), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n314), .B2(new_n308), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n254), .A2(G232), .A3(new_n251), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT69), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT69), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n254), .A2(new_n353), .A3(G232), .A4(new_n251), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OR2_X1    g0155(.A1(KEYINPUT70), .A2(G107), .ZN(new_n356));
  NAND2_X1  g0156(.A1(KEYINPUT70), .A2(G107), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n252), .A2(G238), .B1(new_n250), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n328), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n266), .A2(G244), .A3(new_n267), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n271), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n350), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OR3_X1    g0165(.A1(new_n360), .A2(G179), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(G200), .B1(new_n360), .B2(new_n362), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n350), .C1(new_n363), .C2(new_n340), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n261), .A2(new_n272), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n292), .C1(G169), .C2(new_n371), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n304), .A2(new_n343), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G159), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT74), .B1(new_n305), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n284), .A2(new_n380), .A3(G159), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n280), .A2(new_n240), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n201), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n254), .B2(G20), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n248), .A2(G33), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT7), .B(new_n208), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n387), .B1(new_n393), .B2(G68), .ZN(new_n394));
  AOI211_X1 g0194(.A(KEYINPUT73), .B(new_n240), .C1(new_n389), .C2(new_n392), .ZN(new_n395));
  OAI211_X1 g0195(.A(KEYINPUT16), .B(new_n386), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT7), .B1(new_n250), .B2(new_n208), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n388), .B(G20), .C1(new_n247), .C2(new_n249), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n402), .A3(new_n275), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n278), .A2(new_n281), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(new_n289), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n287), .B2(new_n404), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT75), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n403), .A2(KEYINPUT75), .A3(new_n407), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n254), .A2(G226), .A3(G1698), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n247), .A2(new_n249), .A3(G223), .A4(new_n251), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G87), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n259), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT76), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(KEYINPUT76), .A3(new_n259), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n262), .A2(G232), .A3(new_n265), .A4(new_n267), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n271), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(G179), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n416), .A2(new_n271), .A3(new_n421), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n420), .A2(new_n423), .B1(new_n424), .B2(new_n364), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n410), .A2(new_n411), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT18), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n410), .A2(new_n428), .A3(new_n411), .A4(new_n425), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n422), .A2(G190), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n418), .A2(new_n419), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G200), .ZN(new_n432));
  INV_X1    g0232(.A(new_n416), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n422), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n403), .A2(new_n407), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n403), .A2(new_n435), .A3(KEYINPUT17), .A4(new_n407), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n427), .A2(new_n429), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n377), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n207), .A2(G45), .ZN(new_n444));
  OR2_X1    g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(G274), .A3(new_n262), .A4(new_n265), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  INV_X1    g0250(.A(new_n446), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n453), .A2(new_n262), .A3(G270), .A4(new_n265), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n247), .A2(new_n249), .A3(G264), .A4(G1698), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n247), .A2(new_n249), .A3(G257), .A4(new_n251), .ZN(new_n457));
  INV_X1    g0257(.A(G303), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n254), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n259), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n207), .A2(G33), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n287), .A2(new_n461), .A3(new_n214), .A4(new_n274), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G116), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n207), .A2(new_n465), .A3(G13), .A4(G20), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n466), .B(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n274), .A2(new_n214), .B1(G20), .B2(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n470), .B(new_n208), .C1(G33), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(KEYINPUT20), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT20), .B1(new_n469), .B2(new_n472), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n464), .B(new_n468), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n460), .A2(KEYINPUT81), .A3(G179), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT81), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n459), .A2(new_n259), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(G179), .A3(new_n448), .A4(new_n454), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n466), .A2(new_n467), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n466), .A2(new_n467), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n481), .A2(new_n482), .B1(new_n462), .B2(new_n465), .ZN(new_n483));
  INV_X1    g0283(.A(new_n475), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n473), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n478), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n448), .A2(new_n454), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n479), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT21), .A3(G169), .A4(new_n476), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n477), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n477), .A2(new_n486), .A3(new_n489), .A4(KEYINPUT82), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n460), .A2(new_n485), .A3(new_n364), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n494), .A2(KEYINPUT21), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n476), .B1(new_n488), .B2(G200), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n340), .B2(new_n488), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(new_n493), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G107), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G20), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G13), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G1), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT25), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n462), .A2(new_n500), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g0308(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n254), .A2(new_n509), .A3(new_n208), .A4(G87), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n247), .A2(new_n249), .A3(new_n208), .A4(G87), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT83), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(KEYINPUT22), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT23), .B1(new_n358), .B2(new_n208), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT23), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n502), .A2(new_n516), .B1(new_n282), .B2(G116), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n510), .A2(new_n514), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT24), .ZN(new_n519));
  OAI22_X1  g0319(.A1(KEYINPUT23), .A2(new_n501), .B1(new_n307), .B2(new_n465), .ZN(new_n520));
  INV_X1    g0320(.A(new_n357), .ZN(new_n521));
  NOR2_X1   g0321(.A1(KEYINPUT70), .A2(G107), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G20), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n520), .B1(new_n524), .B2(KEYINPUT23), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT24), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n525), .A2(new_n526), .A3(new_n514), .A4(new_n510), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n508), .B1(new_n528), .B2(new_n275), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n266), .A2(new_n530), .A3(G264), .A4(new_n453), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n453), .A2(new_n262), .A3(G264), .A4(new_n265), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT84), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n254), .A2(G257), .A3(G1698), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n254), .A2(G250), .A3(new_n251), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G294), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n259), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n340), .A2(new_n534), .A3(new_n448), .A4(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n531), .A2(new_n533), .B1(new_n259), .B2(new_n538), .ZN(new_n541));
  AOI21_X1  g0341(.A(G200), .B1(new_n541), .B2(new_n448), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n529), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n448), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n247), .A2(new_n249), .A3(G244), .A4(new_n251), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n470), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n544), .B1(new_n550), .B2(new_n259), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n453), .A2(new_n262), .A3(G257), .A4(new_n265), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT78), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n553), .A3(new_n372), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n462), .A2(G97), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G97), .B2(new_n316), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n555), .B(KEYINPUT77), .C1(G97), .C2(new_n316), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n561), .A2(new_n471), .A3(G107), .ZN(new_n562));
  XNOR2_X1  g0362(.A(G97), .B(G107), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n564), .A2(new_n208), .B1(new_n308), .B2(new_n305), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n523), .B1(new_n389), .B2(new_n392), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n275), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n551), .A2(new_n553), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n554), .B(new_n568), .C1(new_n569), .C2(G169), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(new_n561), .ZN(new_n571));
  INV_X1    g0371(.A(new_n562), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n393), .A2(new_n358), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n275), .B1(new_n558), .B2(new_n559), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n551), .A2(new_n553), .A3(G190), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n578), .C1(new_n569), .C2(new_n432), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n543), .A2(new_n570), .A3(new_n579), .ZN(new_n580));
  AND4_X1   g0380(.A1(G179), .A2(new_n534), .A3(new_n448), .A4(new_n539), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n364), .B1(new_n541), .B2(new_n448), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n276), .B1(new_n519), .B2(new_n527), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n581), .A2(new_n582), .B1(new_n583), .B2(new_n508), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n247), .A2(new_n249), .A3(G244), .A4(G1698), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n247), .A2(new_n249), .A3(G238), .A4(new_n251), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G116), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n259), .ZN(new_n589));
  AOI21_X1  g0389(.A(G250), .B1(new_n207), .B2(G45), .ZN(new_n590));
  INV_X1    g0390(.A(G274), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n450), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n266), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n259), .A2(new_n588), .B1(new_n266), .B2(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G190), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G87), .A2(G97), .ZN(new_n599));
  NAND3_X1  g0399(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n523), .A2(new_n599), .B1(new_n208), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n247), .A2(new_n249), .A3(new_n208), .A4(G68), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT19), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n307), .B2(new_n471), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT79), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n356), .A2(new_n599), .A3(new_n357), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n600), .A2(new_n208), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT79), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n602), .A4(new_n604), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n275), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n345), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(new_n287), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n463), .A2(G87), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n589), .A2(new_n593), .A3(new_n372), .ZN(new_n618));
  AOI21_X1  g0418(.A(G169), .B1(new_n589), .B2(new_n593), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n463), .A2(new_n613), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n612), .A2(new_n621), .A3(new_n615), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n598), .A2(new_n617), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n584), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n580), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n443), .A2(new_n499), .A3(new_n625), .ZN(G372));
  INV_X1    g0426(.A(KEYINPUT88), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n304), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT88), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n408), .A2(new_n425), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT18), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n341), .A2(new_n366), .A3(new_n365), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n338), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n440), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n375), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n443), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n620), .A2(new_n622), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n597), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n609), .A2(new_n602), .A3(new_n604), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n276), .B1(new_n642), .B2(KEYINPUT79), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n614), .B1(new_n643), .B2(new_n611), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n596), .B2(new_n432), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n594), .A2(KEYINPUT85), .A3(G200), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n644), .A2(new_n646), .A3(new_n647), .A4(new_n616), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT86), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n641), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n617), .A2(KEYINPUT86), .A3(new_n646), .A4(new_n647), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n640), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n543), .A2(new_n570), .A3(new_n579), .ZN(new_n653));
  INV_X1    g0453(.A(new_n490), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n495), .A3(new_n584), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT87), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n620), .A2(new_n622), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n620), .B2(new_n622), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n551), .A2(new_n553), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n662), .A2(new_n364), .B1(new_n567), .B2(new_n560), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n644), .A2(new_n616), .A3(new_n595), .A4(new_n597), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n639), .A4(new_n554), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n648), .A2(new_n649), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n651), .A3(new_n597), .ZN(new_n669));
  INV_X1    g0469(.A(new_n570), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n639), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n667), .B1(new_n671), .B2(new_n666), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n661), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n637), .B1(new_n638), .B2(new_n673), .ZN(G369));
  NAND2_X1  g0474(.A1(new_n654), .A2(new_n495), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n504), .A2(new_n208), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n485), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n498), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n584), .A2(new_n682), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT90), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n534), .A2(new_n448), .A3(new_n539), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G169), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n541), .A2(G179), .A3(new_n448), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n528), .A2(new_n275), .ZN(new_n694));
  INV_X1    g0494(.A(new_n508), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n543), .B1(new_n529), .B2(new_n682), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n690), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n688), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n492), .A2(new_n495), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n681), .B1(new_n700), .B2(new_n493), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n698), .A2(new_n701), .B1(new_n696), .B2(new_n682), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n211), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n607), .A2(G116), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n218), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT92), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n664), .A2(new_n639), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n696), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n432), .B1(new_n551), .B2(new_n553), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n568), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n578), .A2(new_n716), .B1(new_n663), .B2(new_n554), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(new_n543), .A4(new_n682), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n712), .B1(new_n718), .B2(new_n498), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n499), .A2(new_n625), .A3(KEYINPUT92), .A4(new_n682), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n682), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n460), .A2(G179), .A3(new_n596), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n662), .A3(new_n691), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n596), .A2(new_n487), .A3(G179), .A4(new_n479), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n569), .A2(new_n728), .A3(KEYINPUT30), .A4(new_n541), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n569), .A2(new_n728), .A3(new_n541), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n724), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n534), .A2(new_n539), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n662), .A2(new_n727), .A3(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n736), .A2(KEYINPUT91), .A3(KEYINPUT30), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT91), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n731), .B2(new_n732), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n730), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n681), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n734), .B1(new_n741), .B2(new_n722), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n711), .B1(new_n721), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n673), .B2(new_n681), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n660), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n492), .A2(new_n493), .A3(new_n495), .A4(new_n584), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT93), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n653), .B(new_n652), .C1(new_n748), .C2(KEYINPUT93), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(KEYINPUT29), .A3(new_n682), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n743), .B1(new_n745), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n710), .B1(new_n754), .B2(G1), .ZN(G364));
  NOR2_X1   g0555(.A1(new_n503), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n207), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n705), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n688), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n686), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n214), .B1(G20), .B2(new_n364), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT95), .B1(new_n372), .B2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n208), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n372), .A2(KEYINPUT95), .A3(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n340), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT96), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT96), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G87), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n208), .A2(G190), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n372), .A3(new_n432), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT32), .B1(new_n777), .B2(new_n378), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n777), .A2(KEYINPUT32), .A3(new_n378), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n208), .A2(new_n372), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G190), .A3(new_n432), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n254), .B1(new_n781), .B2(new_n280), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n779), .B(new_n782), .C1(G68), .C2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n372), .A2(new_n432), .A3(G190), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n471), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n783), .A2(new_n340), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G50), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n776), .A2(G179), .A3(new_n432), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n308), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n768), .A2(G190), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(G107), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n775), .A2(new_n778), .A3(new_n785), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n784), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT33), .B(G317), .Z(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G326), .B2(new_n790), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n788), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n781), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n254), .B(new_n802), .C1(G322), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n792), .ZN(new_n805));
  INV_X1    g0605(.A(new_n777), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n805), .A2(G311), .B1(new_n806), .B2(G329), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n800), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  INV_X1    g0609(.A(new_n794), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n810), .C1(new_n458), .C2(new_n773), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n764), .B1(new_n796), .B2(new_n811), .ZN(new_n812));
  OR3_X1    g0612(.A1(KEYINPUT94), .A2(G13), .A3(G33), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT94), .B1(G13), .B2(G33), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G20), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n763), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n704), .A2(new_n250), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G355), .B1(new_n465), .B2(new_n704), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n704), .A2(new_n254), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(G45), .B2(new_n218), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n244), .A2(new_n449), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n762), .B(new_n812), .C1(new_n818), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n817), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n686), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n761), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n816), .A2(new_n764), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n759), .B1(G77), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n790), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n797), .A2(new_n835), .B1(new_n836), .B2(new_n781), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n834), .B(new_n837), .C1(G159), .C2(new_n805), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n794), .A2(G68), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n254), .B1(new_n788), .B2(new_n280), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G132), .B2(new_n806), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n773), .A2(new_n202), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n773), .A2(new_n500), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n254), .B(new_n789), .C1(G294), .C2(new_n803), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n794), .A2(G87), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n784), .A2(G283), .B1(new_n806), .B2(G311), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n790), .A2(G303), .B1(new_n805), .B2(G116), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n844), .A2(new_n845), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n831), .B1(new_n852), .B2(new_n763), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n681), .B1(new_n347), .B2(new_n349), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n369), .A2(new_n854), .B1(new_n365), .B2(new_n366), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n365), .A2(new_n366), .A3(new_n682), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n853), .B1(new_n858), .B2(new_n816), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT97), .B1(new_n855), .B2(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n369), .A2(new_n854), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n367), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT97), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n856), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n673), .B2(new_n681), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n370), .A2(new_n681), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n661), .B2(new_n672), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n743), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n762), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n873), .A2(KEYINPUT98), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n870), .A2(new_n743), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n873), .B2(KEYINPUT98), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n860), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(G384));
  AOI211_X1 g0679(.A(new_n465), .B(new_n216), .C1(new_n573), .C2(KEYINPUT35), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(KEYINPUT35), .B2(new_n573), .ZN(new_n881));
  XNOR2_X1  g0681(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n881), .B(new_n882), .ZN(new_n883));
  OR3_X1    g0683(.A1(new_n218), .A2(new_n308), .A3(new_n383), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n239), .B(KEYINPUT100), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n207), .B(G13), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n856), .B(KEYINPUT101), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n869), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n869), .A2(KEYINPUT102), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n396), .A2(new_n275), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n393), .A2(new_n387), .A3(G68), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT16), .B1(new_n898), .B2(new_n386), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n407), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n679), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n442), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n385), .B1(new_n896), .B2(new_n897), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n276), .B1(new_n906), .B2(KEYINPUT16), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n386), .B1(new_n394), .B2(new_n395), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n401), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n406), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n436), .B1(new_n910), .B2(new_n679), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n900), .A2(new_n425), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT37), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n410), .A2(new_n411), .A3(new_n901), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n436), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n426), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n905), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n904), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n442), .A2(new_n903), .B1(new_n917), .B2(new_n913), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n920), .B2(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n322), .A2(new_n681), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n338), .A2(new_n341), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n338), .B2(new_n341), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n894), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n632), .A2(new_n679), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n440), .B1(KEYINPUT18), .B2(new_n426), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n902), .B1(new_n929), .B2(new_n429), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n913), .A2(new_n917), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n905), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n410), .A2(new_n411), .A3(new_n901), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n631), .A2(new_n436), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT37), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n917), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n632), .B2(new_n440), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n426), .A2(new_n914), .A3(new_n916), .ZN(new_n940));
  INV_X1    g0740(.A(new_n408), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n941), .A2(new_n435), .B1(new_n900), .B2(new_n901), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n900), .A2(new_n425), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n915), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT38), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT103), .B1(new_n945), .B2(new_n930), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT103), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n904), .A2(new_n918), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n939), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n933), .B1(new_n949), .B2(KEYINPUT39), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n338), .A2(new_n681), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n927), .B(new_n928), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n745), .A2(new_n753), .A3(new_n443), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n637), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n858), .B1(new_n923), .B2(new_n924), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n726), .A2(new_n729), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT91), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n731), .A2(new_n738), .A3(new_n732), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT104), .B1(new_n961), .B2(new_n724), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT104), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n740), .A2(new_n963), .A3(new_n723), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n962), .A2(new_n964), .B1(new_n741), .B2(new_n722), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n957), .B1(new_n965), .B2(new_n721), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT105), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n937), .A2(new_n938), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n905), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n904), .A2(new_n947), .A3(new_n918), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n947), .B1(new_n904), .B2(new_n918), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT40), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n966), .B2(KEYINPUT105), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n967), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n921), .A2(new_n966), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n973), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n721), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n962), .A2(new_n964), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n741), .A2(new_n722), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n443), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n978), .A2(new_n983), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n984), .A2(new_n985), .A3(new_n711), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n956), .A2(new_n986), .B1(new_n207), .B2(new_n756), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n956), .A2(new_n986), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n887), .B1(new_n987), .B2(new_n988), .ZN(G367));
  OAI21_X1  g0789(.A(new_n818), .B1(new_n211), .B2(new_n345), .ZN(new_n990));
  INV_X1    g0790(.A(new_n821), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n234), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n759), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n774), .A2(G58), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n794), .A2(G77), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n254), .B1(new_n781), .B2(new_n835), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G68), .B2(new_n787), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n797), .A2(new_n378), .B1(new_n833), .B2(new_n777), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n832), .A2(new_n836), .B1(new_n792), .B2(new_n202), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n994), .A2(new_n995), .A3(new_n997), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n774), .A2(G116), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT46), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1002), .A2(new_n1003), .B1(G294), .B2(new_n784), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT113), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n254), .B1(new_n787), .B2(new_n358), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1008), .B1(new_n809), .B2(new_n792), .C1(new_n1009), .C2(new_n777), .ZN(new_n1010));
  INV_X1    g0810(.A(G311), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n832), .A2(new_n1011), .B1(new_n458), .B2(new_n781), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1012), .A2(KEYINPUT112), .B1(new_n810), .B2(new_n471), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1010), .B(new_n1013), .C1(KEYINPUT112), .C2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1001), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n993), .B1(new_n1017), .B2(new_n763), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n617), .A2(new_n682), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT106), .Z(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n660), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1023), .A2(KEYINPUT107), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n652), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(KEYINPUT107), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(new_n826), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1018), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT45), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n702), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n717), .B1(new_n577), .B2(new_n682), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT108), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n670), .A2(new_n681), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1030), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n702), .A2(new_n1036), .A3(KEYINPUT45), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1031), .A2(new_n1037), .A3(KEYINPUT44), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT44), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n702), .B2(new_n1036), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n699), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT110), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1045), .A2(KEYINPUT110), .A3(new_n1046), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1040), .A2(new_n699), .A3(new_n1044), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n698), .A2(new_n701), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT111), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n688), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n687), .A2(new_n1054), .A3(new_n1053), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n698), .A2(new_n701), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1058), .B(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n754), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n754), .B1(new_n1052), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n705), .B(KEYINPUT41), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n758), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n699), .A2(new_n1037), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1036), .A2(new_n698), .A3(new_n701), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT42), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n570), .B1(new_n1034), .B2(new_n584), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n682), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(KEYINPUT42), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT109), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1027), .B(KEYINPUT43), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(KEYINPUT109), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1027), .A2(KEYINPUT43), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1066), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1079), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1066), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n1082), .A3(new_n1076), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1029), .B1(new_n1065), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT114), .Z(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(G387));
  AOI21_X1  g0887(.A(new_n706), .B1(new_n1061), .B2(new_n754), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n754), .B2(new_n1061), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n698), .A2(new_n826), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n821), .B1(new_n231), .B2(new_n449), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n819), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n707), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n277), .A2(G50), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT50), .ZN(new_n1095));
  AOI21_X1  g0895(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n707), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1093), .A2(new_n1097), .B1(new_n500), .B2(new_n704), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n818), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n759), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n254), .B1(new_n792), .B2(new_n240), .C1(new_n202), .C2(new_n781), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n613), .A2(new_n787), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n835), .B2(new_n777), .C1(new_n832), .C2(new_n378), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n404), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1101), .B(new_n1103), .C1(new_n1104), .C2(new_n784), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n471), .B2(new_n810), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n773), .A2(new_n308), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT115), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n254), .B1(new_n806), .B2(G326), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G322), .A2(new_n790), .B1(new_n803), .B2(G317), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n458), .B2(new_n792), .C1(new_n1011), .C2(new_n797), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT48), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n809), .B2(new_n788), .C1(new_n801), .C2(new_n773), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT49), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1110), .B1(new_n465), .B2(new_n810), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1109), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT116), .Z(new_n1119));
  AOI21_X1  g0919(.A(new_n1100), .B1(new_n1119), .B2(new_n763), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1061), .A2(new_n758), .B1(new_n1090), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1089), .A2(new_n1121), .ZN(G393));
  NAND3_X1  g0922(.A1(new_n1047), .A2(new_n1051), .A3(new_n758), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n818), .B1(new_n471), .B2(new_n211), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n991), .A2(new_n238), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n759), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n788), .A2(new_n308), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G50), .B2(new_n784), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n277), .B2(new_n792), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n250), .B(new_n1129), .C1(G143), .C2(new_n806), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n832), .A2(new_n835), .B1(new_n378), .B2(new_n781), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT51), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1133), .A2(new_n848), .A3(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1130), .B(new_n1135), .C1(new_n240), .C2(new_n773), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n773), .A2(new_n809), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n784), .A2(G303), .B1(G116), .B2(new_n787), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n801), .B2(new_n792), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n254), .B(new_n1139), .C1(G322), .C2(new_n806), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n832), .A2(new_n1009), .B1(new_n1011), .B2(new_n781), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT52), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1141), .A2(new_n1142), .B1(G107), .B2(new_n794), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1140), .B(new_n1143), .C1(new_n1142), .C2(new_n1141), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1136), .B1(new_n1137), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1126), .B1(new_n1145), .B2(new_n763), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1036), .B2(new_n826), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1123), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT117), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT117), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1123), .A2(new_n1150), .A3(new_n1147), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n754), .A2(new_n1061), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n705), .B1(new_n1052), .B2(new_n1062), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(G390));
  AOI21_X1  g0955(.A(new_n926), .B1(new_n743), .B2(new_n858), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n711), .B(new_n957), .C1(new_n965), .C2(new_n721), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT102), .B1(new_n869), .B2(new_n889), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT26), .B1(new_n652), .B2(new_n670), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n656), .B(new_n660), .C1(new_n1159), .C2(new_n667), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n891), .B(new_n888), .C1(new_n1160), .C2(new_n868), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1156), .A2(new_n1157), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n748), .A2(KEYINPUT93), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1163), .A2(new_n653), .A3(new_n652), .A4(new_n749), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n681), .B1(new_n1164), .B2(new_n747), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n857), .B1(new_n1165), .B2(new_n863), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n743), .A2(new_n858), .A3(new_n926), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n711), .B(new_n866), .C1(new_n965), .C2(new_n721), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1166), .B(new_n1167), .C1(new_n1168), .C2(new_n926), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT118), .ZN(new_n1171));
  OAI211_X1 g0971(.A(G330), .B(new_n443), .C1(new_n979), .C2(new_n982), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n953), .A2(new_n1172), .A3(new_n637), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1171), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n752), .A2(new_n682), .A3(new_n863), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n856), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n866), .ZN(new_n1178));
  OAI211_X1 g0978(.A(G330), .B(new_n1178), .C1(new_n979), .C2(new_n982), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1177), .B1(new_n1179), .B2(new_n925), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n957), .ZN(new_n1181));
  OAI211_X1 g0981(.A(G330), .B(new_n1181), .C1(new_n979), .C2(new_n982), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n858), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n711), .B(new_n1183), .C1(new_n721), .C2(new_n742), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1184), .B2(new_n926), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1180), .A2(new_n1167), .B1(new_n1185), .B2(new_n894), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT118), .B1(new_n1186), .B2(new_n1173), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n926), .B1(new_n1161), .B2(new_n1158), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n951), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n950), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1177), .A2(new_n926), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n972), .A3(new_n951), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1167), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1182), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1175), .B(new_n1187), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT39), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n972), .A2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1197), .A2(new_n933), .B1(new_n951), .B2(new_n1188), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1192), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1157), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n932), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1196), .B2(new_n972), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n951), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n894), .B2(new_n926), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1167), .B(new_n1192), .C1(new_n1202), .C2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1171), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1206));
  AOI211_X1 g1006(.A(KEYINPUT118), .B(new_n1173), .C1(new_n1162), .C2(new_n1169), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1200), .B(new_n1205), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1195), .A2(new_n1208), .A3(new_n705), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n949), .A2(new_n1203), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n950), .A2(new_n1189), .B1(new_n1210), .B2(new_n1191), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1205), .B(new_n758), .C1(new_n1182), .C2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n759), .B1(new_n1104), .B2(new_n830), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n254), .B(new_n1127), .C1(G116), .C2(new_n803), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n797), .A2(new_n523), .B1(new_n777), .B2(new_n801), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n832), .A2(new_n809), .B1(new_n792), .B2(new_n471), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n775), .A2(new_n841), .A3(new_n1214), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n790), .A2(G128), .ZN(new_n1219));
  INV_X1    g1019(.A(G132), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n254), .C1(new_n1220), .C2(new_n781), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(KEYINPUT54), .B(G143), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n805), .A2(new_n1223), .B1(new_n806), .B2(G125), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n833), .B2(new_n797), .C1(new_n378), .C2(new_n788), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1221), .B(new_n1225), .C1(G50), .C2(new_n794), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT53), .B1(new_n773), .B2(new_n835), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n773), .A2(KEYINPUT53), .A3(new_n835), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1218), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1213), .B1(new_n1230), .B2(new_n763), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1202), .B2(new_n816), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1212), .A2(KEYINPUT119), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT119), .B1(new_n1212), .B2(new_n1232), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1209), .B1(new_n1233), .B2(new_n1234), .ZN(G378));
  XNOR2_X1  g1035(.A(new_n1173), .B(KEYINPUT124), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1187), .A2(new_n1175), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n711), .B1(new_n976), .B2(new_n973), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n975), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n630), .A2(new_n374), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n295), .A2(new_n679), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT55), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1247));
  INV_X1    g1047(.A(new_n1245), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n630), .A2(new_n374), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1247), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1248), .B1(new_n630), .B2(new_n374), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n375), .B(new_n1245), .C1(new_n628), .C2(new_n629), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1250), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1242), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n921), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n928), .B1(new_n1188), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1203), .B2(new_n1202), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1241), .A2(new_n975), .A3(new_n1255), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1241), .A2(new_n975), .A3(new_n1255), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1255), .B1(new_n1241), .B2(new_n975), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n952), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(new_n1265), .A3(KEYINPUT57), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n705), .B1(new_n1240), .B2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1205), .B1(new_n1211), .B2(new_n1182), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1236), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT57), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1262), .A2(new_n1265), .A3(new_n758), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n759), .B1(G50), .B2(new_n830), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G33), .A2(G41), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT120), .Z(new_n1277));
  OAI211_X1 g1077(.A(new_n1277), .B(new_n202), .C1(G41), .C2(new_n254), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n805), .A2(new_n613), .B1(new_n806), .B2(G283), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1279), .B1(new_n471), .B2(new_n797), .C1(new_n465), .C2(new_n832), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n810), .A2(new_n280), .ZN(new_n1281));
  AOI211_X1 g1081(.A(G41), .B(new_n254), .C1(new_n803), .C2(G107), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n240), .B2(new_n788), .ZN(new_n1283));
  NOR4_X1   g1083(.A1(new_n1107), .A2(new_n1280), .A3(new_n1281), .A4(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1278), .B1(new_n1284), .B2(KEYINPUT58), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT121), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(KEYINPUT58), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(G132), .A2(new_n784), .B1(new_n803), .B2(G128), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n790), .A2(G125), .B1(G150), .B2(new_n787), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1288), .B(new_n1289), .C1(new_n833), .C2(new_n792), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n774), .B2(new_n1223), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT59), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1277), .B1(G124), .B2(new_n806), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n810), .B2(new_n378), .ZN(new_n1296));
  XOR2_X1   g1096(.A(new_n1296), .B(KEYINPUT122), .Z(new_n1297));
  NAND3_X1  g1097(.A1(new_n1293), .A2(new_n1294), .A3(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1286), .A2(new_n1287), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1275), .B1(new_n1299), .B2(new_n763), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1256), .B2(new_n816), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1274), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1273), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(G375));
  NAND2_X1  g1105(.A1(new_n1186), .A2(new_n1173), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1268), .A2(new_n1064), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n925), .A2(new_n815), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n759), .B1(G68), .B2(new_n830), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n784), .A2(new_n1223), .B1(new_n803), .B2(G137), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1220), .B2(new_n832), .ZN(new_n1311));
  OAI22_X1  g1111(.A1(new_n788), .A2(new_n202), .B1(new_n792), .B2(new_n835), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n250), .B(new_n1312), .C1(G128), .C2(new_n806), .ZN(new_n1313));
  OAI221_X1 g1113(.A(new_n1313), .B1(new_n280), .B2(new_n810), .C1(new_n773), .C2(new_n378), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1311), .B1(new_n1314), .B2(KEYINPUT126), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(KEYINPUT126), .B2(new_n1314), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n790), .A2(G294), .B1(new_n806), .B2(G303), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n254), .B1(new_n803), .B2(G283), .ZN(new_n1318));
  AND4_X1   g1118(.A1(new_n995), .A2(new_n1317), .A3(new_n1102), .A4(new_n1318), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n784), .A2(G116), .B1(new_n805), .B2(new_n358), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(KEYINPUT125), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1319), .B(new_n1321), .C1(new_n773), .C2(new_n471), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1316), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1309), .B1(new_n1323), .B2(new_n763), .ZN(new_n1324));
  AOI22_X1  g1124(.A1(new_n1170), .A2(new_n758), .B1(new_n1308), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1307), .A2(new_n1325), .ZN(G381));
  AND2_X1   g1126(.A1(new_n1212), .A2(new_n1232), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1209), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1089), .A2(new_n1121), .A3(new_n828), .ZN(new_n1329));
  NOR4_X1   g1129(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1086), .A2(new_n1304), .A3(new_n1328), .A4(new_n1330), .ZN(G407));
  NAND2_X1  g1131(.A1(new_n680), .A2(G213), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1304), .A2(new_n1328), .A3(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(G407), .A2(new_n1334), .A3(G213), .ZN(G409));
  INV_X1    g1135(.A(new_n1085), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G393), .A2(G396), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1329), .ZN(new_n1338));
  AOI21_X1  g1138(.A(G390), .B1(new_n1338), .B2(KEYINPUT114), .ZN(new_n1339));
  OR2_X1    g1139(.A1(new_n1154), .A2(new_n1153), .ZN(new_n1340));
  AOI22_X1  g1140(.A1(new_n1340), .A2(new_n1152), .B1(new_n1337), .B2(new_n1329), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1336), .B1(new_n1339), .B2(new_n1341), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1089), .A2(new_n1121), .A3(new_n828), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n828), .B1(new_n1089), .B2(new_n1121), .ZN(new_n1344));
  OAI21_X1  g1144(.A(KEYINPUT114), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(new_n1152), .A3(new_n1340), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1338), .A2(G390), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1346), .A2(new_n1085), .A3(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1342), .A2(new_n1348), .ZN(new_n1349));
  OAI211_X1 g1149(.A(G378), .B(new_n1302), .C1(new_n1267), .C2(new_n1272), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1270), .A2(new_n1271), .A3(new_n1064), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1302), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1328), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1333), .B1(new_n1350), .B2(new_n1353), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n705), .B1(new_n1355), .B2(KEYINPUT60), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1268), .A2(new_n1306), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1356), .B1(new_n1357), .B2(KEYINPUT60), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1325), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n878), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1360), .ZN(new_n1361));
  NOR3_X1   g1161(.A1(new_n1358), .A2(new_n878), .A3(new_n1359), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  AOI21_X1  g1163(.A(KEYINPUT62), .B1(new_n1354), .B2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1350), .A2(new_n1353), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT127), .B1(new_n1365), .B2(new_n1332), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT127), .ZN(new_n1367));
  AOI211_X1 g1167(.A(new_n1367), .B(new_n1333), .C1(new_n1350), .C2(new_n1353), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1366), .A2(new_n1368), .ZN(new_n1369));
  AND2_X1   g1169(.A1(new_n1363), .A2(KEYINPUT62), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1364), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1362), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1372), .A2(G2897), .A3(new_n1333), .A4(new_n1360), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1333), .A2(G2897), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1374), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1373), .A2(new_n1375), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1376), .B1(new_n1366), .B2(new_n1368), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT61), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  OAI21_X1  g1179(.A(new_n1349), .B1(new_n1371), .B2(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1354), .B1(new_n1373), .B2(new_n1375), .ZN(new_n1381));
  NOR3_X1   g1181(.A1(new_n1349), .A2(new_n1381), .A3(KEYINPUT61), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1369), .A2(KEYINPUT63), .A3(new_n1363), .ZN(new_n1383));
  AND2_X1   g1183(.A1(new_n1354), .A2(new_n1363), .ZN(new_n1384));
  OR2_X1    g1184(.A1(new_n1384), .A2(KEYINPUT63), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1382), .A2(new_n1383), .A3(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1380), .A2(new_n1386), .ZN(G405));
  INV_X1    g1187(.A(new_n1328), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1350), .B1(new_n1304), .B2(new_n1388), .ZN(new_n1389));
  XNOR2_X1  g1189(.A(new_n1389), .B(new_n1363), .ZN(new_n1390));
  XNOR2_X1  g1190(.A(new_n1390), .B(new_n1349), .ZN(G402));
endmodule


