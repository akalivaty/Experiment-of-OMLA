//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT69), .B(G128), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n188), .A2(G143), .ZN(new_n195));
  OAI22_X1  g009(.A1(new_n191), .A2(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n193), .B2(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n188), .A2(KEYINPUT65), .A3(G143), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(G146), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n199), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n203), .A2(new_n204), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n196), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G134), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G137), .ZN(new_n211));
  OAI21_X1  g025(.A(G131), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(G134), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT11), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n209), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n214), .A2(KEYINPUT11), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n207), .A2(new_n212), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  OR2_X1    g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n224), .B(new_n225), .C1(new_n194), .C2(new_n195), .ZN(new_n226));
  INV_X1    g040(.A(new_n224), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n198), .A2(new_n199), .A3(new_n202), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n210), .A2(G137), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n211), .B2(new_n218), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n213), .B1(new_n215), .B2(new_n233), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n232), .A2(new_n234), .A3(G131), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n221), .B1(new_n216), .B2(new_n220), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n230), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n223), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT70), .B1(new_n239), .B2(G119), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G116), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n240), .B(new_n243), .C1(G116), .C2(new_n242), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n238), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n248), .B(KEYINPUT28), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n232), .B2(new_n234), .ZN(new_n250));
  AOI211_X1 g064(.A(KEYINPUT67), .B(new_n229), .C1(new_n222), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n222), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n230), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n223), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n246), .ZN(new_n256));
  INV_X1    g070(.A(G237), .ZN(new_n257));
  INV_X1    g071(.A(G953), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G210), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n259), .B(KEYINPUT27), .Z(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n260), .B(new_n261), .Z(new_n262));
  NAND3_X1  g076(.A1(new_n249), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT29), .B1(new_n263), .B2(KEYINPUT75), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT69), .B(G128), .Z(new_n265));
  AOI22_X1  g079(.A1(new_n265), .A2(new_n190), .B1(new_n189), .B2(new_n202), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n203), .A2(new_n204), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n203), .A2(new_n204), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n222), .A2(new_n212), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n237), .B(KEYINPUT30), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n223), .A2(KEYINPUT71), .A3(KEYINPUT30), .A4(new_n237), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n255), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n246), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n273), .A2(new_n274), .B1(new_n255), .B2(new_n276), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT72), .A3(new_n246), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n283), .A2(new_n248), .ZN(new_n284));
  OAI221_X1 g098(.A(new_n264), .B1(KEYINPUT75), .B2(new_n263), .C1(new_n262), .C2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n238), .A2(new_n247), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n249), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n262), .A2(KEYINPUT29), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n187), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n262), .B1(new_n249), .B2(new_n256), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n248), .A2(new_n262), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT31), .B1(new_n283), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  AOI211_X1 g113(.A(new_n299), .B(new_n296), .C1(new_n280), .C2(new_n282), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n295), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n303), .B(new_n295), .C1(new_n298), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT74), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n293), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT32), .B(new_n307), .C1(new_n302), .C2(new_n304), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n292), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT22), .B(G137), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n258), .A2(G221), .A3(G234), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G125), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n319), .B1(new_n323), .B2(KEYINPUT16), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n322), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n318), .B1(new_n326), .B2(new_n316), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n188), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n200), .A2(G119), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n192), .B2(G119), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT24), .B(G110), .Z(new_n331));
  AOI22_X1  g145(.A1(new_n325), .A2(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT23), .B1(new_n200), .B2(G119), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n336), .A2(new_n337), .A3(G110), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n336), .B2(G110), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n332), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n327), .A2(new_n188), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n326), .A2(G146), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n336), .A2(G110), .B1(new_n330), .B2(new_n331), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT78), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n340), .B(new_n350), .C1(new_n346), .C2(new_n347), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n315), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n315), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n312), .B1(new_n355), .B2(G902), .ZN(new_n356));
  INV_X1    g170(.A(G902), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT25), .B(new_n357), .C1(new_n352), .C2(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G217), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(G234), .B2(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n361), .A2(G902), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n355), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n355), .A2(new_n367), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n362), .B(new_n363), .C1(new_n366), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n370), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n366), .B1(new_n373), .B2(new_n368), .ZN(new_n374));
  INV_X1    g188(.A(new_n361), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n356), .B2(new_n358), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT82), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n257), .A2(new_n258), .A3(G214), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n193), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G131), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(G143), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n221), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n341), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n323), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n326), .B(KEYINPUT85), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(new_n386), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n385), .B1(G146), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(KEYINPUT18), .A2(G131), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n391), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n388), .A2(new_n188), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n392), .B(new_n393), .C1(new_n394), .C2(new_n342), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT86), .B(G104), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n328), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT87), .B1(new_n402), .B2(new_n341), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT17), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n382), .A2(new_n384), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n381), .A2(KEYINPUT17), .A3(G131), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n325), .A2(new_n407), .A3(new_n328), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n403), .A2(new_n405), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n395), .A3(new_n399), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n401), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(G475), .A2(G902), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT89), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n418));
  INV_X1    g232(.A(new_n412), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n401), .B2(new_n410), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n420), .B2(new_n415), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n422), .A3(new_n415), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n414), .A2(new_n417), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n409), .A2(new_n395), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(new_n399), .ZN(new_n426));
  OAI21_X1  g240(.A(G475), .B1(new_n426), .B2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT9), .B(G234), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n430), .A2(new_n360), .A3(G953), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n265), .B2(new_n193), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n192), .A2(KEYINPUT90), .A3(G143), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n193), .A2(G128), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n210), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G122), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G116), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n239), .A2(G122), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G107), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G107), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT13), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n436), .B(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n433), .B2(new_n434), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n447), .B1(new_n450), .B2(new_n210), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n438), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT14), .ZN(new_n453));
  OAI21_X1  g267(.A(G107), .B1(new_n441), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n455), .B(new_n456), .C1(KEYINPUT14), .C2(new_n445), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n445), .A2(KEYINPUT14), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT91), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n459), .A3(new_n444), .ZN(new_n460));
  INV_X1    g274(.A(new_n434), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT90), .B1(new_n192), .B2(G143), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n436), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G134), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n464), .B2(new_n437), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n431), .B1(new_n452), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n437), .ZN(new_n467));
  INV_X1    g281(.A(new_n460), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n437), .B(new_n447), .C1(new_n210), .C2(new_n450), .ZN(new_n470));
  INV_X1    g284(.A(new_n431), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n472), .A3(new_n357), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n473), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(G234), .A2(G237), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(G952), .A3(new_n258), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT21), .B(G898), .Z(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT92), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n480), .A2(G902), .A3(G953), .A4(new_n477), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n476), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n429), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT10), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n198), .A2(new_n199), .A3(new_n202), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n190), .A2(G128), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n267), .A2(new_n268), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G104), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G107), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n488), .A2(G107), .ZN(new_n491));
  OAI21_X1  g305(.A(G101), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT3), .B1(new_n488), .B2(G107), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT3), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n443), .A3(G104), .ZN(new_n495));
  INV_X1    g309(.A(G101), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n493), .A2(new_n495), .A3(new_n496), .A4(new_n489), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n484), .B1(new_n487), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n495), .A3(new_n489), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G101), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n503), .A3(G101), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n230), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n498), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n207), .A2(new_n506), .A3(KEYINPUT10), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n499), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n253), .ZN(new_n509));
  INV_X1    g323(.A(new_n253), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n499), .A2(new_n510), .A3(new_n505), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G140), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT83), .ZN(new_n514));
  INV_X1    g328(.A(G227), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(G953), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n514), .B(new_n516), .Z(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n207), .A2(new_n506), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n267), .A2(new_n268), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n486), .A2(new_n485), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n498), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n253), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(KEYINPUT12), .B(new_n253), .C1(new_n520), .C2(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n511), .A2(new_n517), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G469), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n357), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n357), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(new_n511), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n518), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n529), .A2(new_n509), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n533), .B(new_n535), .C1(new_n539), .C2(new_n532), .ZN(new_n540));
  OAI21_X1  g354(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G210), .B1(G237), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n246), .A2(new_n502), .A3(new_n504), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT5), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n242), .A3(G116), .ZN(new_n549));
  OAI211_X1 g363(.A(G113), .B(new_n549), .C1(new_n244), .C2(new_n548), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n244), .A2(new_n245), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n506), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(G110), .B(G122), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n547), .A2(new_n552), .A3(new_n554), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(KEYINPUT6), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n269), .A2(new_n321), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n229), .A2(G125), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G224), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G953), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n559), .B(new_n560), .C1(new_n562), .C2(G953), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT6), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n553), .A2(new_n567), .A3(new_n555), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n558), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT7), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n561), .B1(new_n571), .B2(new_n563), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n550), .A2(new_n551), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n498), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n552), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(new_n554), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n563), .A2(new_n571), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n559), .A2(new_n560), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n572), .A2(new_n578), .A3(new_n557), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n357), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n546), .B1(new_n570), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n569), .A2(new_n357), .A3(new_n545), .A4(new_n581), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n544), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n483), .A2(new_n542), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n311), .A2(new_n379), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  AOI21_X1  g403(.A(KEYINPUT72), .B1(new_n281), .B2(new_n246), .ZN(new_n590));
  AND4_X1   g404(.A1(KEYINPUT72), .A2(new_n275), .A3(new_n246), .A4(new_n277), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n297), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n299), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n283), .A2(KEYINPUT31), .A3(new_n297), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n303), .B1(new_n595), .B2(new_n295), .ZN(new_n596));
  AOI211_X1 g410(.A(KEYINPUT73), .B(new_n294), .C1(new_n593), .C2(new_n594), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n357), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n308), .B1(new_n596), .B2(new_n597), .ZN(new_n600));
  INV_X1    g414(.A(new_n542), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n379), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT93), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n481), .A2(new_n478), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n585), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n473), .A2(new_n474), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n473), .A2(KEYINPUT96), .A3(new_n474), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT95), .B(new_n471), .C1(new_n452), .C2(new_n465), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n471), .A2(KEYINPUT95), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n469), .A2(new_n470), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(KEYINPUT33), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n466), .A2(new_n472), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n616), .A2(new_n618), .A3(G478), .A4(new_n357), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n607), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n473), .A2(KEYINPUT96), .A3(new_n474), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT96), .B1(new_n473), .B2(new_n474), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n607), .B(new_n619), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n603), .A2(new_n428), .A3(new_n606), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NAND3_X1  g442(.A1(new_n414), .A2(new_n421), .A3(new_n416), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n606), .A2(new_n427), .A3(new_n476), .A4(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n603), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n349), .A2(new_n351), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n315), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n635), .A2(new_n638), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n366), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n359), .B2(new_n361), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n542), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n585), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n483), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n599), .A3(new_n600), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT37), .B(G110), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G12));
  NOR2_X1   g464(.A1(new_n258), .A2(G900), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(G902), .A3(new_n477), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT100), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n478), .B(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n629), .A2(new_n427), .A3(new_n476), .A4(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT102), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(KEYINPUT102), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n657), .A2(new_n658), .A3(new_n585), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n643), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n656), .B(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n658), .B1(new_n663), .B2(new_n585), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n311), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(G128), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G30));
  NAND2_X1  g482(.A1(new_n583), .A2(new_n584), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT38), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n642), .A2(new_n543), .A3(new_n428), .A4(new_n476), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n655), .B(KEYINPUT39), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n601), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n671), .B(new_n672), .C1(KEYINPUT40), .C2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n262), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n284), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n248), .A2(new_n676), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n357), .B1(new_n678), .B2(new_n286), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(new_n309), .B2(new_n310), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n675), .B(new_n681), .C1(KEYINPUT40), .C2(new_n674), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  OAI211_X1 g497(.A(new_n428), .B(new_n655), .C1(new_n620), .C2(new_n624), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n644), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n311), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NAND2_X1  g501(.A1(new_n625), .A2(new_n428), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n518), .A2(new_n512), .B1(new_n528), .B2(new_n529), .ZN(new_n689));
  OAI21_X1  g503(.A(G469), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n533), .A3(new_n541), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT105), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n690), .A2(new_n533), .A3(new_n693), .A4(new_n541), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n688), .A2(new_n695), .A3(new_n605), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n311), .A2(new_n379), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT106), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n311), .A2(new_n699), .A3(new_n379), .A4(new_n696), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND2_X1  g517(.A1(new_n600), .A2(KEYINPUT32), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n305), .A2(new_n293), .A3(new_n308), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n291), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n630), .A2(new_n695), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n706), .A2(new_n378), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n239), .ZN(G18));
  INV_X1    g523(.A(new_n642), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n585), .A2(new_n541), .A3(new_n533), .A4(new_n690), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n646), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n242), .ZN(G21));
  NAND3_X1  g529(.A1(new_n692), .A2(new_n604), .A3(new_n694), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n428), .A2(new_n585), .A3(new_n476), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n428), .A2(KEYINPUT107), .A3(new_n585), .A4(new_n476), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n374), .A2(new_n376), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n595), .B1(new_n262), .B2(new_n288), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n308), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n599), .A2(new_n721), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR3_X1   g540(.A1(new_n684), .A2(new_n642), .A3(new_n711), .ZN(new_n727));
  AOI21_X1  g541(.A(G902), .B1(new_n302), .B2(new_n304), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n727), .B(new_n724), .C1(new_n187), .C2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n599), .A2(KEYINPUT108), .A3(new_n724), .A4(new_n727), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(new_n722), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n706), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n669), .A2(new_n544), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n542), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n684), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n311), .A2(new_n379), .A3(new_n741), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n744));
  AND3_X1   g558(.A1(new_n743), .A2(KEYINPUT110), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT110), .B1(new_n743), .B2(new_n744), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  NAND4_X1  g562(.A1(new_n311), .A2(new_n379), .A3(new_n663), .A4(new_n739), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n532), .B1(new_n539), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n537), .A2(KEYINPUT45), .A3(new_n538), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n534), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n533), .B1(new_n754), .B2(KEYINPUT46), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n541), .B(new_n673), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n599), .A2(new_n600), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n625), .A2(new_n429), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n625), .A2(new_n761), .A3(new_n429), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n758), .A2(new_n710), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n738), .B(new_n757), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n764), .B2(new_n763), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  OAI21_X1  g581(.A(new_n541), .B1(new_n755), .B2(new_n756), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(KEYINPUT47), .B(new_n541), .C1(new_n755), .C2(new_n756), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n379), .A2(new_n684), .A3(new_n738), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n706), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NAND2_X1  g589(.A1(new_n588), .A2(new_n647), .ZN(new_n776));
  INV_X1    g590(.A(new_n476), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n688), .B1(new_n428), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n606), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n603), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n725), .B1(new_n706), .B2(new_n713), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n708), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n783), .B1(new_n701), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n701), .A2(new_n785), .A3(new_n783), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n719), .A2(new_n720), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n655), .B(KEYINPUT113), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n601), .A2(new_n790), .A3(new_n642), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n681), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n733), .A2(new_n666), .A3(new_n686), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n731), .A2(new_n732), .B1(new_n665), .B2(new_n311), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(KEYINPUT52), .A3(new_n686), .A4(new_n793), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n749), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n598), .A2(G472), .B1(new_n308), .B2(new_n723), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n710), .A3(new_n741), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n427), .A2(new_n777), .A3(new_n629), .A4(new_n655), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n739), .A2(new_n710), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n802), .B1(new_n706), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT112), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n706), .A2(new_n804), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n749), .A4(new_n802), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n799), .A2(new_n747), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT53), .B1(new_n789), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n701), .A2(new_n783), .A3(new_n785), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n781), .B1(new_n813), .B2(new_n786), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n799), .A2(new_n810), .A3(new_n747), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n797), .A2(new_n795), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT54), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n654), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n760), .A2(new_n821), .A3(new_n762), .ZN(new_n822));
  INV_X1    g636(.A(new_n691), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n737), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n736), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT48), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n681), .A2(new_n378), .A3(new_n478), .A4(new_n824), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n428), .A3(new_n625), .ZN(new_n829));
  INV_X1    g643(.A(G952), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n599), .A2(new_n722), .A3(new_n724), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n822), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n830), .B(G953), .C1(new_n832), .C2(new_n712), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n760), .A2(new_n821), .A3(new_n762), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n823), .A2(new_n544), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n669), .B(KEYINPUT38), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n671), .A2(KEYINPUT114), .A3(new_n544), .A4(new_n823), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n835), .A2(new_n722), .A3(new_n842), .A4(new_n801), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT50), .B1(new_n843), .B2(KEYINPUT115), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n832), .A2(new_n845), .A3(new_n842), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(KEYINPUT116), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n625), .A2(new_n428), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n801), .A2(new_n710), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n828), .A2(new_n848), .B1(new_n850), .B2(new_n825), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n843), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n846), .B2(new_n844), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n690), .A2(new_n533), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n770), .B(new_n771), .C1(new_n541), .C2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n860), .A2(new_n832), .A3(new_n737), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(new_n861), .B2(KEYINPUT51), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n834), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n844), .A2(new_n846), .ZN(new_n864));
  INV_X1    g678(.A(new_n855), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n847), .A3(new_n851), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n863), .B(KEYINPUT118), .C1(KEYINPUT51), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n817), .B1(new_n814), .B2(new_n815), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n701), .A2(new_n785), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n781), .A2(KEYINPUT53), .A3(new_n816), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n811), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n868), .B1(new_n852), .B2(new_n856), .ZN(new_n878));
  INV_X1    g692(.A(new_n861), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT51), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n866), .A2(new_n862), .A3(new_n847), .A4(new_n851), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n829), .A3(new_n833), .A4(new_n827), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n877), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n820), .A2(new_n870), .A3(new_n876), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n830), .A2(new_n258), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n541), .A2(new_n543), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n859), .B2(KEYINPUT49), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(KEYINPUT49), .B2(new_n859), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n722), .A2(new_n671), .ZN(new_n890));
  OR4_X1    g704(.A1(new_n681), .A2(new_n759), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n886), .A2(KEYINPUT119), .A3(new_n891), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(G75));
  AOI21_X1  g710(.A(new_n357), .B1(new_n871), .B2(new_n874), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(G210), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n558), .A2(new_n568), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n566), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n258), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n903), .A2(new_n908), .ZN(G51));
  NAND2_X1  g723(.A1(new_n871), .A2(new_n874), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n876), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n534), .B(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n531), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n897), .A2(new_n753), .A3(new_n752), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n904), .B1(new_n915), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n410), .A3(new_n401), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(new_n411), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n905), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n919), .A2(KEYINPUT121), .A3(new_n905), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G60));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n820), .B2(new_n876), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n616), .B2(new_n618), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n616), .A2(new_n618), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n930), .B(new_n927), .C1(new_n911), .C2(new_n876), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n929), .A2(new_n904), .A3(new_n931), .ZN(G63));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT122), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT60), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n910), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n371), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n905), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n639), .A2(new_n640), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n934), .B(new_n935), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n942), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n904), .B1(new_n938), .B2(new_n371), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT122), .A4(new_n933), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n943), .A2(new_n946), .ZN(G66));
  XNOR2_X1  g761(.A(new_n814), .B(KEYINPUT123), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n258), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n480), .B2(new_n562), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n900), .B1(G898), .B2(new_n258), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  INV_X1    g767(.A(G900), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n515), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n766), .A2(new_n774), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n797), .A2(new_n686), .ZN(new_n958));
  INV_X1    g772(.A(new_n757), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n736), .A2(new_n959), .A3(new_n790), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n749), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n747), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n258), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n281), .B(new_n389), .Z(new_n965));
  XNOR2_X1  g779(.A(new_n651), .B(KEYINPUT125), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n706), .A2(new_n378), .A3(new_n740), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n673), .A3(new_n778), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n797), .A2(new_n682), .A3(new_n686), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n957), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(KEYINPUT62), .B2(new_n971), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n965), .A2(G953), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n956), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n955), .A2(KEYINPUT126), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n977), .B(new_n978), .Z(G72));
  NOR2_X1   g793(.A1(new_n948), .A2(new_n974), .ZN(new_n980));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT63), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n677), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n678), .B1(new_n280), .B2(new_n282), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n948), .A2(new_n963), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n982), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n812), .A2(new_n819), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n284), .A2(new_n262), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n990));
  AOI22_X1  g804(.A1(new_n989), .A2(KEYINPUT127), .B1(new_n283), .B2(new_n297), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n982), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n904), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n983), .A2(new_n986), .A3(new_n993), .ZN(G57));
endmodule


