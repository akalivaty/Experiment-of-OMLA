

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(n771), .ZN(n739) );
  NOR2_X2 U555 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X2 U556 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U557 ( .A1(n748), .A2(n961), .ZN(n730) );
  XNOR2_X1 U558 ( .A(KEYINPUT66), .B(n550), .ZN(n645) );
  XNOR2_X1 U559 ( .A(n793), .B(n792), .ZN(n794) );
  NAND2_X1 U560 ( .A1(n791), .A2(n790), .ZN(n793) );
  AND2_X1 U561 ( .A1(n528), .A2(n527), .ZN(n521) );
  XNOR2_X1 U562 ( .A(KEYINPUT23), .B(n531), .ZN(n522) );
  INV_X1 U563 ( .A(KEYINPUT30), .ZN(n761) );
  XNOR2_X1 U564 ( .A(n761), .B(KEYINPUT107), .ZN(n762) );
  XNOR2_X1 U565 ( .A(n763), .B(n762), .ZN(n764) );
  INV_X1 U566 ( .A(KEYINPUT64), .ZN(n792) );
  NAND2_X1 U567 ( .A1(n723), .A2(n722), .ZN(n771) );
  NAND2_X1 U568 ( .A1(G8), .A2(n771), .ZN(n806) );
  XNOR2_X1 U569 ( .A(KEYINPUT68), .B(n551), .ZN(n655) );
  NOR2_X1 U570 ( .A1(G2105), .A2(n530), .ZN(n901) );
  NOR2_X1 U571 ( .A1(G651), .A2(n645), .ZN(n664) );
  NOR2_X1 U572 ( .A1(n578), .A2(n577), .ZN(n954) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U574 ( .A(KEYINPUT17), .B(n523), .Z(n900) );
  NAND2_X1 U575 ( .A1(G137), .A2(n900), .ZN(n525) );
  INV_X1 U576 ( .A(KEYINPUT65), .ZN(n524) );
  XNOR2_X1 U577 ( .A(n525), .B(n524), .ZN(n529) );
  INV_X1 U578 ( .A(G2105), .ZN(n526) );
  INV_X1 U579 ( .A(G2104), .ZN(n530) );
  NOR2_X1 U580 ( .A1(n526), .A2(n530), .ZN(n906) );
  NAND2_X1 U581 ( .A1(G113), .A2(n906), .ZN(n528) );
  NOR2_X1 U582 ( .A1(G2104), .A2(n526), .ZN(n904) );
  NAND2_X1 U583 ( .A1(G125), .A2(n904), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n529), .A2(n521), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G101), .A2(n901), .ZN(n531) );
  NOR2_X2 U586 ( .A1(n532), .A2(n522), .ZN(G160) );
  XOR2_X1 U587 ( .A(G2443), .B(G2446), .Z(n534) );
  XNOR2_X1 U588 ( .A(G2427), .B(G2451), .ZN(n533) );
  XNOR2_X1 U589 ( .A(n534), .B(n533), .ZN(n540) );
  XOR2_X1 U590 ( .A(G2430), .B(G2454), .Z(n536) );
  XNOR2_X1 U591 ( .A(G1348), .B(G1341), .ZN(n535) );
  XNOR2_X1 U592 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U593 ( .A(G2435), .B(G2438), .Z(n537) );
  XNOR2_X1 U594 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U595 ( .A(n540), .B(n539), .Z(n541) );
  AND2_X1 U596 ( .A1(G14), .A2(n541), .ZN(G401) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U598 ( .A1(G135), .A2(n900), .ZN(n543) );
  NAND2_X1 U599 ( .A1(G111), .A2(n906), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n904), .A2(G123), .ZN(n544) );
  XOR2_X1 U602 ( .A(KEYINPUT18), .B(n544), .Z(n545) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n901), .A2(G99), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n927) );
  XNOR2_X1 U606 ( .A(G2096), .B(n927), .ZN(n549) );
  OR2_X1 U607 ( .A1(G2100), .A2(n549), .ZN(G156) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  XOR2_X1 U611 ( .A(G543), .B(KEYINPUT0), .Z(n550) );
  XNOR2_X1 U612 ( .A(KEYINPUT67), .B(G651), .ZN(n557) );
  NOR2_X1 U613 ( .A1(n645), .A2(n557), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n655), .A2(G76), .ZN(n552) );
  XNOR2_X1 U615 ( .A(KEYINPUT82), .B(n552), .ZN(n555) );
  NOR2_X1 U616 ( .A1(G543), .A2(G651), .ZN(n657) );
  NAND2_X1 U617 ( .A1(n657), .A2(G89), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT4), .B(n553), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n556), .B(KEYINPUT5), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G51), .A2(n664), .ZN(n560) );
  NOR2_X1 U622 ( .A1(G543), .A2(n557), .ZN(n558) );
  XOR2_X2 U623 ( .A(KEYINPUT1), .B(n558), .Z(n658) );
  NAND2_X1 U624 ( .A1(G63), .A2(n658), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n561), .Z(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U632 ( .A(G223), .ZN(n841) );
  NAND2_X1 U633 ( .A1(n841), .A2(G567), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT11), .ZN(n567) );
  XNOR2_X1 U635 ( .A(KEYINPUT77), .B(n567), .ZN(G234) );
  XOR2_X1 U636 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n569) );
  NAND2_X1 U637 ( .A1(G56), .A2(n658), .ZN(n568) );
  XNOR2_X1 U638 ( .A(n569), .B(n568), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n657), .A2(G81), .ZN(n570) );
  XNOR2_X1 U640 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G68), .A2(n655), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U643 ( .A(n573), .B(KEYINPUT13), .Z(n574) );
  INV_X1 U644 ( .A(n574), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G43), .A2(n664), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n954), .A2(G860), .ZN(G153) );
  NAND2_X1 U648 ( .A1(G52), .A2(n664), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G64), .A2(n658), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT72), .B(KEYINPUT9), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n655), .A2(G77), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n657), .A2(G90), .ZN(n581) );
  XOR2_X1 U654 ( .A(KEYINPUT71), .B(n581), .Z(n582) );
  NAND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U656 ( .A(n585), .B(n584), .Z(n586) );
  NOR2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U658 ( .A(KEYINPUT73), .B(n588), .Z(G171) );
  INV_X1 U659 ( .A(G171), .ZN(G301) );
  NAND2_X1 U660 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U661 ( .A1(G66), .A2(n658), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n657), .A2(G92), .ZN(n589) );
  XOR2_X1 U663 ( .A(KEYINPUT79), .B(n589), .Z(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n592), .B(KEYINPUT80), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G54), .A2(n664), .ZN(n593) );
  XNOR2_X1 U667 ( .A(KEYINPUT81), .B(n593), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n655), .A2(G79), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X2 U671 ( .A(KEYINPUT15), .B(n598), .Z(n960) );
  INV_X1 U672 ( .A(G868), .ZN(n675) );
  NAND2_X1 U673 ( .A1(n960), .A2(n675), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G53), .A2(n664), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G65), .A2(n658), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT75), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G78), .A2(n655), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n657), .A2(G91), .ZN(n606) );
  XOR2_X1 U682 ( .A(KEYINPUT74), .B(n606), .Z(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U684 ( .A(KEYINPUT76), .B(n609), .Z(G299) );
  INV_X1 U685 ( .A(G299), .ZN(n961) );
  NAND2_X1 U686 ( .A1(n961), .A2(n675), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT83), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n675), .A2(G286), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n612), .A2(n611), .ZN(G297) );
  INV_X1 U690 ( .A(G860), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n613), .A2(G559), .ZN(n614) );
  INV_X1 U692 ( .A(n960), .ZN(n731) );
  NAND2_X1 U693 ( .A1(n614), .A2(n731), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n615), .B(KEYINPUT16), .ZN(n616) );
  XNOR2_X1 U695 ( .A(KEYINPUT84), .B(n616), .ZN(G148) );
  NAND2_X1 U696 ( .A1(n954), .A2(n675), .ZN(n617) );
  XNOR2_X1 U697 ( .A(KEYINPUT85), .B(n617), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G868), .A2(n731), .ZN(n618) );
  NOR2_X1 U699 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U701 ( .A1(G80), .A2(n655), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G93), .A2(n657), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U704 ( .A(KEYINPUT88), .B(n623), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G55), .A2(n664), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G67), .A2(n658), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n676) );
  NAND2_X1 U709 ( .A1(G559), .A2(n731), .ZN(n628) );
  XNOR2_X1 U710 ( .A(n628), .B(n954), .ZN(n673) );
  XOR2_X1 U711 ( .A(n673), .B(KEYINPUT86), .Z(n629) );
  NOR2_X1 U712 ( .A1(G860), .A2(n629), .ZN(n630) );
  XOR2_X1 U713 ( .A(KEYINPUT87), .B(n630), .Z(n631) );
  XOR2_X1 U714 ( .A(n676), .B(n631), .Z(G145) );
  NAND2_X1 U715 ( .A1(G47), .A2(n664), .ZN(n632) );
  XOR2_X1 U716 ( .A(KEYINPUT70), .B(n632), .Z(n637) );
  NAND2_X1 U717 ( .A1(G72), .A2(n655), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G85), .A2(n657), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U720 ( .A(KEYINPUT69), .B(n635), .Z(n636) );
  NOR2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G60), .A2(n658), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U724 ( .A1(n664), .A2(G49), .ZN(n640) );
  XOR2_X1 U725 ( .A(KEYINPUT89), .B(n640), .Z(n642) );
  NAND2_X1 U726 ( .A1(G651), .A2(G74), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U728 ( .A1(n658), .A2(n643), .ZN(n644) );
  XNOR2_X1 U729 ( .A(n644), .B(KEYINPUT90), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G87), .A2(n645), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U732 ( .A1(G50), .A2(n664), .ZN(n649) );
  NAND2_X1 U733 ( .A1(G62), .A2(n658), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U735 ( .A(KEYINPUT92), .B(n650), .Z(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(G75), .ZN(n652) );
  NAND2_X1 U737 ( .A1(G88), .A2(n657), .ZN(n651) );
  AND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U739 ( .A1(n654), .A2(n653), .ZN(G303) );
  INV_X1 U740 ( .A(G303), .ZN(G166) );
  NAND2_X1 U741 ( .A1(n655), .A2(G73), .ZN(n656) );
  XOR2_X1 U742 ( .A(KEYINPUT2), .B(n656), .Z(n663) );
  NAND2_X1 U743 ( .A1(n657), .A2(G86), .ZN(n660) );
  NAND2_X1 U744 ( .A1(G61), .A2(n658), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U746 ( .A(KEYINPUT91), .B(n661), .Z(n662) );
  NOR2_X1 U747 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U748 ( .A1(n664), .A2(G48), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n666), .A2(n665), .ZN(G305) );
  XOR2_X1 U750 ( .A(n676), .B(G290), .Z(n672) );
  XOR2_X1 U751 ( .A(KEYINPUT19), .B(KEYINPUT93), .Z(n668) );
  XNOR2_X1 U752 ( .A(G299), .B(G166), .ZN(n667) );
  XNOR2_X1 U753 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U754 ( .A(n669), .B(G305), .Z(n670) );
  XNOR2_X1 U755 ( .A(G288), .B(n670), .ZN(n671) );
  XNOR2_X1 U756 ( .A(n672), .B(n671), .ZN(n848) );
  XOR2_X1 U757 ( .A(n848), .B(n673), .Z(n674) );
  NOR2_X1 U758 ( .A1(n675), .A2(n674), .ZN(n678) );
  NOR2_X1 U759 ( .A1(G868), .A2(n676), .ZN(n677) );
  NOR2_X1 U760 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2078), .A2(G2084), .ZN(n680) );
  XOR2_X1 U762 ( .A(KEYINPUT20), .B(KEYINPUT94), .Z(n679) );
  XNOR2_X1 U763 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n683), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U767 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U768 ( .A1(G220), .A2(G219), .ZN(n684) );
  XNOR2_X1 U769 ( .A(KEYINPUT22), .B(n684), .ZN(n685) );
  NAND2_X1 U770 ( .A1(n685), .A2(G96), .ZN(n686) );
  NOR2_X1 U771 ( .A1(n686), .A2(G218), .ZN(n687) );
  XNOR2_X1 U772 ( .A(n687), .B(KEYINPUT95), .ZN(n846) );
  NAND2_X1 U773 ( .A1(n846), .A2(G2106), .ZN(n691) );
  NAND2_X1 U774 ( .A1(G69), .A2(G120), .ZN(n688) );
  NOR2_X1 U775 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U776 ( .A1(G108), .A2(n689), .ZN(n845) );
  NAND2_X1 U777 ( .A1(n845), .A2(G567), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n691), .A2(n690), .ZN(n923) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n923), .A2(n692), .ZN(n844) );
  NAND2_X1 U781 ( .A1(n844), .A2(G36), .ZN(G176) );
  NAND2_X1 U782 ( .A1(G138), .A2(n900), .ZN(n694) );
  NAND2_X1 U783 ( .A1(G102), .A2(n901), .ZN(n693) );
  NAND2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n698) );
  NAND2_X1 U785 ( .A1(G114), .A2(n906), .ZN(n696) );
  NAND2_X1 U786 ( .A1(G126), .A2(n904), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U788 ( .A1(n698), .A2(n697), .ZN(G164) );
  XNOR2_X1 U789 ( .A(G1986), .B(G290), .ZN(n969) );
  NOR2_X1 U790 ( .A1(G164), .A2(G1384), .ZN(n722) );
  NAND2_X1 U791 ( .A1(G160), .A2(G40), .ZN(n721) );
  NOR2_X1 U792 ( .A1(n722), .A2(n721), .ZN(n836) );
  NAND2_X1 U793 ( .A1(n969), .A2(n836), .ZN(n699) );
  XNOR2_X1 U794 ( .A(n699), .B(KEYINPUT96), .ZN(n720) );
  NAND2_X1 U795 ( .A1(G141), .A2(n900), .ZN(n701) );
  NAND2_X1 U796 ( .A1(G117), .A2(n906), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n901), .A2(G105), .ZN(n702) );
  XOR2_X1 U799 ( .A(KEYINPUT38), .B(n702), .Z(n703) );
  NOR2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n904), .A2(G129), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n889) );
  NAND2_X1 U803 ( .A1(G1996), .A2(n889), .ZN(n707) );
  XOR2_X1 U804 ( .A(KEYINPUT100), .B(n707), .Z(n717) );
  INV_X1 U805 ( .A(G1991), .ZN(n1005) );
  NAND2_X1 U806 ( .A1(G131), .A2(n900), .ZN(n709) );
  NAND2_X1 U807 ( .A1(G95), .A2(n901), .ZN(n708) );
  NAND2_X1 U808 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U809 ( .A(KEYINPUT98), .B(n710), .ZN(n714) );
  NAND2_X1 U810 ( .A1(G107), .A2(n906), .ZN(n712) );
  NAND2_X1 U811 ( .A1(G119), .A2(n904), .ZN(n711) );
  NAND2_X1 U812 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U813 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U814 ( .A(KEYINPUT99), .B(n715), .Z(n895) );
  NOR2_X1 U815 ( .A1(n1005), .A2(n895), .ZN(n716) );
  NOR2_X1 U816 ( .A1(n717), .A2(n716), .ZN(n936) );
  INV_X1 U817 ( .A(n836), .ZN(n718) );
  NOR2_X1 U818 ( .A1(n936), .A2(n718), .ZN(n828) );
  INV_X1 U819 ( .A(n828), .ZN(n719) );
  NAND2_X1 U820 ( .A1(n720), .A2(n719), .ZN(n812) );
  INV_X1 U821 ( .A(n721), .ZN(n723) );
  NAND2_X1 U822 ( .A1(n739), .A2(G2072), .ZN(n725) );
  INV_X1 U823 ( .A(KEYINPUT27), .ZN(n724) );
  XNOR2_X1 U824 ( .A(n725), .B(n724), .ZN(n728) );
  NAND2_X1 U825 ( .A1(G1956), .A2(n771), .ZN(n726) );
  XNOR2_X1 U826 ( .A(n726), .B(KEYINPUT102), .ZN(n727) );
  NAND2_X1 U827 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U828 ( .A(n729), .B(KEYINPUT103), .ZN(n748) );
  XNOR2_X1 U829 ( .A(n730), .B(KEYINPUT28), .ZN(n752) );
  AND2_X1 U830 ( .A1(n731), .A2(n954), .ZN(n737) );
  INV_X1 U831 ( .A(KEYINPUT104), .ZN(n736) );
  NAND2_X1 U832 ( .A1(G1996), .A2(n739), .ZN(n732) );
  XNOR2_X1 U833 ( .A(n732), .B(KEYINPUT26), .ZN(n734) );
  NAND2_X1 U834 ( .A1(G1341), .A2(n771), .ZN(n733) );
  NAND2_X1 U835 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U836 ( .A(n736), .B(n735), .ZN(n744) );
  NAND2_X1 U837 ( .A1(n737), .A2(n744), .ZN(n743) );
  INV_X1 U838 ( .A(G1348), .ZN(n959) );
  NOR2_X1 U839 ( .A1(n739), .A2(n959), .ZN(n738) );
  XNOR2_X1 U840 ( .A(n738), .B(KEYINPUT105), .ZN(n741) );
  NAND2_X1 U841 ( .A1(n739), .A2(G2067), .ZN(n740) );
  NAND2_X1 U842 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U843 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U844 ( .A1(n744), .A2(n954), .ZN(n745) );
  NAND2_X1 U845 ( .A1(n745), .A2(n960), .ZN(n746) );
  NAND2_X1 U846 ( .A1(n747), .A2(n746), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n748), .A2(n961), .ZN(n749) );
  NAND2_X1 U848 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n754) );
  XOR2_X1 U850 ( .A(KEYINPUT106), .B(KEYINPUT29), .Z(n753) );
  XNOR2_X1 U851 ( .A(n754), .B(n753), .ZN(n759) );
  XOR2_X1 U852 ( .A(G2078), .B(KEYINPUT25), .Z(n1009) );
  NOR2_X1 U853 ( .A1(n1009), .A2(n771), .ZN(n755) );
  XNOR2_X1 U854 ( .A(n755), .B(KEYINPUT101), .ZN(n757) );
  INV_X1 U855 ( .A(G1961), .ZN(n977) );
  NAND2_X1 U856 ( .A1(n977), .A2(n771), .ZN(n756) );
  NAND2_X1 U857 ( .A1(n757), .A2(n756), .ZN(n765) );
  NAND2_X1 U858 ( .A1(n765), .A2(G171), .ZN(n758) );
  NAND2_X1 U859 ( .A1(n759), .A2(n758), .ZN(n770) );
  NOR2_X1 U860 ( .A1(G1966), .A2(n806), .ZN(n783) );
  NOR2_X1 U861 ( .A1(G2084), .A2(n771), .ZN(n780) );
  NOR2_X1 U862 ( .A1(n783), .A2(n780), .ZN(n760) );
  NAND2_X1 U863 ( .A1(G8), .A2(n760), .ZN(n763) );
  NOR2_X1 U864 ( .A1(G168), .A2(n764), .ZN(n767) );
  NOR2_X1 U865 ( .A1(G171), .A2(n765), .ZN(n766) );
  NOR2_X1 U866 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U867 ( .A(KEYINPUT31), .B(n768), .Z(n769) );
  NAND2_X1 U868 ( .A1(n770), .A2(n769), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n781), .A2(G286), .ZN(n778) );
  INV_X1 U870 ( .A(G8), .ZN(n776) );
  NOR2_X1 U871 ( .A1(G1971), .A2(n806), .ZN(n773) );
  NOR2_X1 U872 ( .A1(G2090), .A2(n771), .ZN(n772) );
  NOR2_X1 U873 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U874 ( .A1(n774), .A2(G303), .ZN(n775) );
  OR2_X1 U875 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U876 ( .A(n779), .B(KEYINPUT32), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G8), .A2(n780), .ZN(n785) );
  INV_X1 U878 ( .A(n781), .ZN(n782) );
  NOR2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n800) );
  NOR2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n795) );
  NOR2_X1 U883 ( .A1(G1971), .A2(G303), .ZN(n788) );
  NOR2_X1 U884 ( .A1(n795), .A2(n788), .ZN(n956) );
  NAND2_X1 U885 ( .A1(n800), .A2(n956), .ZN(n791) );
  NAND2_X1 U886 ( .A1(G1976), .A2(G288), .ZN(n955) );
  INV_X1 U887 ( .A(n955), .ZN(n789) );
  NOR2_X1 U888 ( .A1(n806), .A2(n789), .ZN(n790) );
  NOR2_X1 U889 ( .A1(KEYINPUT33), .A2(n794), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n795), .A2(KEYINPUT33), .ZN(n796) );
  NOR2_X1 U891 ( .A1(n796), .A2(n806), .ZN(n797) );
  XOR2_X1 U892 ( .A(G1981), .B(G305), .Z(n950) );
  NAND2_X1 U893 ( .A1(n799), .A2(n950), .ZN(n810) );
  NOR2_X1 U894 ( .A1(G2090), .A2(G303), .ZN(n801) );
  NAND2_X1 U895 ( .A1(G8), .A2(n801), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n800), .A2(n802), .ZN(n803) );
  AND2_X1 U897 ( .A1(n803), .A2(n806), .ZN(n808) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n804) );
  XOR2_X1 U899 ( .A(n804), .B(KEYINPUT24), .Z(n805) );
  NOR2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  AND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n824) );
  XOR2_X1 U904 ( .A(G2067), .B(KEYINPUT37), .Z(n813) );
  XNOR2_X1 U905 ( .A(KEYINPUT97), .B(n813), .ZN(n834) );
  NAND2_X1 U906 ( .A1(G140), .A2(n900), .ZN(n815) );
  NAND2_X1 U907 ( .A1(G104), .A2(n901), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U909 ( .A(KEYINPUT34), .B(n816), .ZN(n821) );
  NAND2_X1 U910 ( .A1(G116), .A2(n906), .ZN(n818) );
  NAND2_X1 U911 ( .A1(G128), .A2(n904), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U913 ( .A(KEYINPUT35), .B(n819), .Z(n820) );
  NOR2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U915 ( .A(KEYINPUT36), .B(n822), .ZN(n913) );
  NOR2_X1 U916 ( .A1(n834), .A2(n913), .ZN(n930) );
  NAND2_X1 U917 ( .A1(n930), .A2(n836), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n839) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n889), .ZN(n925) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n826) );
  INV_X1 U921 ( .A(n895), .ZN(n825) );
  NOR2_X1 U922 ( .A1(G1991), .A2(n825), .ZN(n934) );
  NOR2_X1 U923 ( .A1(n826), .A2(n934), .ZN(n827) );
  NOR2_X1 U924 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n829), .B(KEYINPUT108), .ZN(n830) );
  NOR2_X1 U926 ( .A1(n925), .A2(n830), .ZN(n831) );
  XNOR2_X1 U927 ( .A(n831), .B(KEYINPUT39), .ZN(n833) );
  INV_X1 U928 ( .A(n930), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n834), .A2(n913), .ZN(n938) );
  NAND2_X1 U931 ( .A1(n835), .A2(n938), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U934 ( .A(KEYINPUT40), .B(n840), .ZN(G329) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n841), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U939 ( .A1(n844), .A2(n843), .ZN(G188) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n847), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U946 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U947 ( .A(G286), .B(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n960), .B(n954), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(G171), .B(n851), .Z(n852) );
  NOR2_X1 U951 ( .A1(G37), .A2(n852), .ZN(n853) );
  XOR2_X1 U952 ( .A(KEYINPUT117), .B(n853), .Z(G397) );
  XNOR2_X1 U953 ( .A(G1996), .B(KEYINPUT41), .ZN(n863) );
  XOR2_X1 U954 ( .A(G1981), .B(G1956), .Z(n855) );
  XNOR2_X1 U955 ( .A(G1991), .B(G1961), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U957 ( .A(G1976), .B(G1971), .Z(n857) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1966), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U961 ( .A(KEYINPUT110), .B(G2474), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G229) );
  XOR2_X1 U964 ( .A(G2100), .B(G2096), .Z(n865) );
  XNOR2_X1 U965 ( .A(KEYINPUT42), .B(G2678), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U967 ( .A(KEYINPUT43), .B(G2090), .Z(n867) );
  XNOR2_X1 U968 ( .A(G2067), .B(G2072), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U970 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U971 ( .A(G2078), .B(G2084), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(G227) );
  NAND2_X1 U973 ( .A1(G100), .A2(n901), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G112), .A2(n906), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G136), .A2(n900), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(KEYINPUT112), .ZN(n878) );
  XOR2_X1 U978 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n876) );
  NAND2_X1 U979 ( .A1(G124), .A2(n904), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U982 ( .A1(n880), .A2(n879), .ZN(G162) );
  NAND2_X1 U983 ( .A1(G142), .A2(n900), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G106), .A2(n901), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U986 ( .A(n883), .B(KEYINPUT45), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G118), .A2(n906), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G130), .A2(n904), .ZN(n886) );
  XNOR2_X1 U990 ( .A(KEYINPUT113), .B(n886), .ZN(n887) );
  NOR2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n899) );
  XNOR2_X1 U992 ( .A(G162), .B(n889), .ZN(n890) );
  XNOR2_X1 U993 ( .A(n890), .B(n927), .ZN(n894) );
  XOR2_X1 U994 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n892) );
  XNOR2_X1 U995 ( .A(G164), .B(KEYINPUT46), .ZN(n891) );
  XNOR2_X1 U996 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U997 ( .A(n894), .B(n893), .Z(n897) );
  XNOR2_X1 U998 ( .A(G160), .B(n895), .ZN(n896) );
  XNOR2_X1 U999 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n915) );
  NAND2_X1 U1001 ( .A1(G139), .A2(n900), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(G103), .A2(n901), .ZN(n902) );
  NAND2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n912) );
  NAND2_X1 U1004 ( .A1(n904), .A2(G127), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n905), .B(KEYINPUT114), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(G115), .A2(n906), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT115), .B(n909), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(KEYINPUT47), .B(n910), .ZN(n911) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n940) );
  XNOR2_X1 U1011 ( .A(n913), .B(n940), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n916), .ZN(G395) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(G397), .A2(n918), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(n923), .A2(G401), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT118), .B(n919), .Z(n920) );
  NOR2_X1 U1019 ( .A1(G395), .A2(n920), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(n923), .ZN(G319) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n926), .Z(n932) );
  XNOR2_X1 U1027 ( .A(G160), .B(G2084), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n937), .B(KEYINPUT119), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1035 ( .A(G2072), .B(n940), .Z(n942) );
  XOR2_X1 U1036 ( .A(G164), .B(G2078), .Z(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1038 ( .A(KEYINPUT50), .B(n943), .Z(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n946), .ZN(n948) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n949), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1044 ( .A(KEYINPUT56), .B(G16), .ZN(n976) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G168), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n952), .B(KEYINPUT57), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT122), .B(n953), .ZN(n974) );
  XOR2_X1 U1049 ( .A(n954), .B(G1341), .Z(n972) );
  AND2_X1 U1050 ( .A1(G303), .A2(G1971), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n967) );
  XNOR2_X1 U1053 ( .A(n960), .B(n959), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(n961), .B(G1956), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(G1961), .B(G301), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(KEYINPUT123), .B(n970), .ZN(n971) );
  NOR2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1062 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1063 ( .A1(n976), .A2(n975), .ZN(n1004) );
  XOR2_X1 U1064 ( .A(KEYINPUT124), .B(G16), .Z(n1002) );
  XNOR2_X1 U1065 ( .A(G5), .B(n977), .ZN(n991) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G21), .ZN(n989) );
  XNOR2_X1 U1067 ( .A(KEYINPUT59), .B(G4), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n978), .B(KEYINPUT125), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n979), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n985) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G20), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(G1981), .B(G6), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n986), .B(KEYINPUT60), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(KEYINPUT126), .B(n987), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n998) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G23), .B(G1976), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n995) );
  XOR2_X1 U1083 ( .A(G1986), .B(G24), .Z(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(KEYINPUT58), .B(n996), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n999) );
  XNOR2_X1 U1088 ( .A(n1000), .B(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1028) );
  XOR2_X1 U1091 ( .A(G29), .B(KEYINPUT120), .Z(n1024) );
  XNOR2_X1 U1092 ( .A(G25), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(G28), .ZN(n1015) );
  XNOR2_X1 U1094 ( .A(G2067), .B(G26), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G33), .B(G2072), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G1996), .B(G32), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G27), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(KEYINPUT53), .B(n1016), .Z(n1019) );
  XOR2_X1 U1103 ( .A(KEYINPUT54), .B(G34), .Z(n1017) );
  XNOR2_X1 U1104 ( .A(G2084), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(G35), .B(G2090), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(n1022), .B(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(G11), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(KEYINPUT121), .B(n1026), .Z(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

