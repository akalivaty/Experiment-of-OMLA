

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767;

  NAND2_X1 U371 ( .A1(n364), .A2(n571), .ZN(n614) );
  NAND2_X1 U372 ( .A1(n557), .A2(n558), .ZN(n737) );
  AND2_X2 U373 ( .A1(n381), .A2(n409), .ZN(n355) );
  AND2_X2 U374 ( .A1(n643), .A2(n642), .ZN(n647) );
  NOR2_X2 U375 ( .A1(n607), .A2(n408), .ZN(n396) );
  OR2_X2 U376 ( .A1(n657), .A2(n411), .ZN(n381) );
  XNOR2_X2 U377 ( .A(n747), .B(n527), .ZN(n657) );
  NOR2_X1 U378 ( .A1(n766), .A2(n767), .ZN(n366) );
  XNOR2_X1 U379 ( .A(n414), .B(KEYINPUT85), .ZN(n624) );
  NOR2_X1 U380 ( .A1(n579), .A2(n695), .ZN(n580) );
  AND2_X1 U381 ( .A1(n378), .A2(n371), .ZN(n370) );
  NOR2_X1 U382 ( .A1(n723), .A2(n585), .ZN(n586) );
  NOR2_X1 U383 ( .A1(n362), .A2(n620), .ZN(n739) );
  AND2_X1 U384 ( .A1(n545), .A2(n360), .ZN(n551) );
  XNOR2_X1 U385 ( .A(n584), .B(n583), .ZN(n723) );
  XNOR2_X1 U386 ( .A(n624), .B(KEYINPUT19), .ZN(n620) );
  OR2_X1 U387 ( .A1(n695), .A2(n579), .ZN(n562) );
  XNOR2_X1 U388 ( .A(n618), .B(KEYINPUT1), .ZN(n579) );
  XNOR2_X1 U389 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U390 ( .A1(n410), .A2(n535), .ZN(n409) );
  XNOR2_X1 U391 ( .A(n752), .B(G146), .ZN(n464) );
  XNOR2_X1 U392 ( .A(n506), .B(n421), .ZN(n754) );
  XNOR2_X1 U393 ( .A(n452), .B(n451), .ZN(n517) );
  XNOR2_X1 U394 ( .A(n492), .B(n491), .ZN(n505) );
  XNOR2_X1 U395 ( .A(n450), .B(KEYINPUT3), .ZN(n452) );
  XNOR2_X1 U396 ( .A(G113), .B(KEYINPUT67), .ZN(n451) );
  XOR2_X1 U397 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n492) );
  BUF_X1 U398 ( .A(n673), .Z(n680) );
  INV_X1 U399 ( .A(n479), .ZN(n421) );
  XNOR2_X1 U400 ( .A(n629), .B(n401), .ZN(n634) );
  INV_X1 U401 ( .A(KEYINPUT38), .ZN(n401) );
  XNOR2_X1 U402 ( .A(n455), .B(G472), .ZN(n699) );
  XNOR2_X1 U403 ( .A(n513), .B(n352), .ZN(n693) );
  NOR2_X1 U404 ( .A1(n372), .A2(n375), .ZN(n371) );
  INV_X1 U405 ( .A(n628), .ZN(n372) );
  AND2_X1 U406 ( .A1(n365), .A2(n353), .ZN(n641) );
  XNOR2_X1 U407 ( .A(n366), .B(KEYINPUT46), .ZN(n365) );
  AND2_X1 U408 ( .A1(n376), .A2(n375), .ZN(n374) );
  NOR2_X1 U409 ( .A1(n641), .A2(KEYINPUT48), .ZN(n377) );
  OR2_X1 U410 ( .A1(n596), .A2(n595), .ZN(n609) );
  NOR2_X1 U411 ( .A1(n408), .A2(n608), .ZN(n405) );
  XNOR2_X1 U412 ( .A(n524), .B(n388), .ZN(n387) );
  INV_X1 U413 ( .A(G137), .ZN(n388) );
  XNOR2_X1 U414 ( .A(n573), .B(KEYINPUT105), .ZN(n626) );
  NAND2_X1 U415 ( .A1(n626), .A2(n439), .ZN(n438) );
  AND2_X1 U416 ( .A1(n625), .A2(n627), .ZN(n439) );
  NOR2_X1 U417 ( .A1(n696), .A2(n437), .ZN(n436) );
  NOR2_X1 U418 ( .A1(n625), .A2(n627), .ZN(n437) );
  INV_X1 U419 ( .A(KEYINPUT110), .ZN(n431) );
  NAND2_X1 U420 ( .A1(n532), .A2(n528), .ZN(n412) );
  OR2_X1 U421 ( .A1(n532), .A2(n528), .ZN(n411) );
  XNOR2_X1 U422 ( .A(n399), .B(n398), .ZN(n722) );
  INV_X1 U423 ( .A(KEYINPUT41), .ZN(n398) );
  NAND2_X1 U424 ( .A1(n711), .A2(n400), .ZN(n399) );
  NOR2_X1 U425 ( .A1(n713), .A2(n535), .ZN(n400) );
  AND2_X1 U426 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X1 U427 ( .A1(n619), .A2(n618), .ZN(n362) );
  XNOR2_X1 U428 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n616) );
  BUF_X1 U429 ( .A(n579), .Z(n696) );
  XNOR2_X1 U430 ( .A(n391), .B(n546), .ZN(n567) );
  NAND2_X1 U431 ( .A1(n545), .A2(n544), .ZN(n391) );
  XNOR2_X1 U432 ( .A(n508), .B(n509), .ZN(n674) );
  XNOR2_X1 U433 ( .A(n504), .B(n367), .ZN(n509) );
  XNOR2_X1 U434 ( .A(n425), .B(n656), .ZN(n424) );
  NAND2_X1 U435 ( .A1(n673), .A2(G475), .ZN(n425) );
  NOR2_X1 U436 ( .A1(n756), .A2(G952), .ZN(n686) );
  INV_X1 U437 ( .A(KEYINPUT48), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n764), .B(KEYINPUT80), .ZN(n378) );
  INV_X1 U439 ( .A(G237), .ZN(n456) );
  INV_X1 U440 ( .A(n412), .ZN(n410) );
  XNOR2_X1 U441 ( .A(G131), .B(G101), .ZN(n447) );
  XOR2_X1 U442 ( .A(KEYINPUT5), .B(KEYINPUT70), .Z(n448) );
  NOR2_X1 U443 ( .A1(n377), .A2(n374), .ZN(n373) );
  NAND2_X1 U444 ( .A1(n641), .A2(n370), .ZN(n369) );
  XNOR2_X1 U445 ( .A(G113), .B(G143), .ZN(n483) );
  NAND2_X1 U446 ( .A1(G234), .A2(G237), .ZN(n469) );
  XNOR2_X1 U447 ( .A(n444), .B(n442), .ZN(n552) );
  XNOR2_X1 U448 ( .A(n488), .B(n443), .ZN(n442) );
  OR2_X1 U449 ( .A1(n655), .A2(G902), .ZN(n444) );
  INV_X1 U450 ( .A(G475), .ZN(n443) );
  NAND2_X1 U451 ( .A1(n406), .A2(n612), .ZN(n384) );
  XNOR2_X1 U452 ( .A(G119), .B(G110), .ZN(n502) );
  INV_X1 U453 ( .A(KEYINPUT10), .ZN(n478) );
  XNOR2_X1 U454 ( .A(n503), .B(n368), .ZN(n367) );
  XNOR2_X1 U455 ( .A(G128), .B(G137), .ZN(n503) );
  XNOR2_X1 U456 ( .A(KEYINPUT23), .B(G140), .ZN(n368) );
  INV_X1 U457 ( .A(G134), .ZN(n446) );
  XNOR2_X1 U458 ( .A(G116), .B(G107), .ZN(n489) );
  INV_X1 U459 ( .A(n755), .ZN(n380) );
  NOR2_X1 U460 ( .A1(n627), .A2(n431), .ZN(n430) );
  AND2_X1 U461 ( .A1(n357), .A2(n438), .ZN(n379) );
  NOR2_X1 U462 ( .A1(n696), .A2(n693), .ZN(n568) );
  NAND2_X1 U463 ( .A1(n356), .A2(n413), .ZN(n629) );
  AND2_X1 U464 ( .A1(n393), .A2(n477), .ZN(n631) );
  INV_X1 U465 ( .A(n693), .ZN(n364) );
  XNOR2_X1 U466 ( .A(n552), .B(n441), .ZN(n557) );
  INV_X1 U467 ( .A(KEYINPUT98), .ZN(n441) );
  XOR2_X1 U468 ( .A(KEYINPUT62), .B(n666), .Z(n667) );
  NOR2_X1 U469 ( .A1(n722), .A2(n362), .ZN(n635) );
  NAND2_X1 U470 ( .A1(n428), .A2(n427), .ZN(n764) );
  NAND2_X1 U471 ( .A1(n426), .A2(n379), .ZN(n427) );
  AND2_X1 U472 ( .A1(n432), .A2(n429), .ZN(n428) );
  NAND2_X1 U473 ( .A1(n434), .A2(n433), .ZN(n426) );
  INV_X1 U474 ( .A(G122), .ZN(n591) );
  XNOR2_X1 U475 ( .A(n354), .B(n563), .ZN(n597) );
  XNOR2_X1 U476 ( .A(n551), .B(n550), .ZN(n598) );
  XNOR2_X1 U477 ( .A(n594), .B(KEYINPUT103), .ZN(n408) );
  XNOR2_X1 U478 ( .A(n395), .B(n394), .ZN(n675) );
  INV_X1 U479 ( .A(n674), .ZN(n394) );
  NAND2_X1 U480 ( .A1(n680), .A2(G217), .ZN(n395) );
  INV_X1 U481 ( .A(KEYINPUT60), .ZN(n422) );
  INV_X1 U482 ( .A(n686), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n408), .B(n382), .ZN(G3) );
  INV_X1 U484 ( .A(G101), .ZN(n382) );
  XOR2_X1 U485 ( .A(KEYINPUT72), .B(n646), .Z(n350) );
  AND2_X1 U486 ( .A1(n350), .A2(KEYINPUT78), .ZN(n351) );
  XOR2_X1 U487 ( .A(n512), .B(KEYINPUT25), .Z(n352) );
  XOR2_X1 U488 ( .A(KEYINPUT74), .B(n640), .Z(n353) );
  AND2_X1 U489 ( .A1(n385), .A2(n545), .ZN(n354) );
  NAND2_X1 U490 ( .A1(n386), .A2(n649), .ZN(n650) );
  AND2_X1 U491 ( .A1(n381), .A2(n412), .ZN(n356) );
  AND2_X1 U492 ( .A1(n436), .A2(n431), .ZN(n357) );
  AND2_X1 U493 ( .A1(n566), .A2(n696), .ZN(n358) );
  AND2_X1 U494 ( .A1(n383), .A2(n380), .ZN(n359) );
  AND2_X1 U495 ( .A1(n615), .A2(n549), .ZN(n360) );
  AND2_X1 U496 ( .A1(n568), .A2(n566), .ZN(n361) );
  XNOR2_X1 U497 ( .A(KEYINPUT15), .B(G902), .ZN(n651) );
  INV_X1 U498 ( .A(KEYINPUT78), .ZN(n440) );
  NAND2_X1 U499 ( .A1(n693), .A2(n363), .ZN(n695) );
  INV_X1 U500 ( .A(n692), .ZN(n363) );
  NOR2_X1 U501 ( .A1(n634), .A2(n364), .ZN(n630) );
  OR2_X1 U502 ( .A1(n587), .A2(n364), .ZN(n533) );
  AND2_X1 U503 ( .A1(n696), .A2(n364), .ZN(n547) );
  NAND2_X1 U504 ( .A1(n373), .A2(n369), .ZN(n643) );
  NAND2_X1 U505 ( .A1(n378), .A2(n628), .ZN(n376) );
  NAND2_X1 U506 ( .A1(n380), .A2(n528), .ZN(n419) );
  XNOR2_X2 U507 ( .A(n523), .B(n446), .ZN(n497) );
  XNOR2_X2 U508 ( .A(G143), .B(G128), .ZN(n523) );
  NAND2_X1 U509 ( .A1(n397), .A2(n653), .ZN(n416) );
  OR2_X2 U510 ( .A1(n383), .A2(n741), .ZN(n397) );
  XNOR2_X2 U511 ( .A(n384), .B(n613), .ZN(n741) );
  INV_X1 U512 ( .A(n650), .ZN(n383) );
  INV_X1 U513 ( .A(n545), .ZN(n585) );
  XNOR2_X2 U514 ( .A(n542), .B(KEYINPUT0), .ZN(n545) );
  INV_X1 U515 ( .A(n704), .ZN(n385) );
  NOR2_X1 U516 ( .A1(n662), .A2(n686), .ZN(n665) );
  NOR2_X1 U517 ( .A1(n669), .A2(n686), .ZN(n672) );
  NAND2_X1 U518 ( .A1(n567), .A2(n358), .ZN(n592) );
  NAND2_X1 U519 ( .A1(n392), .A2(n603), .ZN(n607) );
  NAND2_X1 U520 ( .A1(n648), .A2(n440), .ZN(n386) );
  XNOR2_X2 U521 ( .A(n497), .B(n387), .ZN(n752) );
  INV_X1 U522 ( .A(n699), .ZN(n615) );
  NAND2_X1 U523 ( .A1(n699), .A2(n710), .ZN(n457) );
  NAND2_X1 U524 ( .A1(n420), .A2(n359), .ZN(n688) );
  XNOR2_X1 U525 ( .A(n389), .B(n422), .ZN(G60) );
  NAND2_X1 U526 ( .A1(n424), .A2(n423), .ZN(n389) );
  NAND2_X1 U527 ( .A1(n597), .A2(n598), .ZN(n599) );
  NAND2_X1 U528 ( .A1(n390), .A2(n608), .ZN(n404) );
  NAND2_X1 U529 ( .A1(n396), .A2(n407), .ZN(n390) );
  XNOR2_X1 U530 ( .A(n602), .B(n601), .ZN(n392) );
  XNOR2_X1 U531 ( .A(n457), .B(n458), .ZN(n393) );
  NOR2_X1 U532 ( .A1(n650), .A2(n419), .ZN(n418) );
  NAND2_X1 U533 ( .A1(n355), .A2(n413), .ZN(n414) );
  NAND2_X1 U534 ( .A1(n397), .A2(n689), .ZN(n690) );
  NAND2_X1 U535 ( .A1(n711), .A2(n710), .ZN(n707) );
  NAND2_X1 U536 ( .A1(n404), .A2(n402), .ZN(n406) );
  NAND2_X1 U537 ( .A1(n405), .A2(n403), .ZN(n402) );
  NOR2_X1 U538 ( .A1(n607), .A2(n606), .ZN(n403) );
  INV_X1 U539 ( .A(n606), .ZN(n407) );
  NAND2_X1 U540 ( .A1(n657), .A2(n532), .ZN(n413) );
  XNOR2_X1 U541 ( .A(n415), .B(n478), .ZN(n506) );
  XNOR2_X1 U542 ( .A(n519), .B(n415), .ZN(n522) );
  XNOR2_X2 U543 ( .A(G146), .B(G125), .ZN(n415) );
  NAND2_X2 U544 ( .A1(n416), .A2(n417), .ZN(n673) );
  NAND2_X1 U545 ( .A1(n418), .A2(n420), .ZN(n417) );
  INV_X1 U546 ( .A(n741), .ZN(n420) );
  NAND2_X1 U547 ( .A1(n567), .A2(n361), .ZN(n570) );
  NAND2_X1 U548 ( .A1(n438), .A2(n436), .ZN(n435) );
  NAND2_X1 U549 ( .A1(n434), .A2(n430), .ZN(n429) );
  NAND2_X1 U550 ( .A1(n435), .A2(KEYINPUT110), .ZN(n432) );
  INV_X1 U551 ( .A(n627), .ZN(n433) );
  INV_X1 U552 ( .A(n626), .ZN(n434) );
  NAND2_X1 U553 ( .A1(n647), .A2(n351), .ZN(n649) );
  NAND2_X1 U554 ( .A1(n647), .A2(n350), .ZN(n648) );
  AND2_X1 U555 ( .A1(n480), .A2(G210), .ZN(n445) );
  INV_X1 U556 ( .A(KEYINPUT101), .ZN(n601) );
  XNOR2_X1 U557 ( .A(n449), .B(n445), .ZN(n453) );
  INV_X1 U558 ( .A(KEYINPUT82), .ZN(n608) );
  XNOR2_X1 U559 ( .A(n516), .B(n461), .ZN(n462) );
  XNOR2_X1 U560 ( .A(n453), .B(n517), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n462), .B(n479), .ZN(n463) );
  OR2_X1 U562 ( .A1(n615), .A2(n562), .ZN(n704) );
  XNOR2_X1 U563 ( .A(n464), .B(n454), .ZN(n666) );
  XNOR2_X1 U564 ( .A(n464), .B(n463), .ZN(n681) );
  INV_X1 U565 ( .A(KEYINPUT94), .ZN(n550) );
  XOR2_X1 U566 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n458) );
  XNOR2_X2 U567 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n524) );
  XNOR2_X1 U568 ( .A(n448), .B(n447), .ZN(n449) );
  NOR2_X1 U569 ( .A1(G953), .A2(G237), .ZN(n480) );
  XNOR2_X2 U570 ( .A(G119), .B(G116), .ZN(n450) );
  INV_X1 U571 ( .A(G902), .ZN(n510) );
  NAND2_X1 U572 ( .A1(n666), .A2(n510), .ZN(n455) );
  NAND2_X1 U573 ( .A1(n510), .A2(n456), .ZN(n529) );
  NAND2_X1 U574 ( .A1(n529), .A2(G214), .ZN(n710) );
  XNOR2_X2 U575 ( .A(G104), .B(G101), .ZN(n460) );
  XNOR2_X2 U576 ( .A(G110), .B(G107), .ZN(n459) );
  XNOR2_X2 U577 ( .A(n460), .B(n459), .ZN(n516) );
  INV_X2 U578 ( .A(G953), .ZN(n756) );
  NAND2_X1 U579 ( .A1(G227), .A2(n756), .ZN(n461) );
  XOR2_X1 U580 ( .A(G131), .B(G140), .Z(n479) );
  NOR2_X1 U581 ( .A1(n681), .A2(G902), .ZN(n465) );
  XNOR2_X2 U582 ( .A(n465), .B(G469), .ZN(n618) );
  XOR2_X1 U583 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n467) );
  NAND2_X1 U584 ( .A1(G234), .A2(n651), .ZN(n466) );
  XNOR2_X1 U585 ( .A(n467), .B(n466), .ZN(n511) );
  NAND2_X1 U586 ( .A1(n511), .A2(G221), .ZN(n468) );
  XNOR2_X1 U587 ( .A(KEYINPUT21), .B(n468), .ZN(n692) );
  XNOR2_X1 U588 ( .A(n469), .B(KEYINPUT90), .ZN(n470) );
  XNOR2_X1 U589 ( .A(KEYINPUT14), .B(n470), .ZN(n472) );
  NAND2_X1 U590 ( .A1(n472), .A2(G952), .ZN(n471) );
  XOR2_X1 U591 ( .A(KEYINPUT91), .B(n471), .Z(n721) );
  NOR2_X1 U592 ( .A1(G953), .A2(n721), .ZN(n538) );
  AND2_X1 U593 ( .A1(n472), .A2(G953), .ZN(n473) );
  NAND2_X1 U594 ( .A1(G902), .A2(n473), .ZN(n536) );
  NOR2_X1 U595 ( .A1(n536), .A2(G900), .ZN(n474) );
  NOR2_X1 U596 ( .A1(n538), .A2(n474), .ZN(n475) );
  NOR2_X1 U597 ( .A1(n692), .A2(n475), .ZN(n571) );
  INV_X1 U598 ( .A(n571), .ZN(n476) );
  NOR2_X1 U599 ( .A1(n618), .A2(n476), .ZN(n477) );
  XOR2_X1 U600 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n482) );
  NAND2_X1 U601 ( .A1(G214), .A2(n480), .ZN(n481) );
  XNOR2_X1 U602 ( .A(n482), .B(n481), .ZN(n486) );
  XOR2_X1 U603 ( .A(G122), .B(G104), .Z(n484) );
  XNOR2_X1 U604 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U605 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U606 ( .A(n754), .B(n487), .ZN(n655) );
  XNOR2_X1 U607 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n488) );
  INV_X1 U608 ( .A(n552), .ZN(n501) );
  XOR2_X1 U609 ( .A(KEYINPUT9), .B(G122), .Z(n490) );
  XNOR2_X1 U610 ( .A(n490), .B(n489), .ZN(n496) );
  XOR2_X1 U611 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n494) );
  NAND2_X1 U612 ( .A1(G234), .A2(n756), .ZN(n491) );
  NAND2_X1 U613 ( .A1(G217), .A2(n505), .ZN(n493) );
  XNOR2_X1 U614 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U615 ( .A(n496), .B(n495), .ZN(n498) );
  XNOR2_X1 U616 ( .A(n498), .B(n497), .ZN(n676) );
  NOR2_X1 U617 ( .A1(n676), .A2(G902), .ZN(n499) );
  XNOR2_X1 U618 ( .A(n499), .B(G478), .ZN(n558) );
  INV_X1 U619 ( .A(n558), .ZN(n500) );
  NAND2_X1 U620 ( .A1(n501), .A2(n500), .ZN(n587) );
  XNOR2_X1 U621 ( .A(n502), .B(KEYINPUT24), .ZN(n504) );
  NAND2_X1 U622 ( .A1(n505), .A2(G221), .ZN(n507) );
  XNOR2_X1 U623 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U624 ( .A1(n674), .A2(n510), .ZN(n513) );
  NAND2_X1 U625 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U626 ( .A(KEYINPUT68), .B(KEYINPUT16), .ZN(n514) );
  XNOR2_X1 U627 ( .A(n514), .B(n591), .ZN(n515) );
  XNOR2_X1 U628 ( .A(n516), .B(n515), .ZN(n518) );
  XNOR2_X1 U629 ( .A(n518), .B(n517), .ZN(n747) );
  XNOR2_X1 U630 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n519) );
  NAND2_X1 U631 ( .A1(n756), .A2(G224), .ZN(n520) );
  XNOR2_X1 U632 ( .A(n520), .B(KEYINPUT88), .ZN(n521) );
  XNOR2_X1 U633 ( .A(n522), .B(n521), .ZN(n526) );
  XNOR2_X1 U634 ( .A(n523), .B(n524), .ZN(n525) );
  XNOR2_X1 U635 ( .A(n526), .B(n525), .ZN(n527) );
  INV_X1 U636 ( .A(n651), .ZN(n528) );
  NAND2_X1 U637 ( .A1(n529), .A2(G210), .ZN(n531) );
  INV_X1 U638 ( .A(KEYINPUT89), .ZN(n530) );
  XNOR2_X1 U639 ( .A(n531), .B(n530), .ZN(n532) );
  NOR2_X1 U640 ( .A1(n533), .A2(n629), .ZN(n534) );
  NAND2_X1 U641 ( .A1(n631), .A2(n534), .ZN(n638) );
  XNOR2_X1 U642 ( .A(n638), .B(G143), .ZN(G45) );
  INV_X1 U643 ( .A(n710), .ZN(n535) );
  NOR2_X1 U644 ( .A1(G898), .A2(n536), .ZN(n537) );
  OR2_X1 U645 ( .A1(n538), .A2(n537), .ZN(n540) );
  INV_X1 U646 ( .A(KEYINPUT92), .ZN(n539) );
  NOR2_X2 U647 ( .A1(n620), .A2(n541), .ZN(n542) );
  NAND2_X1 U648 ( .A1(n552), .A2(n558), .ZN(n713) );
  NOR2_X1 U649 ( .A1(n692), .A2(n713), .ZN(n543) );
  XNOR2_X1 U650 ( .A(n543), .B(KEYINPUT102), .ZN(n544) );
  XNOR2_X1 U651 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n546) );
  AND2_X1 U652 ( .A1(n615), .A2(n547), .ZN(n548) );
  AND2_X1 U653 ( .A1(n567), .A2(n548), .ZN(n595) );
  XOR2_X1 U654 ( .A(G110), .B(n595), .Z(G12) );
  NOR2_X1 U655 ( .A1(n695), .A2(n618), .ZN(n549) );
  NOR2_X1 U656 ( .A1(n598), .A2(n737), .ZN(n554) );
  XNOR2_X1 U657 ( .A(G104), .B(KEYINPUT113), .ZN(n553) );
  XNOR2_X1 U658 ( .A(n554), .B(n553), .ZN(G6) );
  XOR2_X1 U659 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n556) );
  XNOR2_X1 U660 ( .A(G107), .B(KEYINPUT26), .ZN(n555) );
  XNOR2_X1 U661 ( .A(n556), .B(n555), .ZN(n561) );
  OR2_X1 U662 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U663 ( .A(KEYINPUT100), .B(n559), .ZN(n732) );
  NOR2_X1 U664 ( .A1(n598), .A2(n732), .ZN(n560) );
  XOR2_X1 U665 ( .A(n561), .B(n560), .Z(G9) );
  XOR2_X1 U666 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n563) );
  NOR2_X1 U667 ( .A1(n597), .A2(n737), .ZN(n564) );
  XOR2_X1 U668 ( .A(G113), .B(n564), .Z(G15) );
  NOR2_X1 U669 ( .A1(n597), .A2(n732), .ZN(n565) );
  XOR2_X1 U670 ( .A(G116), .B(n565), .Z(G18) );
  XNOR2_X1 U671 ( .A(n615), .B(KEYINPUT6), .ZN(n581) );
  INV_X1 U672 ( .A(n581), .ZN(n566) );
  INV_X1 U673 ( .A(KEYINPUT32), .ZN(n569) );
  XNOR2_X1 U674 ( .A(n570), .B(n569), .ZN(n596) );
  XOR2_X1 U675 ( .A(n596), .B(G119), .Z(G21) );
  XOR2_X1 U676 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n576) );
  NOR2_X1 U677 ( .A1(n737), .A2(n614), .ZN(n572) );
  NAND2_X1 U678 ( .A1(n572), .A2(n581), .ZN(n573) );
  AND2_X1 U679 ( .A1(n696), .A2(n626), .ZN(n574) );
  NAND2_X1 U680 ( .A1(n574), .A2(n710), .ZN(n575) );
  XNOR2_X1 U681 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U682 ( .A(n577), .B(KEYINPUT43), .ZN(n578) );
  NAND2_X1 U683 ( .A1(n578), .A2(n629), .ZN(n642) );
  XNOR2_X1 U684 ( .A(n642), .B(G140), .ZN(G42) );
  XNOR2_X1 U685 ( .A(n580), .B(KEYINPUT104), .ZN(n582) );
  NAND2_X1 U686 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U687 ( .A(KEYINPUT87), .B(KEYINPUT33), .ZN(n583) );
  XNOR2_X1 U688 ( .A(n586), .B(KEYINPUT34), .ZN(n589) );
  XNOR2_X1 U689 ( .A(n587), .B(KEYINPUT71), .ZN(n588) );
  NAND2_X1 U690 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X2 U691 ( .A(n590), .B(KEYINPUT35), .ZN(n604) );
  XNOR2_X1 U692 ( .A(n604), .B(n591), .ZN(G24) );
  XNOR2_X1 U693 ( .A(n592), .B(KEYINPUT81), .ZN(n593) );
  NAND2_X1 U694 ( .A1(n593), .A2(n693), .ZN(n594) );
  NAND2_X1 U695 ( .A1(n609), .A2(KEYINPUT44), .ZN(n603) );
  XNOR2_X1 U696 ( .A(n599), .B(KEYINPUT96), .ZN(n600) );
  NAND2_X1 U697 ( .A1(n737), .A2(n732), .ZN(n636) );
  NAND2_X1 U698 ( .A1(n600), .A2(n636), .ZN(n602) );
  NAND2_X1 U699 ( .A1(n604), .A2(KEYINPUT44), .ZN(n605) );
  XNOR2_X1 U700 ( .A(n605), .B(KEYINPUT83), .ZN(n606) );
  NOR2_X1 U701 ( .A1(n604), .A2(KEYINPUT44), .ZN(n611) );
  INV_X1 U702 ( .A(n609), .ZN(n610) );
  NAND2_X1 U703 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U704 ( .A(KEYINPUT77), .B(KEYINPUT45), .ZN(n613) );
  NOR2_X1 U705 ( .A1(n615), .A2(n614), .ZN(n617) );
  XNOR2_X1 U706 ( .A(n617), .B(n616), .ZN(n619) );
  INV_X1 U707 ( .A(n739), .ZN(n623) );
  INV_X1 U708 ( .A(n636), .ZN(n708) );
  NOR2_X1 U709 ( .A1(n708), .A2(KEYINPUT47), .ZN(n621) );
  XNOR2_X1 U710 ( .A(n621), .B(KEYINPUT69), .ZN(n622) );
  OR2_X1 U711 ( .A1(n623), .A2(n622), .ZN(n628) );
  BUF_X1 U712 ( .A(n624), .Z(n625) );
  XOR2_X1 U713 ( .A(KEYINPUT36), .B(KEYINPUT84), .Z(n627) );
  XNOR2_X1 U714 ( .A(n632), .B(KEYINPUT39), .ZN(n644) );
  NOR2_X1 U715 ( .A1(n644), .A2(n737), .ZN(n633) );
  XNOR2_X1 U716 ( .A(n633), .B(KEYINPUT40), .ZN(n767) );
  INV_X1 U717 ( .A(n634), .ZN(n711) );
  XNOR2_X1 U718 ( .A(KEYINPUT42), .B(n635), .ZN(n766) );
  NAND2_X1 U719 ( .A1(n739), .A2(n636), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n637), .A2(KEYINPUT47), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U722 ( .A1(n644), .A2(n732), .ZN(n645) );
  XNOR2_X1 U723 ( .A(n645), .B(KEYINPUT111), .ZN(n763) );
  NAND2_X1 U724 ( .A1(n647), .A2(n763), .ZN(n755) );
  NAND2_X1 U725 ( .A1(KEYINPUT2), .A2(n763), .ZN(n646) );
  XOR2_X1 U726 ( .A(KEYINPUT76), .B(n651), .Z(n652) );
  AND2_X1 U727 ( .A1(n652), .A2(KEYINPUT2), .ZN(n653) );
  XNOR2_X1 U728 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n654) );
  XOR2_X1 U729 ( .A(n655), .B(n654), .Z(n656) );
  NAND2_X1 U730 ( .A1(n673), .A2(G210), .ZN(n661) );
  XNOR2_X1 U731 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n658) );
  XOR2_X1 U732 ( .A(n658), .B(KEYINPUT55), .Z(n659) );
  XNOR2_X1 U733 ( .A(n657), .B(n659), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U735 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n663), .B(KEYINPUT79), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(G51) );
  NAND2_X1 U738 ( .A1(n673), .A2(G472), .ZN(n668) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U740 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n670) );
  XOR2_X1 U741 ( .A(n670), .B(KEYINPUT86), .Z(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G57) );
  NOR2_X1 U743 ( .A1(n675), .A2(n686), .ZN(G66) );
  NAND2_X1 U744 ( .A1(n680), .A2(G478), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n676), .B(KEYINPUT124), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n679), .A2(n686), .ZN(G63) );
  NAND2_X1 U748 ( .A1(n680), .A2(G469), .ZN(n685) );
  XOR2_X1 U749 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n682) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT58), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n681), .B(n683), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n685), .B(n684), .ZN(n687) );
  NOR2_X1 U753 ( .A1(n687), .A2(n686), .ZN(G54) );
  XOR2_X1 U754 ( .A(KEYINPUT2), .B(KEYINPUT73), .Z(n689) );
  NAND2_X1 U755 ( .A1(n688), .A2(n690), .ZN(n691) );
  XNOR2_X1 U756 ( .A(n691), .B(KEYINPUT75), .ZN(n730) );
  NOR2_X1 U757 ( .A1(n693), .A2(n363), .ZN(n694) );
  XNOR2_X1 U758 ( .A(KEYINPUT49), .B(n694), .ZN(n702) );
  XOR2_X1 U759 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n698) );
  NAND2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U761 ( .A(n698), .B(n697), .ZN(n700) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U765 ( .A(KEYINPUT51), .B(n705), .ZN(n706) );
  NOR2_X1 U766 ( .A1(n722), .A2(n706), .ZN(n718) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U768 ( .A(KEYINPUT117), .B(n709), .Z(n715) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U770 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U771 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U772 ( .A1(n723), .A2(n716), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n719), .B(KEYINPUT52), .ZN(n720) );
  NOR2_X1 U775 ( .A1(n721), .A2(n720), .ZN(n726) );
  NOR2_X1 U776 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U777 ( .A(n724), .B(KEYINPUT118), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n727), .B(KEYINPUT119), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U782 ( .A(KEYINPUT53), .B(n731), .Z(G75) );
  XOR2_X1 U783 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n735) );
  INV_X1 U784 ( .A(n732), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n739), .A2(n733), .ZN(n734) );
  XNOR2_X1 U786 ( .A(n735), .B(n734), .ZN(n736) );
  XOR2_X1 U787 ( .A(G128), .B(n736), .Z(G30) );
  INV_X1 U788 ( .A(n737), .ZN(n738) );
  NAND2_X1 U789 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U790 ( .A(n740), .B(G146), .ZN(G48) );
  NOR2_X1 U791 ( .A1(n741), .A2(G953), .ZN(n746) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n742) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n742), .ZN(n743) );
  NAND2_X1 U794 ( .A1(n743), .A2(G898), .ZN(n744) );
  XNOR2_X1 U795 ( .A(n744), .B(KEYINPUT125), .ZN(n745) );
  NOR2_X1 U796 ( .A1(n746), .A2(n745), .ZN(n751) );
  NOR2_X1 U797 ( .A1(G898), .A2(n756), .ZN(n748) );
  NOR2_X1 U798 ( .A1(n747), .A2(n748), .ZN(n749) );
  XOR2_X1 U799 ( .A(KEYINPUT126), .B(n749), .Z(n750) );
  XNOR2_X1 U800 ( .A(n751), .B(n750), .ZN(G69) );
  XOR2_X1 U801 ( .A(KEYINPUT127), .B(n752), .Z(n753) );
  XNOR2_X1 U802 ( .A(n754), .B(n753), .ZN(n758) );
  XNOR2_X1 U803 ( .A(n758), .B(n755), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n757), .A2(n756), .ZN(n762) );
  XNOR2_X1 U805 ( .A(G227), .B(n758), .ZN(n759) );
  NAND2_X1 U806 ( .A1(n759), .A2(G900), .ZN(n760) );
  NAND2_X1 U807 ( .A1(G953), .A2(n760), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n762), .A2(n761), .ZN(G72) );
  XNOR2_X1 U809 ( .A(G134), .B(n763), .ZN(G36) );
  XOR2_X1 U810 ( .A(n764), .B(G125), .Z(n765) );
  XNOR2_X1 U811 ( .A(KEYINPUT37), .B(n765), .ZN(G27) );
  XOR2_X1 U812 ( .A(G137), .B(n766), .Z(G39) );
  XOR2_X1 U813 ( .A(n767), .B(G131), .Z(G33) );
endmodule

