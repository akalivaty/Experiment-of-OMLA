//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923;
  INV_X1    g000(.A(KEYINPUT2), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G148gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n205), .A2(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT78), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n203), .A2(new_n204), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n206), .B(new_n214), .C1(new_n211), .C2(KEYINPUT2), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G120gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G113gat), .ZN(new_n219));
  INV_X1    g018(.A(G113gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G120gat), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT1), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G127gat), .B(G134gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT72), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT72), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(new_n223), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n225), .B1(new_n219), .B2(new_n221), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n224), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n217), .A2(new_n236), .A3(KEYINPUT4), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n232), .A2(new_n234), .B1(new_n223), .B2(new_n222), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n213), .A2(new_n244), .A3(new_n215), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n216), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n237), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n247), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n250), .A2(KEYINPUT79), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT79), .B1(new_n250), .B2(new_n251), .ZN(new_n253));
  OAI221_X1 g052(.A(KEYINPUT5), .B1(new_n241), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n239), .A2(KEYINPUT81), .A3(new_n240), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT81), .B1(new_n239), .B2(new_n240), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n246), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G1gat), .B(G29gat), .Z(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G57gat), .B(G85gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT6), .ZN(new_n266));
  INV_X1    g065(.A(new_n264), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n254), .A2(new_n258), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n259), .A2(KEYINPUT6), .A3(new_n264), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT26), .ZN(new_n273));
  NOR3_X1   g072(.A1(KEYINPUT70), .A2(G169gat), .A3(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n273), .A2(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n274), .A2(new_n273), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n283));
  INV_X1    g082(.A(G183gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT27), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G183gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(G183gat), .ZN(new_n289));
  AOI21_X1  g088(.A(G190gat), .B1(new_n289), .B2(KEYINPUT68), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n282), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(KEYINPUT27), .ZN(new_n292));
  INV_X1    g091(.A(G190gat), .ZN(new_n293));
  AND4_X1   g092(.A1(KEYINPUT28), .A2(new_n289), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n272), .B(new_n281), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  AND2_X1   g095(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(new_n297), .B2(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n272), .A2(KEYINPUT64), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT64), .B1(new_n272), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n298), .B(KEYINPUT65), .C1(new_n300), .C2(new_n301), .ZN(new_n305));
  INV_X1    g104(.A(G169gat), .ZN(new_n306));
  INV_X1    g105(.A(G176gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT23), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(G169gat), .B2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n278), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n308), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT25), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n304), .A2(new_n305), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n308), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n277), .A2(new_n278), .ZN(new_n317));
  INV_X1    g116(.A(new_n296), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT67), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n316), .B(new_n317), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n295), .A2(new_n315), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(G226gat), .A2(G233gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(KEYINPUT29), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  NOR2_X1   g128(.A1(G197gat), .A2(G204gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(G197gat), .A2(G204gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G211gat), .A2(G218gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n330), .A2(new_n332), .B1(new_n334), .B2(KEYINPUT22), .ZN(new_n335));
  NOR2_X1   g134(.A1(G211gat), .A2(G218gat), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT76), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n338));
  INV_X1    g137(.A(G211gat), .ZN(new_n339));
  INV_X1    g138(.A(G218gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n338), .B1(new_n341), .B2(new_n333), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n335), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT22), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n344), .A2(new_n331), .B1(new_n345), .B2(new_n333), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT76), .B1(new_n334), .B2(new_n336), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n338), .A3(new_n333), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n343), .A2(KEYINPUT77), .A3(new_n349), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n329), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n354), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n355), .A2(new_n356), .A3(new_n360), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(KEYINPUT30), .A3(new_n363), .ZN(new_n364));
  OR3_X1    g163(.A1(new_n357), .A2(KEYINPUT30), .A3(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n271), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT88), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n295), .A2(new_n315), .A3(new_n236), .A4(new_n325), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT73), .ZN(new_n370));
  INV_X1    g169(.A(new_n294), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT68), .B1(new_n289), .B2(new_n292), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT68), .B1(new_n284), .B2(KEYINPUT27), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n293), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n371), .B1(new_n375), .B2(new_n282), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n279), .A2(new_n280), .B1(G183gat), .B2(G190gat), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n376), .A2(new_n377), .B1(KEYINPUT25), .B2(new_n324), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT73), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n378), .A2(new_n379), .A3(new_n236), .A4(new_n315), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n326), .A2(new_n243), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n370), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n382), .A2(KEYINPUT74), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT74), .B1(new_n382), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT32), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n384), .B2(new_n385), .ZN(new_n388));
  XOR2_X1   g187(.A(G15gat), .B(G43gat), .Z(new_n389));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n391), .ZN(new_n393));
  OAI221_X1 g192(.A(KEYINPUT32), .B1(new_n387), .B2(new_n393), .C1(new_n384), .C2(new_n385), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n382), .A2(new_n383), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT34), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n392), .A3(new_n394), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(KEYINPUT75), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n395), .A2(new_n402), .A3(new_n397), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT82), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n343), .A2(new_n407), .A3(new_n349), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT3), .B1(new_n408), .B2(KEYINPUT83), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n343), .A2(new_n410), .A3(new_n349), .A4(new_n407), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n217), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n352), .A2(new_n353), .B1(new_n407), .B2(new_n245), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n245), .A2(new_n407), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n245), .A2(KEYINPUT84), .A3(new_n407), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n354), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n405), .B1(new_n216), .B2(KEYINPUT3), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n216), .A2(new_n407), .A3(new_n349), .A4(new_n343), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G22gat), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n414), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n414), .B2(new_n423), .ZN(new_n426));
  OAI21_X1  g225(.A(G78gat), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n414), .A2(new_n423), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G22gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n423), .A3(new_n424), .ZN(new_n430));
  INV_X1    g229(.A(G78gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT31), .B(G50gat), .ZN(new_n433));
  INV_X1    g232(.A(G106gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n427), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n427), .B2(new_n432), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n439), .A2(KEYINPUT35), .ZN(new_n440));
  OR3_X1    g239(.A1(new_n368), .A2(new_n404), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n398), .A2(new_n438), .A3(new_n400), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT89), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n367), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n398), .A2(new_n438), .A3(KEYINPUT89), .A4(new_n400), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n447), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT90), .B1(new_n447), .B2(KEYINPUT35), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n441), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT36), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n398), .B2(new_n400), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n401), .A2(new_n403), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(new_n451), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n438), .B1(new_n271), .B2(new_n366), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n366), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n246), .B1(new_n256), .B2(new_n257), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n251), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n463), .A2(new_n267), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n461), .A2(new_n251), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT39), .B1(new_n250), .B2(new_n251), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n460), .A2(new_n265), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n464), .B(KEYINPUT40), .C1(new_n465), .C2(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n355), .A2(new_n356), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n360), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n329), .A2(KEYINPUT87), .A3(new_n354), .ZN(new_n478));
  OAI211_X1 g277(.A(KEYINPUT37), .B(new_n478), .C1(new_n357), .C2(KEYINPUT87), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT38), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT38), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n357), .B2(KEYINPUT37), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n480), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n271), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n363), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n438), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n474), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n459), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT36), .B1(new_n401), .B2(new_n403), .ZN(new_n490));
  NOR4_X1   g289(.A1(new_n490), .A2(new_n458), .A3(new_n455), .A4(new_n452), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n450), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493));
  INV_X1    g292(.A(G1gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT16), .A3(new_n494), .ZN(new_n495));
  OR2_X1    g294(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n495), .B(new_n496), .C1(new_n494), .C2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n497), .B(new_n498), .Z(new_n499));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT15), .ZN(new_n501));
  INV_X1    g300(.A(G29gat), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT14), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT14), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n500), .A2(KEYINPUT15), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n508), .A2(KEYINPUT91), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n508), .A2(KEYINPUT91), .B1(G29gat), .B2(G36gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n499), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n516), .B(KEYINPUT13), .Z(new_n517));
  AOI21_X1  g316(.A(KEYINPUT94), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n515), .A2(KEYINPUT94), .A3(new_n517), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n514), .A2(KEYINPUT17), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n514), .A2(KEYINPUT17), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n499), .A3(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n499), .A2(new_n514), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n522), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  AOI211_X1 g323(.A(new_n518), .B(new_n519), .C1(KEYINPUT18), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT93), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G197gat), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT11), .B(G169gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n525), .B1(KEYINPUT18), .B2(new_n524), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n532), .B(new_n533), .Z(new_n534));
  AND2_X1   g333(.A1(new_n492), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  INV_X1    g337(.A(G85gat), .ZN(new_n539));
  INV_X1    g338(.A(G92gat), .ZN(new_n540));
  AOI22_X1  g339(.A1(KEYINPUT8), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(G99gat), .B(G106gat), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT97), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n542), .A2(new_n543), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n520), .A2(new_n521), .A3(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT98), .Z(new_n549));
  INV_X1    g348(.A(KEYINPUT41), .ZN(new_n550));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551));
  OAI221_X1 g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .C1(new_n514), .C2(new_n547), .ZN(new_n552));
  XOR2_X1   g351(.A(G190gat), .B(G218gat), .Z(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n550), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT96), .ZN(new_n558));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT99), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n560), .B(KEYINPUT99), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n554), .A2(new_n555), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G57gat), .B(G64gat), .Z(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(new_n431), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(KEYINPUT9), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n499), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT95), .Z(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n203), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n575), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G127gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n566), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n547), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n572), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n572), .A2(new_n546), .A3(new_n544), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(new_n591), .B2(new_n572), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n592), .B1(new_n594), .B2(KEYINPUT10), .ZN(new_n595));
  INV_X1    g394(.A(G230gat), .ZN(new_n596));
  INV_X1    g395(.A(G233gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n598), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G120gat), .B(G148gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT100), .ZN(new_n604));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n604), .B(new_n605), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OR3_X1    g406(.A1(new_n600), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n607), .B1(new_n600), .B2(new_n602), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(KEYINPUT101), .A3(new_n609), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n590), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n535), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(new_n271), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n494), .ZN(G1324gat));
  NAND3_X1  g417(.A1(new_n535), .A2(new_n460), .A3(new_n615), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n619), .A2(G8gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT16), .B(G8gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT42), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(KEYINPUT42), .B2(new_n622), .ZN(G1325gat));
  OAI21_X1  g423(.A(G15gat), .B1(new_n616), .B2(new_n454), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n404), .A2(G15gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(new_n616), .B2(new_n626), .ZN(G1326gat));
  NOR2_X1   g426(.A1(new_n616), .A2(new_n438), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT43), .B(G22gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1327gat));
  NOR3_X1   g429(.A1(new_n368), .A2(new_n404), .A3(new_n440), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n447), .A2(KEYINPUT35), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT90), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n447), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n457), .A2(new_n487), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n565), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n566), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n638), .A2(new_n639), .B1(new_n492), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n614), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n588), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n532), .B(new_n533), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n271), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n502), .B1(new_n648), .B2(KEYINPUT102), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(KEYINPUT102), .B2(new_n648), .ZN(new_n650));
  AND4_X1   g449(.A1(new_n535), .A2(new_n588), .A3(new_n565), .A4(new_n642), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n502), .A3(new_n484), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT45), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(G1328gat));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n503), .A3(new_n460), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(KEYINPUT46), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT103), .ZN(new_n657));
  OAI21_X1  g456(.A(G36gat), .B1(new_n646), .B2(new_n366), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(KEYINPUT46), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(G1329gat));
  NOR2_X1   g459(.A1(new_n404), .A2(G43gat), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n651), .A2(new_n661), .B1(KEYINPUT104), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G43gat), .B1(new_n646), .B2(new_n454), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n662), .A2(KEYINPUT104), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(G1330gat));
  NOR2_X1   g466(.A1(new_n438), .A2(G50gat), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n641), .A2(new_n439), .A3(new_n645), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n651), .A2(new_n668), .B1(new_n669), .B2(G50gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g470(.A1(new_n457), .A2(new_n487), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n450), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n590), .A2(new_n534), .A3(new_n642), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n484), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G57gat), .ZN(G1332gat));
  INV_X1    g476(.A(KEYINPUT49), .ZN(new_n678));
  INV_X1    g477(.A(G64gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n460), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT105), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1333gat));
  INV_X1    g483(.A(new_n454), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n568), .B1(new_n675), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n404), .A2(G71gat), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n675), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g488(.A1(new_n675), .A2(new_n439), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G78gat), .ZN(G1335gat));
  INV_X1    g490(.A(KEYINPUT51), .ZN(new_n692));
  OAI211_X1 g491(.A(KEYINPUT107), .B(new_n565), .C1(new_n636), .C2(new_n637), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n644), .A2(new_n588), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT107), .B1(new_n673), .B2(new_n565), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n692), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n566), .B1(new_n450), .B2(new_n672), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n694), .B1(new_n699), .B2(KEYINPUT107), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n638), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(KEYINPUT51), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n642), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n539), .A3(new_n484), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT85), .B1(new_n454), .B2(new_n456), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(new_n491), .A3(new_n487), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n640), .B1(new_n636), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n694), .A2(new_n642), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n708), .B(new_n709), .C1(new_n699), .C2(KEYINPUT44), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n638), .A2(new_n639), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n713), .A2(KEYINPUT106), .A3(new_n708), .A4(new_n709), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G85gat), .B1(new_n715), .B2(new_n271), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n705), .A2(new_n716), .ZN(G1336gat));
  NAND3_X1  g516(.A1(new_n704), .A2(new_n540), .A3(new_n460), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719));
  OAI21_X1  g518(.A(G92gat), .B1(new_n710), .B2(new_n366), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G92gat), .B1(new_n715), .B2(new_n366), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n723), .B2(new_n719), .ZN(G1337gat));
  INV_X1    g523(.A(G99gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n704), .A2(new_n725), .A3(new_n453), .ZN(new_n726));
  OAI21_X1  g525(.A(G99gat), .B1(new_n715), .B2(new_n454), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1338gat));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n712), .A2(new_n439), .A3(new_n714), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G106gat), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n698), .A2(new_n703), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n614), .A2(new_n434), .A3(new_n439), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT109), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n731), .A2(KEYINPUT108), .A3(G106gat), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n730), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n710), .B2(new_n438), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n641), .A2(KEYINPUT110), .A3(new_n439), .A4(new_n709), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n743), .A3(G106gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n696), .A2(new_n697), .A3(new_n692), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT51), .B1(new_n700), .B2(new_n702), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n737), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n744), .A2(new_n747), .A3(new_n730), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT53), .B1(new_n734), .B2(new_n737), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(new_n751), .A3(new_n744), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n729), .B1(new_n740), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n732), .A2(new_n733), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n739), .A3(new_n747), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT53), .ZN(new_n757));
  AND4_X1   g556(.A1(new_n751), .A2(new_n744), .A3(new_n747), .A4(new_n730), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n751), .B1(new_n750), .B2(new_n744), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n760), .A3(KEYINPUT112), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n754), .A2(new_n761), .ZN(G1339gat));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n600), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n599), .B2(new_n595), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n606), .B1(new_n600), .B2(new_n763), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(KEYINPUT55), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n608), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n765), .A2(new_n766), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n534), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n533), .A2(new_n531), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n515), .A2(new_n517), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n773), .B1(new_n530), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n614), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n566), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n771), .A2(new_n565), .A3(new_n777), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n589), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n590), .A2(new_n534), .A3(new_n614), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n460), .A2(new_n271), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n444), .A2(new_n446), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n220), .B1(new_n789), .B2(new_n644), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n782), .A2(new_n783), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(KEYINPUT113), .A3(new_n438), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n784), .B2(new_n439), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n792), .A2(new_n794), .A3(new_n453), .A4(new_n785), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n534), .A2(G113gat), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(G1340gat));
  OAI21_X1  g597(.A(G120gat), .B1(new_n795), .B2(new_n642), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n787), .A2(new_n218), .A3(new_n788), .A4(new_n614), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT114), .Z(G1341gat));
  OAI21_X1  g601(.A(G127gat), .B1(new_n795), .B2(new_n588), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n588), .A2(G127gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n789), .B2(new_n804), .ZN(G1342gat));
  NOR3_X1   g604(.A1(new_n789), .A2(G134gat), .A3(new_n566), .ZN(new_n806));
  XOR2_X1   g605(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n807));
  OR2_X1    g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G134gat), .B1(new_n795), .B2(new_n566), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(G1343gat));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n685), .B2(new_n438), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n454), .A2(KEYINPUT119), .A3(new_n439), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n787), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(G141gat), .A3(new_n644), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(KEYINPUT58), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n685), .A2(new_n786), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n791), .A2(new_n439), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(KEYINPUT57), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821));
  INV_X1    g620(.A(new_n783), .ZN(new_n822));
  INV_X1    g621(.A(new_n781), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n770), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n608), .A3(new_n767), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n778), .B1(new_n644), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n565), .B1(new_n827), .B2(KEYINPUT117), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n822), .B1(new_n830), .B2(new_n589), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n821), .B1(new_n831), .B2(new_n439), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n820), .A2(new_n644), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n817), .B1(new_n207), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n820), .ZN(new_n835));
  INV_X1    g634(.A(new_n832), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(KEYINPUT118), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n820), .B2(new_n832), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n534), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n816), .B1(new_n840), .B2(G141gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n834), .B1(new_n841), .B2(new_n842), .ZN(G1344gat));
  INV_X1    g642(.A(new_n815), .ZN(new_n844));
  INV_X1    g643(.A(G148gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n614), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n837), .A2(new_n614), .A3(new_n839), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n845), .A2(KEYINPUT59), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g648(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n850));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n831), .B2(new_n439), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n784), .A2(new_n821), .A3(new_n438), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n614), .A3(new_n818), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n850), .B1(new_n854), .B2(G148gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n846), .B1(new_n849), .B2(new_n855), .ZN(G1345gat));
  NAND4_X1  g655(.A1(new_n837), .A2(G155gat), .A3(new_n839), .A4(new_n589), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n203), .B1(new_n815), .B2(new_n588), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(KEYINPUT121), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1346gat));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n204), .A3(new_n565), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n837), .A2(new_n565), .A3(new_n839), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n204), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n484), .A2(new_n366), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n792), .A2(new_n794), .A3(new_n453), .A4(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n306), .A3(new_n644), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n791), .A2(new_n788), .A3(new_n867), .ZN(new_n870));
  AOI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n534), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n869), .A2(new_n871), .ZN(G1348gat));
  OAI21_X1  g671(.A(G176gat), .B1(new_n868), .B2(new_n642), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n307), .A3(new_n614), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1349gat));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(KEYINPUT60), .ZN(new_n877));
  OAI21_X1  g676(.A(G183gat), .B1(new_n868), .B2(new_n588), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n870), .A2(new_n289), .A3(new_n292), .A4(new_n589), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(KEYINPUT60), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n880), .B(new_n881), .Z(G1350gat));
  NAND3_X1  g681(.A1(new_n870), .A2(new_n293), .A3(new_n565), .ZN(new_n883));
  OAI21_X1  g682(.A(G190gat), .B1(new_n868), .B2(new_n566), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT61), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n884), .A2(KEYINPUT61), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(G1351gat));
  NAND2_X1  g687(.A1(new_n454), .A2(new_n867), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n819), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(KEYINPUT123), .B(G197gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n534), .A3(new_n891), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n889), .B(KEYINPUT124), .Z(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n853), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n644), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n891), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n853), .A2(new_n534), .A3(new_n894), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(KEYINPUT125), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n892), .B1(new_n898), .B2(new_n901), .ZN(G1352gat));
  INV_X1    g701(.A(G204gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n890), .A2(new_n903), .A3(new_n614), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT126), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(KEYINPUT126), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(KEYINPUT62), .A3(new_n906), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n853), .A2(new_n614), .A3(new_n894), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n909), .B(new_n910), .C1(new_n903), .C2(new_n911), .ZN(G1353gat));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n339), .A3(new_n589), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n589), .B(new_n894), .C1(new_n851), .C2(new_n852), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n914), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT63), .B1(new_n914), .B2(G211gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n913), .B(KEYINPUT127), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1354gat));
  OAI21_X1  g720(.A(G218gat), .B1(new_n895), .B2(new_n566), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n890), .A2(new_n340), .A3(new_n565), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1355gat));
endmodule


