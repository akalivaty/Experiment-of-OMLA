//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(KEYINPUT68), .A3(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n463), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n469), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n478));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n472), .A2(KEYINPUT67), .A3(new_n473), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G125), .ZN(new_n483));
  NAND2_X1  g058(.A1(G113), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n475), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n477), .A2(new_n485), .ZN(G160));
  INV_X1    g061(.A(new_n476), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n474), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(G162));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n475), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI22_X1  g072(.A1(new_n489), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n481), .A2(new_n482), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n475), .C1(new_n479), .C2(new_n480), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n502), .B1(KEYINPUT4), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT69), .A4(new_n500), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n498), .B1(new_n504), .B2(new_n505), .ZN(G164));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  XOR2_X1   g082(.A(KEYINPUT5), .B(G543), .Z(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G88), .B1(new_n518), .B2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(G166));
  NAND2_X1  g097(.A1(new_n518), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n513), .A2(new_n514), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT5), .B(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n523), .B(new_n525), .C1(new_n526), .C2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT71), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n527), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n534), .A2(new_n535), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G651), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n542), .A2(new_n535), .B1(new_n529), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n539), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n518), .B2(G53), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n518), .A2(new_n553), .A3(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n508), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n539), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n563), .B1(new_n562), .B2(new_n561), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n554), .A2(new_n555), .B1(G91), .B2(new_n516), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n558), .A2(new_n564), .A3(new_n565), .ZN(G299));
  OR2_X1    g141(.A1(new_n537), .A2(new_n540), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT74), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n537), .A2(KEYINPUT74), .A3(new_n540), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT75), .B1(new_n529), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n516), .A2(new_n576), .A3(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n528), .A2(G74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n518), .B2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n516), .A2(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n518), .A2(G48), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n539), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n589), .A2(new_n535), .B1(new_n529), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n539), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(KEYINPUT76), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(KEYINPUT76), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(new_n516), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n508), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n518), .B2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT78), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n605), .A2(new_n606), .B1(new_n607), .B2(KEYINPUT77), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(KEYINPUT77), .B2(new_n607), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(KEYINPUT77), .B2(new_n607), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  INV_X1    g186(.A(G299), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G297));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G280));
  INV_X1    g189(.A(new_n605), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  INV_X1    g192(.A(new_n547), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n606), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n605), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n487), .A2(G135), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT79), .Z(new_n624));
  OAI21_X1  g199(.A(KEYINPUT80), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G111), .B2(new_n475), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n475), .A2(G111), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n463), .B1(new_n627), .B2(KEYINPUT80), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n490), .A2(G123), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT81), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2096), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n481), .A2(new_n482), .A3(new_n464), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(G401));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n656), .B(KEYINPUT17), .Z(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n654), .B2(new_n662), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n664), .B2(new_n655), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(G2100), .Z(new_n666));
  XOR2_X1   g241(.A(KEYINPUT85), .B(G2096), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1981), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G4), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n615), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1348), .ZN(new_n690));
  NOR2_X1   g265(.A1(G29), .A2(G35), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G162), .B2(G29), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT29), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G2090), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G26), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  OR2_X1    g273(.A1(G104), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT93), .ZN(new_n701));
  INV_X1    g276(.A(G128), .ZN(new_n702));
  INV_X1    g277(.A(G140), .ZN(new_n703));
  OAI22_X1  g278(.A1(new_n702), .A2(new_n489), .B1(new_n476), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n698), .B1(new_n705), .B2(new_n696), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G2067), .ZN(new_n707));
  INV_X1    g282(.A(G32), .ZN(new_n708));
  AOI21_X1  g283(.A(KEYINPUT95), .B1(new_n696), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n487), .A2(G141), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT26), .Z(new_n713));
  INV_X1    g288(.A(G129), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n489), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n464), .A2(G105), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n711), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G29), .ZN(new_n718));
  MUX2_X1   g293(.A(KEYINPUT95), .B(new_n709), .S(new_n718), .Z(new_n719));
  XOR2_X1   g294(.A(KEYINPUT27), .B(G1996), .Z(new_n720));
  AOI21_X1  g295(.A(new_n707), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n696), .B1(new_n722), .B2(G34), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G160), .B2(G29), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n721), .B(new_n727), .C1(new_n720), .C2(new_n719), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G33), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n481), .A2(new_n482), .A3(G127), .ZN(new_n732));
  INV_X1    g307(.A(G115), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n463), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2105), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n487), .A2(G139), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n730), .B(new_n731), .C1(new_n741), .C2(new_n696), .ZN(new_n742));
  INV_X1    g317(.A(G2072), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n687), .A2(G19), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n547), .B2(new_n687), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1341), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n742), .A2(new_n743), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n687), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n687), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n749), .C1(G1961), .C2(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n728), .A2(new_n744), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n687), .A2(G20), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1956), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n696), .A2(G27), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G164), .B2(new_n696), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2078), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n631), .A2(G29), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n765), .A2(KEYINPUT96), .A3(G28), .ZN(new_n766));
  AOI21_X1  g341(.A(KEYINPUT96), .B1(new_n765), .B2(G28), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n696), .B1(new_n765), .B2(G28), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n751), .B2(G1961), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n687), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n687), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n764), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT97), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n695), .A2(new_n753), .A3(new_n763), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G166), .A2(new_n687), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n687), .A2(G22), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G1971), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n779), .A2(G1971), .A3(new_n780), .ZN(new_n785));
  OR3_X1    g360(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n784), .B1(new_n783), .B2(new_n785), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n687), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(G288), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n687), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT33), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1976), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n687), .A2(G6), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n587), .B2(new_n687), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT90), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n788), .A2(new_n789), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n794), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n786), .A2(new_n787), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT34), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n687), .A2(G24), .ZN(new_n804));
  INV_X1    g379(.A(G290), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n687), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1986), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n696), .A2(G25), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT87), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n487), .A2(G131), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n490), .A2(G119), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n475), .A2(G107), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT88), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT88), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n809), .B1(new_n817), .B2(G29), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT89), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n807), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n800), .A2(new_n803), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n800), .A2(new_n803), .A3(new_n825), .A4(new_n822), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n778), .B1(new_n824), .B2(new_n826), .ZN(G311));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n828));
  XNOR2_X1  g403(.A(G311), .B(new_n828), .ZN(G150));
  NOR2_X1   g404(.A1(new_n605), .A2(new_n616), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n832), .A2(new_n535), .B1(new_n529), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n539), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n547), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n831), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  AOI21_X1  g416(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  INV_X1    g418(.A(new_n837), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(G145));
  NAND2_X1  g422(.A1(new_n501), .A2(new_n502), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n505), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n498), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n705), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(new_n717), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n741), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n717), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n735), .A2(KEYINPUT100), .A3(new_n740), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n490), .A2(G130), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n475), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(G142), .B2(new_n487), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(new_n634), .Z(new_n866));
  INV_X1    g441(.A(new_n817), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n860), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n631), .B(G162), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G160), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n871), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g451(.A(new_n620), .B(new_n838), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n599), .A2(new_n603), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(G299), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n612), .A2(new_n604), .A3(KEYINPUT102), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(G299), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT101), .B1(new_n879), .B2(G299), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n612), .A2(new_n604), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n881), .B(new_n880), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n889), .B2(new_n884), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n877), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n889), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n877), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n805), .A2(new_n791), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n791), .B1(new_n595), .B2(new_n596), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(KEYINPUT103), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  NOR2_X1   g475(.A1(G290), .A2(G288), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(new_n897), .ZN(new_n902));
  XNOR2_X1  g477(.A(G166), .B(new_n587), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n905), .B(new_n900), .C1(new_n901), .C2(new_n897), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n894), .B1(new_n891), .B2(new_n893), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n895), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n895), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g488(.A(G868), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n844), .A2(new_n606), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(G295));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n915), .ZN(G331));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  OR3_X1    g493(.A1(G168), .A2(new_n567), .A3(KEYINPUT105), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n568), .A2(G168), .A3(new_n569), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT105), .B1(G168), .B2(new_n567), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n839), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n919), .A2(new_n838), .A3(new_n920), .A4(new_n921), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n880), .A2(new_n881), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n882), .A2(new_n887), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n879), .A2(KEYINPUT101), .A3(G299), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n926), .A2(new_n929), .B1(new_n839), .B2(new_n922), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n924), .B(KEYINPUT106), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n890), .A2(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n932), .B2(new_n907), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n923), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n883), .A2(KEYINPUT41), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n926), .A2(new_n929), .A3(new_n884), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n924), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n933), .B(new_n934), .C1(new_n940), .C2(new_n907), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n890), .A2(new_n925), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n930), .A2(new_n931), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n908), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n934), .B1(new_n933), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI211_X1 g523(.A(KEYINPUT107), .B(new_n934), .C1(new_n933), .C2(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n918), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n942), .A2(new_n943), .A3(new_n907), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n873), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n907), .B1(new_n938), .B2(new_n939), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n933), .A2(new_n945), .A3(new_n934), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n950), .B1(new_n958), .B2(new_n959), .ZN(G397));
  AOI21_X1  g535(.A(G1384), .B1(new_n850), .B2(new_n851), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n477), .A2(new_n485), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G2067), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n705), .A2(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n701), .A2(new_n704), .A3(G2067), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n717), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G1996), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n966), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n966), .A2(G1996), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT109), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n976), .B2(new_n717), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n817), .B(new_n820), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n977), .B1(new_n966), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n966), .ZN(new_n980));
  XNOR2_X1  g555(.A(G290), .B(G1986), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n587), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT113), .B1(new_n582), .B2(new_n583), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n586), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n582), .A2(KEYINPUT113), .A3(new_n583), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n988), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n992), .A2(new_n586), .A3(new_n986), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n993), .A2(KEYINPUT114), .A3(new_n984), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n983), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n990), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT114), .B1(new_n993), .B2(new_n984), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n997), .A3(KEYINPUT49), .A4(new_n985), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n961), .A2(new_n965), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G8), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(G1976), .B2(new_n791), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1001), .B(new_n1007), .C1(new_n1006), .C2(G288), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1010), .B(new_n965), .C1(new_n961), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n852), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1016), .B2(new_n965), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1015), .A2(new_n1017), .A3(G2090), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n487), .A2(G137), .B1(new_n467), .B2(new_n468), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n483), .A2(new_n484), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1019), .B(G40), .C1(new_n1020), .C2(new_n475), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n963), .B1(G164), .B2(G1384), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1971), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT116), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1016), .A2(new_n965), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1014), .A4(new_n1012), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1024), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(G8), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G166), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT55), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1009), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1021), .A2(G2084), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1016), .A2(new_n1014), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n962), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1966), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1046), .A2(new_n1034), .A3(G286), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1021), .A2(G2090), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(KEYINPUT111), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1024), .B1(new_n1050), .B2(KEYINPUT111), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(G8), .A4(new_n1036), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1034), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1054), .B1(new_n1057), .B2(new_n1036), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1038), .B(new_n1047), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(KEYINPUT111), .A3(new_n1048), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1031), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1050), .A2(KEYINPUT111), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(new_n1036), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT112), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1055), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1057), .A2(new_n1036), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1009), .A2(new_n1060), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1068), .A2(new_n1047), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1061), .A2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1044), .A2(G286), .A3(new_n1045), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n1073), .B2(new_n1034), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1062), .A2(new_n1039), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1045), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1078), .B2(G286), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(G168), .A3(new_n1077), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G8), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1074), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT123), .B1(new_n1082), .B2(KEYINPUT62), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1074), .B(new_n1084), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1062), .A2(new_n965), .ZN(new_n1086));
  INV_X1    g661(.A(G1961), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1089));
  INV_X1    g664(.A(G2078), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1023), .A2(new_n1089), .A3(new_n1090), .A4(new_n965), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1022), .A2(KEYINPUT53), .A3(new_n1090), .A4(new_n1023), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(G301), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1085), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1083), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1068), .A2(new_n1038), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1082), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1068), .A2(new_n1009), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1002), .A2(new_n1006), .A3(new_n791), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1000), .B1(new_n1103), .B2(new_n985), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1072), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1961), .B1(new_n1062), .B2(new_n965), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n570), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1107), .B1(new_n1096), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT122), .B(new_n1107), .C1(new_n1096), .C2(new_n1110), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(G171), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT51), .B1(new_n1046), .B2(G168), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(G8), .A3(new_n1080), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1117), .A2(new_n1118), .B1(new_n1120), .B2(new_n1074), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1115), .A2(new_n1068), .A3(new_n1038), .A4(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n758), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1123));
  XOR2_X1   g698(.A(G299), .B(KEYINPUT57), .Z(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1022), .A2(new_n1023), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n999), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n967), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1021), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(G1348), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(KEYINPUT117), .A3(new_n879), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1124), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT117), .B1(new_n1131), .B2(new_n879), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1127), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1127), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1135), .A2(KEYINPUT118), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1133), .A2(new_n1142), .A3(new_n1134), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1140), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1139), .B1(new_n1144), .B2(KEYINPUT61), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1143), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1142), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1127), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(KEYINPUT119), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1135), .A2(KEYINPUT61), .A3(new_n1127), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1135), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n1127), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT60), .B(new_n1129), .C1(new_n1130), .C2(G1348), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(G1996), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1022), .A2(new_n1158), .A3(new_n1023), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT58), .B(G1341), .Z(new_n1160));
  NAND2_X1  g735(.A1(new_n999), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1157), .B1(new_n1162), .B2(new_n547), .ZN(new_n1163));
  AOI211_X1 g738(.A(KEYINPUT59), .B(new_n618), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1156), .A2(new_n879), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1131), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1156), .A2(new_n879), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1145), .A2(new_n1150), .A3(new_n1155), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1122), .B1(new_n1138), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n982), .B1(new_n1106), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n970), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n980), .B1(new_n1173), .B2(new_n971), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n975), .A2(KEYINPUT46), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n975), .A2(KEYINPUT46), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n867), .A2(new_n820), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT124), .Z(new_n1184));
  AOI21_X1  g759(.A(new_n969), .B1(new_n977), .B2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n966), .A2(G290), .A3(G1986), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT127), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT48), .ZN(new_n1188));
  OAI22_X1  g763(.A1(new_n1185), .A2(new_n966), .B1(new_n979), .B2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1181), .A2(new_n1182), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1172), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g766(.A1(G229), .A2(G227), .A3(new_n461), .A4(G401), .ZN(new_n1193));
  OAI211_X1 g767(.A(new_n875), .B(new_n1193), .C1(new_n948), .C2(new_n949), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


