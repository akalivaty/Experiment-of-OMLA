//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n191));
  INV_X1    g005(.A(G113), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(KEYINPUT66), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(KEYINPUT2), .B2(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT2), .A2(G113), .ZN(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G119), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n196), .B2(new_n197), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n190), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n194), .A2(KEYINPUT2), .A3(G113), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT66), .B1(new_n191), .B2(new_n192), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n198), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(KEYINPUT67), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT4), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT77), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G107), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT77), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n210), .B(G101), .C1(new_n216), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(G101), .B1(new_n216), .B2(new_n222), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n218), .A2(KEYINPUT77), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n219), .B1(new_n225), .B2(new_n221), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n212), .A2(new_n214), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n217), .A4(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n209), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n232), .B(G113), .C1(KEYINPUT5), .C2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT79), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n221), .A2(new_n217), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G101), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n229), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n236), .B1(new_n229), .B2(new_n238), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n207), .B(new_n235), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT6), .ZN(new_n243));
  XNOR2_X1  g057(.A(G110), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n231), .A2(new_n241), .A3(new_n244), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT6), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n244), .B1(new_n231), .B2(new_n241), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n189), .B(new_n246), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n249), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n251), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n247), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G224), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G953), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(G128), .ZN(new_n258));
  INV_X1    g072(.A(G125), .ZN(new_n259));
  OR2_X1    g073(.A1(KEYINPUT65), .A2(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT65), .A2(G128), .ZN(new_n261));
  INV_X1    g075(.A(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G143), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n260), .A2(new_n261), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n258), .B(new_n259), .C1(new_n264), .C2(new_n256), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT0), .B(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n256), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n265), .A2(new_n266), .B1(new_n274), .B2(G125), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n273), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n276), .A2(KEYINPUT85), .A3(new_n259), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n255), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n265), .A2(new_n266), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(G125), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n255), .ZN(new_n282));
  INV_X1    g096(.A(new_n277), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n253), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G210), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n278), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n281), .A2(new_n289), .A3(new_n282), .A4(new_n283), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n293), .A2(new_n247), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n244), .B(KEYINPUT8), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OR2_X1    g110(.A1(new_n241), .A2(KEYINPUT86), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n229), .A2(new_n238), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n235), .A2(new_n207), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n241), .A2(KEYINPUT86), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(G902), .B1(new_n294), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(new_n288), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n288), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n285), .B1(new_n250), .B2(new_n252), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n293), .A2(new_n247), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n301), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n305), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n188), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT87), .ZN(new_n312));
  NOR2_X1   g126(.A1(G475), .A2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G113), .B(G122), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(new_n213), .ZN(new_n316));
  OR2_X1    g130(.A1(KEYINPUT68), .A2(G953), .ZN(new_n317));
  INV_X1    g131(.A(G237), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT68), .A2(G953), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n317), .A2(G214), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n267), .ZN(new_n321));
  AND2_X1   g135(.A1(KEYINPUT68), .A2(G953), .ZN(new_n322));
  NOR2_X1   g136(.A1(KEYINPUT68), .A2(G953), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(G143), .A3(G214), .A4(new_n318), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(KEYINPUT18), .A2(G131), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(new_n262), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n326), .B2(new_n327), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n321), .B2(new_n325), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n321), .A2(new_n325), .A3(new_n334), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n259), .A2(G140), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT16), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n259), .A2(KEYINPUT16), .A3(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n262), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(G146), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(KEYINPUT72), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n345), .A2(new_n349), .A3(new_n262), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n348), .A2(new_n350), .B1(new_n335), .B2(KEYINPUT17), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n339), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n326), .A2(KEYINPUT17), .A3(G131), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n347), .A2(KEYINPUT72), .ZN(new_n355));
  AOI21_X1  g169(.A(G146), .B1(new_n343), .B2(new_n344), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n350), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n354), .B(new_n352), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n316), .B(new_n333), .C1(new_n353), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n316), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n329), .B(KEYINPUT19), .Z(new_n363));
  OAI21_X1  g177(.A(new_n347), .B1(new_n363), .B2(G146), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n336), .B2(new_n338), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n362), .B1(new_n365), .B2(new_n332), .ZN(new_n366));
  AOI211_X1 g180(.A(KEYINPUT20), .B(new_n314), .C1(new_n361), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n366), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n361), .A2(KEYINPUT89), .A3(new_n366), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n313), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n367), .B1(new_n372), .B2(KEYINPUT20), .ZN(new_n373));
  INV_X1    g187(.A(G475), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT88), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n359), .A3(new_n339), .ZN(new_n377));
  AOI211_X1 g191(.A(KEYINPUT90), .B(new_n316), .C1(new_n377), .C2(new_n333), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n333), .B1(new_n353), .B2(new_n360), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n362), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n361), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n374), .B1(new_n382), .B2(new_n307), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G478), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT15), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(KEYINPUT15), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT9), .B(G234), .ZN(new_n393));
  INV_X1    g207(.A(G217), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n393), .A2(new_n394), .A3(G953), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n260), .A2(G143), .A3(new_n261), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n267), .A2(G128), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G134), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(G134), .A3(new_n398), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT13), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n404), .A2(KEYINPUT92), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n400), .B1(KEYINPUT92), .B2(new_n404), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n397), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT91), .ZN(new_n410));
  INV_X1    g224(.A(G122), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(G116), .ZN(new_n412));
  INV_X1    g226(.A(G116), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT91), .A3(G122), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n413), .A2(G122), .ZN(new_n417));
  OAI21_X1  g231(.A(G107), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n415), .B(new_n220), .C1(new_n413), .C2(G122), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n401), .A2(new_n402), .A3(new_n407), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n409), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n401), .A2(new_n402), .A3(new_n419), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT14), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n412), .B2(new_n414), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(new_n417), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT93), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n425), .B2(new_n417), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n416), .A2(new_n424), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n423), .B1(new_n431), .B2(G107), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n396), .B1(new_n422), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n409), .A2(new_n420), .A3(new_n421), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n426), .A2(KEYINPUT93), .B1(new_n416), .B2(new_n424), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n220), .B1(new_n435), .B2(new_n429), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n434), .B(new_n395), .C1(new_n436), .C2(new_n423), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n392), .B1(new_n438), .B2(new_n307), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI211_X1 g254(.A(G902), .B(new_n391), .C1(new_n433), .C2(new_n437), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n385), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G953), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G952), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(G234), .B2(G237), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n307), .B(new_n324), .C1(G234), .C2(G237), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(G898), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n312), .A2(new_n444), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n324), .A2(G221), .A3(G234), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G137), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n329), .A2(new_n262), .ZN(new_n456));
  INV_X1    g270(.A(G128), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G119), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT23), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n233), .B2(G128), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n260), .A2(G119), .A3(new_n261), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n459), .B(new_n461), .C1(new_n462), .C2(new_n460), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G110), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT24), .B(G110), .Z(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n462), .B2(new_n459), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n456), .B(new_n347), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n462), .A3(new_n459), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(G110), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n348), .A2(new_n350), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n467), .A2(new_n470), .A3(KEYINPUT73), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT73), .B1(new_n467), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n455), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n455), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n470), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT73), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n307), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT25), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n473), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n477), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n394), .B1(G234), .B2(new_n307), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n473), .A2(new_n477), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n485), .A2(G902), .A3(new_n483), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(KEYINPUT74), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT74), .ZN(new_n489));
  INV_X1    g303(.A(new_n483), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n480), .B2(new_n481), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n489), .B1(new_n491), .B2(new_n486), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G472), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n324), .A2(G210), .A3(new_n318), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT27), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G101), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n495), .A2(KEYINPUT27), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(KEYINPUT27), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT64), .ZN(new_n505));
  INV_X1    g319(.A(G137), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(KEYINPUT11), .A2(G134), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT64), .A2(G137), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(KEYINPUT11), .A2(G134), .ZN(new_n511));
  NOR2_X1   g325(.A1(KEYINPUT11), .A2(G134), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(G137), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n510), .A2(new_n334), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n334), .B1(new_n510), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n276), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n513), .A3(new_n334), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n507), .A2(new_n400), .A3(new_n509), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n334), .B1(G134), .B2(G137), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n260), .A2(new_n261), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT1), .B1(new_n267), .B2(G146), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n256), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND4_X1   g337(.A1(new_n257), .A2(new_n263), .A3(new_n268), .A4(G128), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n517), .B(new_n520), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n201), .A2(new_n516), .A3(new_n208), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n503), .B1(new_n504), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT29), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n516), .A2(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n209), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n504), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n307), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n530), .A2(new_n533), .A3(new_n526), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT28), .B1(new_n530), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n527), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT29), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n529), .A2(KEYINPUT30), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n516), .A2(new_n525), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n538), .A2(new_n540), .B1(new_n201), .B2(new_n208), .ZN(new_n541));
  INV_X1    g355(.A(new_n526), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n503), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n536), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n532), .B1(new_n544), .B2(KEYINPUT70), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n536), .A2(new_n546), .A3(new_n543), .A4(new_n537), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n494), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n516), .A2(new_n525), .A3(new_n539), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n539), .B1(new_n516), .B2(new_n525), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n209), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n503), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n526), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT31), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n552), .A2(new_n556), .A3(new_n553), .A4(new_n526), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n542), .A2(KEYINPUT28), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n209), .A2(new_n529), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n504), .B1(new_n559), .B2(KEYINPUT69), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n530), .A2(new_n533), .A3(new_n526), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n555), .B(new_n557), .C1(new_n562), .C2(new_n553), .ZN(new_n563));
  NOR2_X1   g377(.A1(G472), .A2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT32), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT32), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n548), .A2(new_n549), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n544), .A2(KEYINPUT70), .ZN(new_n570));
  INV_X1    g384(.A(new_n532), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n547), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G472), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT71), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n493), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(KEYINPUT80), .A2(KEYINPUT12), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n298), .A2(KEYINPUT79), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n229), .A2(new_n236), .A3(new_n238), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n258), .B1(new_n264), .B2(new_n256), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n522), .A2(KEYINPUT78), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n263), .A2(new_n586), .A3(KEYINPUT1), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(G128), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n524), .B1(new_n588), .B2(new_n269), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n589), .A2(new_n298), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n514), .A2(new_n515), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n579), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n579), .ZN(new_n597));
  AOI211_X1 g411(.A(new_n597), .B(new_n594), .C1(new_n584), .C2(new_n590), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(KEYINPUT10), .B(new_n582), .C1(new_n239), .C2(new_n240), .ZN(new_n600));
  INV_X1    g414(.A(new_n592), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n230), .A2(new_n223), .A3(new_n276), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n589), .B2(new_n298), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n324), .A2(G227), .ZN(new_n606));
  XNOR2_X1  g420(.A(G110), .B(G140), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n599), .A2(KEYINPUT82), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT82), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n239), .A2(new_n240), .A3(new_n582), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n589), .A2(new_n298), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n595), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n597), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n591), .A2(new_n579), .A3(new_n595), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n611), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n613), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n602), .A2(new_n604), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n582), .A2(KEYINPUT10), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n580), .B2(new_n581), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n592), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n605), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT83), .ZN(new_n627));
  INV_X1    g441(.A(new_n610), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n631));
  OAI22_X1  g445(.A1(new_n612), .A2(new_n621), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(G469), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n307), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n307), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n620), .A2(new_n625), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n622), .A2(new_n624), .A3(new_n592), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n617), .B2(new_n618), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n637), .B1(new_n639), .B2(new_n610), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT81), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n628), .B1(new_n599), .B2(new_n638), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT81), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n637), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n641), .A2(G469), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n634), .A2(new_n636), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(G221), .B1(new_n393), .B2(G902), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n576), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n452), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G101), .ZN(G3));
  AND2_X1   g465(.A1(new_n488), .A2(new_n492), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n563), .A2(new_n307), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(G472), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n565), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n652), .A2(new_n647), .A3(new_n646), .A4(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT33), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n438), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT95), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n437), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n437), .A2(new_n660), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT33), .A4(new_n433), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT95), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n438), .A2(new_n664), .A3(new_n657), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n386), .A2(G902), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n659), .A2(new_n663), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n438), .A2(new_n307), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n386), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n373), .B2(new_n383), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n288), .B1(new_n287), .B2(new_n303), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n306), .A2(new_n309), .A3(new_n305), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n451), .B(new_n187), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n656), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n213), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  NAND2_X1  g492(.A1(new_n382), .A2(new_n307), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G475), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n361), .A2(KEYINPUT89), .A3(new_n366), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT89), .B1(new_n361), .B2(new_n366), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n681), .A2(new_n682), .A3(new_n314), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n372), .A2(KEYINPUT20), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n680), .B(new_n443), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n656), .A2(new_n674), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT35), .B(G107), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G9));
  INV_X1    g504(.A(new_n648), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n474), .A2(KEYINPUT36), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n475), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n483), .A2(G902), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n484), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n691), .A2(new_n655), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n452), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  INV_X1    g515(.A(new_n447), .ZN(new_n702));
  INV_X1    g516(.A(new_n448), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(G900), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT98), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n687), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n691), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n566), .A2(new_n568), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n572), .A2(new_n549), .A3(G472), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n548), .A2(new_n549), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n311), .B(new_n696), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n701), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n712), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(KEYINPUT99), .A3(new_n691), .A4(new_n706), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  NOR2_X1   g531(.A1(new_n541), .A2(new_n542), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n503), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n503), .A2(new_n530), .A3(new_n526), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n307), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n708), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n188), .A3(new_n696), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n443), .B1(new_n373), .B2(new_n383), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n304), .A2(new_n310), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n727), .B1(new_n304), .B2(new_n310), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n724), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT101), .Z(new_n733));
  XOR2_X1   g547(.A(new_n705), .B(KEYINPUT39), .Z(new_n734));
  NAND2_X1  g548(.A1(new_n691), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT40), .Z(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT102), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G143), .ZN(G45));
  INV_X1    g553(.A(new_n705), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n670), .B(new_n740), .C1(new_n373), .C2(new_n383), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n648), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n714), .A2(KEYINPUT103), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  INV_X1    g558(.A(new_n741), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n646), .A3(new_n647), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n746), .B2(new_n712), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G146), .ZN(G48));
  NOR2_X1   g563(.A1(new_n674), .A2(new_n671), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT82), .B1(new_n599), .B2(new_n611), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n619), .A2(new_n620), .A3(new_n613), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n626), .A2(new_n628), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT83), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n751), .A2(new_n752), .B1(new_n754), .B2(new_n629), .ZN(new_n755));
  OAI21_X1  g569(.A(G469), .B1(new_n755), .B2(G902), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n634), .A3(new_n757), .A4(new_n647), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n647), .A3(new_n634), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT104), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n575), .A2(new_n750), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT41), .B(G113), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G15));
  NOR2_X1   g577(.A1(new_n674), .A2(new_n687), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n575), .A2(new_n764), .A3(new_n758), .A4(new_n760), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G116), .ZN(G18));
  NAND3_X1  g580(.A1(new_n760), .A2(new_n311), .A3(new_n758), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT105), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT105), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n760), .A2(new_n769), .A3(new_n311), .A4(new_n758), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n710), .A2(new_n711), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n491), .B1(new_n694), .B2(new_n693), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n444), .A3(new_n451), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G119), .ZN(G21));
  OAI21_X1  g591(.A(new_n187), .B1(new_n672), .B2(new_n673), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n725), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n491), .A2(new_n486), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n503), .B1(new_n558), .B2(new_n531), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n555), .A2(new_n557), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n564), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n654), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n450), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n760), .A2(new_n779), .A3(new_n758), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G122), .ZN(G24));
  NAND2_X1  g601(.A1(new_n654), .A2(new_n783), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n741), .A2(new_n773), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n771), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G125), .ZN(G27));
  NAND3_X1  g605(.A1(new_n574), .A2(new_n708), .A3(new_n709), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n780), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n633), .B1(new_n640), .B2(new_n307), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n751), .A2(new_n752), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n754), .A2(new_n629), .ZN(new_n797));
  AOI21_X1  g611(.A(G902), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n795), .B1(new_n798), .B2(new_n633), .ZN(new_n799));
  INV_X1    g613(.A(new_n647), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n188), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n304), .A2(new_n310), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n794), .A2(KEYINPUT42), .A3(new_n745), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n792), .A3(new_n745), .A4(new_n652), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(KEYINPUT106), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT42), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n805), .B2(KEYINPUT106), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n804), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G131), .ZN(G33));
  NAND3_X1  g624(.A1(new_n575), .A2(new_n706), .A3(new_n803), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT107), .B(G134), .Z(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G36));
  OR3_X1    g627(.A1(new_n655), .A2(KEYINPUT109), .A3(new_n773), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT109), .B1(new_n655), .B2(new_n773), .ZN(new_n815));
  INV_X1    g629(.A(new_n367), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n683), .B2(new_n684), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n680), .A3(new_n670), .ZN(new_n818));
  AND2_X1   g632(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n819));
  NOR2_X1   g633(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n820), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n384), .A2(new_n670), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n814), .A2(new_n815), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT44), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT110), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT45), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n640), .A2(KEYINPUT81), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n643), .B1(new_n642), .B2(new_n637), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n640), .A2(new_n829), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n633), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n635), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n634), .B1(new_n835), .B2(KEYINPUT46), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n832), .A2(new_n834), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n837), .A2(KEYINPUT46), .A3(new_n636), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n647), .B(new_n734), .C1(new_n836), .C2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n826), .A2(KEYINPUT44), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n672), .A2(new_n673), .A3(new_n188), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n828), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G137), .ZN(G39));
  OAI21_X1  g658(.A(new_n647), .B1(new_n836), .B2(new_n838), .ZN(new_n845));
  XNOR2_X1  g659(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n647), .B(new_n846), .C1(new_n836), .C2(new_n838), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n842), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n792), .A3(new_n652), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n745), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G140), .ZN(G42));
  NAND2_X1  g668(.A1(new_n761), .A2(new_n765), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT113), .B1(new_n440), .B2(new_n442), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n439), .A2(new_n441), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n817), .A3(new_n680), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n671), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n311), .A2(KEYINPUT87), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT87), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n863), .B(new_n188), .C1(new_n304), .C2(new_n310), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n451), .B(new_n861), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n786), .B1(new_n865), .B2(new_n656), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n855), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n452), .B1(new_n649), .B2(new_n697), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n776), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n685), .A2(new_n686), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n859), .A2(new_n705), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n680), .A2(new_n842), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n774), .A2(new_n872), .A3(new_n691), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n789), .A2(new_n803), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n873), .A2(new_n811), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n809), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n771), .A2(new_n789), .B1(new_n713), .B2(new_n715), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n773), .A2(new_n647), .A3(new_n740), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n723), .A2(new_n879), .A3(new_n799), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n743), .A2(new_n747), .B1(new_n779), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT52), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(KEYINPUT52), .A2(new_n790), .A3(new_n716), .A4(new_n881), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n877), .B(KEYINPUT53), .C1(new_n882), .C2(new_n883), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n884), .A2(KEYINPUT114), .A3(new_n885), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(new_n892), .A3(new_n888), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n756), .A2(new_n800), .A3(new_n634), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n848), .A2(new_n849), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n784), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n821), .B1(new_n384), .B2(new_n670), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n680), .A2(new_n817), .A3(new_n670), .A4(new_n824), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n447), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n851), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT50), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n760), .A2(new_n730), .A3(new_n188), .A4(new_n758), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n903), .B1(new_n904), .B2(new_n900), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n900), .A3(new_n903), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT115), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n760), .A2(new_n758), .A3(new_n842), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n447), .B1(new_n898), .B2(new_n899), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n773), .A2(new_n788), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n652), .A2(new_n723), .A3(new_n447), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n385), .A2(new_n670), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  OR3_X1    g732(.A1(new_n904), .A2(new_n900), .A3(new_n903), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT115), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n905), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n902), .A2(new_n908), .A3(new_n918), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n900), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n771), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n671), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n446), .B1(new_n915), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT48), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n911), .B2(new_n794), .ZN(new_n930));
  NOR4_X1   g744(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT48), .A4(new_n793), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n926), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT116), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n702), .B1(new_n823), .B2(new_n825), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n935), .A2(new_n758), .A3(new_n760), .A4(new_n842), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT48), .B1(new_n936), .B2(new_n793), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n911), .A2(new_n929), .A3(new_n794), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(KEYINPUT116), .A3(new_n926), .A4(new_n928), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n913), .A2(new_n917), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n896), .B2(new_n901), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n923), .B1(new_n919), .B2(new_n905), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND4_X1   g759(.A1(new_n894), .A2(new_n924), .A3(new_n941), .A4(new_n945), .ZN(new_n946));
  AOI22_X1  g760(.A1(new_n934), .A2(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n894), .B1(new_n947), .B2(new_n924), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n891), .A2(new_n893), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(G952), .A2(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n756), .A2(new_n634), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT49), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n730), .A2(new_n723), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n780), .A2(new_n801), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT112), .ZN(new_n957));
  OR4_X1    g771(.A1(new_n818), .A2(new_n954), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT118), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n952), .A2(KEYINPUT118), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G75));
  NOR2_X1   g777(.A1(new_n324), .A2(G952), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n886), .A2(new_n888), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(G902), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT56), .B1(new_n968), .B2(G210), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n253), .B(new_n286), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT55), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n965), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n969), .B2(new_n972), .ZN(G51));
  NAND2_X1  g788(.A1(new_n966), .A2(KEYINPUT54), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(KEYINPUT119), .A3(new_n893), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT119), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n966), .A2(new_n977), .A3(KEYINPUT54), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n635), .B(KEYINPUT57), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n632), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n837), .B(KEYINPUT120), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n968), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n964), .B1(new_n981), .B2(new_n983), .ZN(G54));
  NAND2_X1  g798(.A1(new_n370), .A2(new_n371), .ZN(new_n985));
  NAND2_X1  g799(.A1(KEYINPUT58), .A2(G475), .ZN(new_n986));
  OR3_X1    g800(.A1(new_n967), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n967), .B2(new_n986), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n965), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT121), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT121), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n987), .A2(new_n991), .A3(new_n965), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(G60));
  NAND3_X1  g807(.A1(new_n659), .A2(new_n663), .A3(new_n665), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  XOR2_X1   g809(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n996));
  NOR2_X1   g810(.A1(new_n386), .A2(new_n307), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  AND4_X1   g812(.A1(new_n995), .A2(new_n976), .A3(new_n978), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n891), .A2(new_n893), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n995), .B1(new_n1000), .B2(new_n998), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n999), .A2(new_n1001), .A3(new_n964), .ZN(G63));
  INV_X1    g816(.A(KEYINPUT124), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n965), .B1(new_n1003), .B2(KEYINPUT61), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G217), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT60), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n966), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1004), .B1(new_n1007), .B2(new_n485), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n966), .A2(new_n693), .A3(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(KEYINPUT123), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT123), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n966), .A2(new_n1011), .A3(new_n693), .A4(new_n1006), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1003), .A2(KEYINPUT61), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(G66));
  OAI21_X1  g829(.A(G953), .B1(new_n449), .B2(new_n254), .ZN(new_n1016));
  INV_X1    g830(.A(new_n869), .ZN(new_n1017));
  INV_X1    g831(.A(new_n324), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n250), .B(new_n252), .C1(G898), .C2(new_n324), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT125), .Z(new_n1021));
  XNOR2_X1  g835(.A(new_n1019), .B(new_n1021), .ZN(G69));
  NOR2_X1   g836(.A1(new_n550), .A2(new_n551), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(new_n363), .Z(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n878), .A2(new_n748), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n738), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT62), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n738), .A2(new_n1029), .A3(new_n1026), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n735), .B1(new_n671), .B2(new_n860), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1031), .A2(new_n575), .A3(new_n842), .ZN(new_n1032));
  AND3_X1   g846(.A1(new_n843), .A2(new_n853), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1028), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1025), .B1(new_n1034), .B2(new_n324), .ZN(new_n1035));
  INV_X1    g849(.A(G900), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1025), .B1(new_n1036), .B2(new_n324), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n843), .A2(new_n1026), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n840), .A2(new_n779), .A3(new_n794), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n853), .A2(new_n809), .A3(new_n811), .A4(new_n1039), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1037), .B1(new_n1041), .B2(new_n324), .ZN(new_n1042));
  AND2_X1   g856(.A1(new_n1025), .A2(KEYINPUT126), .ZN(new_n1043));
  AOI211_X1 g857(.A(new_n324), .B(new_n1043), .C1(G227), .C2(G900), .ZN(new_n1044));
  OR3_X1    g858(.A1(new_n1035), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1044), .B1(new_n1035), .B2(new_n1042), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1045), .A2(new_n1046), .ZN(G72));
  NAND2_X1  g861(.A1(G472), .A2(G902), .ZN(new_n1048));
  XOR2_X1   g862(.A(new_n1048), .B(KEYINPUT63), .Z(new_n1049));
  INV_X1    g863(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1050), .B1(new_n543), .B2(new_n554), .ZN(new_n1051));
  AND3_X1   g865(.A1(new_n889), .A2(new_n890), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1050), .B1(new_n1041), .B2(new_n1017), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n718), .A2(new_n503), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n965), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1049), .B1(new_n1034), .B2(new_n869), .ZN(new_n1056));
  AOI211_X1 g870(.A(new_n1052), .B(new_n1055), .C1(new_n1056), .C2(new_n719), .ZN(G57));
endmodule


