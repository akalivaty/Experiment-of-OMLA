

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X2 U323 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n318) );
  XNOR2_X1 U324 ( .A(n480), .B(KEYINPUT125), .ZN(n585) );
  XOR2_X1 U325 ( .A(n306), .B(n305), .Z(n514) );
  XOR2_X1 U326 ( .A(KEYINPUT94), .B(n372), .Z(n512) );
  NOR2_X1 U327 ( .A1(n570), .A2(n569), .ZN(n291) );
  XOR2_X1 U328 ( .A(KEYINPUT45), .B(n464), .Z(n292) );
  XNOR2_X1 U329 ( .A(n386), .B(G218GAT), .ZN(n387) );
  XNOR2_X1 U330 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U331 ( .A(n423), .B(n300), .ZN(n301) );
  XNOR2_X1 U332 ( .A(n347), .B(n301), .ZN(n302) );
  NOR2_X1 U333 ( .A1(n478), .A2(n512), .ZN(n554) );
  INV_X1 U334 ( .A(KEYINPUT102), .ZN(n418) );
  INV_X1 U335 ( .A(G218GAT), .ZN(n481) );
  INV_X1 U336 ( .A(G78GAT), .ZN(n460) );
  INV_X1 U337 ( .A(G15GAT), .ZN(n454) );
  XNOR2_X1 U338 ( .A(n481), .B(KEYINPUT62), .ZN(n482) );
  XNOR2_X1 U339 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U340 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U341 ( .A(n483), .B(n482), .ZN(G1355GAT) );
  XNOR2_X1 U342 ( .A(n463), .B(n462), .ZN(G1335GAT) );
  XOR2_X1 U343 ( .A(G183GAT), .B(KEYINPUT19), .Z(n294) );
  XNOR2_X1 U344 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n341) );
  XOR2_X1 U346 ( .A(G64GAT), .B(G92GAT), .Z(n296) );
  XNOR2_X1 U347 ( .A(G176GAT), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n441) );
  XNOR2_X1 U349 ( .A(n341), .B(n441), .ZN(n306) );
  XOR2_X1 U350 ( .A(G36GAT), .B(G190GAT), .Z(n379) );
  XOR2_X1 U351 ( .A(KEYINPUT21), .B(G218GAT), .Z(n298) );
  XNOR2_X1 U352 ( .A(KEYINPUT90), .B(G211GAT), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U354 ( .A(n299), .B(G197GAT), .Z(n347) );
  XOR2_X1 U355 ( .A(G169GAT), .B(G8GAT), .Z(n423) );
  XOR2_X1 U356 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n300) );
  XOR2_X1 U357 ( .A(n379), .B(n302), .Z(n304) );
  NAND2_X1 U358 ( .A1(G226GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U360 ( .A(n514), .B(KEYINPUT97), .Z(n307) );
  XNOR2_X1 U361 ( .A(n307), .B(KEYINPUT27), .ZN(n366) );
  XOR2_X1 U362 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n309) );
  XNOR2_X1 U363 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U365 ( .A(G1GAT), .B(G127GAT), .Z(n407) );
  XOR2_X1 U366 ( .A(G85GAT), .B(n407), .Z(n311) );
  XOR2_X1 U367 ( .A(G120GAT), .B(G57GAT), .Z(n442) );
  XNOR2_X1 U368 ( .A(G148GAT), .B(n442), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U370 ( .A(n313), .B(n312), .Z(n315) );
  NAND2_X1 U371 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n317) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(G134GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n316), .B(KEYINPUT77), .ZN(n393) );
  XOR2_X1 U375 ( .A(n317), .B(n393), .Z(n324) );
  XNOR2_X1 U376 ( .A(n318), .B(KEYINPUT82), .ZN(n334) );
  XNOR2_X1 U377 ( .A(G155GAT), .B(KEYINPUT91), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n319), .B(KEYINPUT3), .ZN(n320) );
  XOR2_X1 U379 ( .A(n320), .B(KEYINPUT2), .Z(n322) );
  XNOR2_X1 U380 ( .A(G141GAT), .B(G162GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n346) );
  XNOR2_X1 U382 ( .A(n334), .B(n346), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n372) );
  NAND2_X1 U384 ( .A1(n366), .A2(n512), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n325), .B(KEYINPUT98), .ZN(n522) );
  XOR2_X1 U386 ( .A(G176GAT), .B(KEYINPUT87), .Z(n327) );
  XNOR2_X1 U387 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n345) );
  XOR2_X1 U389 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n329) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U392 ( .A(KEYINPUT83), .B(G71GAT), .Z(n331) );
  XNOR2_X1 U393 ( .A(G169GAT), .B(G120GAT), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U395 ( .A(n333), .B(n332), .Z(n339) );
  XOR2_X1 U396 ( .A(n334), .B(G99GAT), .Z(n336) );
  NAND2_X1 U397 ( .A1(G227GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U399 ( .A(G134GAT), .B(n337), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U401 ( .A(n340), .B(G127GAT), .Z(n343) );
  XNOR2_X1 U402 ( .A(G15GAT), .B(n341), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X2 U404 ( .A(n345), .B(n344), .Z(n568) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U406 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n349) );
  XNOR2_X1 U407 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U409 ( .A(KEYINPUT88), .B(n350), .Z(n352) );
  NAND2_X1 U410 ( .A1(G228GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U412 ( .A(n353), .B(KEYINPUT89), .Z(n360) );
  XOR2_X1 U413 ( .A(G78GAT), .B(G148GAT), .Z(n355) );
  XNOR2_X1 U414 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n443) );
  XOR2_X1 U416 ( .A(n443), .B(KEYINPUT24), .Z(n357) );
  XOR2_X1 U417 ( .A(G50GAT), .B(KEYINPUT74), .Z(n380) );
  XNOR2_X1 U418 ( .A(n380), .B(KEYINPUT93), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U420 ( .A(G22GAT), .B(n358), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n555) );
  XOR2_X1 U423 ( .A(n555), .B(KEYINPUT28), .Z(n525) );
  OR2_X1 U424 ( .A1(n568), .A2(n525), .ZN(n363) );
  NOR2_X1 U425 ( .A1(n522), .A2(n363), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n364), .B(KEYINPUT99), .ZN(n375) );
  NOR2_X1 U427 ( .A1(n555), .A2(n568), .ZN(n365) );
  XOR2_X1 U428 ( .A(n365), .B(KEYINPUT26), .Z(n541) );
  INV_X1 U429 ( .A(n541), .ZN(n479) );
  NAND2_X1 U430 ( .A1(n479), .A2(n366), .ZN(n371) );
  AND2_X1 U431 ( .A1(n514), .A2(n568), .ZN(n367) );
  XOR2_X1 U432 ( .A(KEYINPUT100), .B(n367), .Z(n368) );
  NAND2_X1 U433 ( .A1(n555), .A2(n368), .ZN(n369) );
  XOR2_X1 U434 ( .A(KEYINPUT25), .B(n369), .Z(n370) );
  NAND2_X1 U435 ( .A1(n371), .A2(n370), .ZN(n373) );
  NAND2_X1 U436 ( .A1(n373), .A2(n372), .ZN(n374) );
  NAND2_X1 U437 ( .A1(n375), .A2(n374), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n376), .B(KEYINPUT101), .ZN(n491) );
  XOR2_X1 U439 ( .A(KEYINPUT75), .B(KEYINPUT9), .Z(n378) );
  XNOR2_X1 U440 ( .A(G162GAT), .B(KEYINPUT76), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n397) );
  XOR2_X1 U442 ( .A(n379), .B(G92GAT), .Z(n382) );
  XNOR2_X1 U443 ( .A(n380), .B(G106GAT), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U445 ( .A(n383), .B(KEYINPUT10), .Z(n390) );
  XOR2_X1 U446 ( .A(G99GAT), .B(G85GAT), .Z(n449) );
  XOR2_X1 U447 ( .A(G43GAT), .B(KEYINPUT7), .Z(n385) );
  XNOR2_X1 U448 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n427) );
  XOR2_X1 U450 ( .A(n449), .B(n427), .Z(n388) );
  NAND2_X1 U451 ( .A1(G232GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n392) );
  INV_X1 U453 ( .A(KEYINPUT65), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n393), .B(KEYINPUT11), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X2 U457 ( .A(n397), .B(n396), .Z(n570) );
  XOR2_X1 U458 ( .A(KEYINPUT78), .B(KEYINPUT81), .Z(n399) );
  NAND2_X1 U459 ( .A1(G231GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U461 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n401) );
  XNOR2_X1 U462 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U464 ( .A(n403), .B(n402), .Z(n409) );
  XOR2_X1 U465 ( .A(KEYINPUT79), .B(G64GAT), .Z(n405) );
  XNOR2_X1 U466 ( .A(G8GAT), .B(G57GAT), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U470 ( .A(G78GAT), .B(G155GAT), .Z(n411) );
  XNOR2_X1 U471 ( .A(G183GAT), .B(G211GAT), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U473 ( .A(n413), .B(n412), .Z(n415) );
  XOR2_X1 U474 ( .A(G15GAT), .B(G22GAT), .Z(n426) );
  XOR2_X1 U475 ( .A(G71GAT), .B(KEYINPUT13), .Z(n440) );
  XNOR2_X1 U476 ( .A(n426), .B(n440), .ZN(n414) );
  XOR2_X1 U477 ( .A(n415), .B(n414), .Z(n565) );
  INV_X1 U478 ( .A(n565), .ZN(n584) );
  NAND2_X1 U479 ( .A1(n570), .A2(n584), .ZN(n416) );
  XNOR2_X1 U480 ( .A(KEYINPUT16), .B(n416), .ZN(n417) );
  NOR2_X1 U481 ( .A1(n491), .A2(n417), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n459) );
  XOR2_X1 U483 ( .A(G141GAT), .B(G197GAT), .Z(n421) );
  XNOR2_X1 U484 ( .A(G50GAT), .B(G113GAT), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U486 ( .A(n422), .B(G36GAT), .Z(n425) );
  XNOR2_X1 U487 ( .A(n423), .B(G29GAT), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U489 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U490 ( .A1(G229GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U492 ( .A(n431), .B(n430), .Z(n439) );
  XOR2_X1 U493 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n433) );
  XNOR2_X1 U494 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U496 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n435) );
  XNOR2_X1 U497 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U500 ( .A(n439), .B(n438), .Z(n542) );
  INV_X1 U501 ( .A(n542), .ZN(n578) );
  XOR2_X1 U502 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n447) );
  XNOR2_X1 U506 ( .A(KEYINPUT31), .B(KEYINPUT72), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U508 ( .A(n449), .B(n448), .Z(n451) );
  NAND2_X1 U509 ( .A1(G230GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U511 ( .A(n453), .B(n452), .Z(n581) );
  OR2_X1 U512 ( .A1(n578), .A2(n581), .ZN(n493) );
  NOR2_X1 U513 ( .A1(n459), .A2(n493), .ZN(n487) );
  NAND2_X1 U514 ( .A1(n487), .A2(n568), .ZN(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n455) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(G1326GAT) );
  XNOR2_X1 U517 ( .A(n581), .B(KEYINPUT41), .ZN(n544) );
  XNOR2_X1 U518 ( .A(KEYINPUT106), .B(n544), .ZN(n559) );
  NOR2_X1 U519 ( .A1(n559), .A2(n542), .ZN(n458) );
  XNOR2_X1 U520 ( .A(KEYINPUT107), .B(n458), .ZN(n510) );
  NOR2_X1 U521 ( .A1(n459), .A2(n510), .ZN(n508) );
  NAND2_X1 U522 ( .A1(n508), .A2(n525), .ZN(n463) );
  XOR2_X1 U523 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n461) );
  XNOR2_X1 U524 ( .A(KEYINPUT36), .B(n570), .ZN(n489) );
  NOR2_X1 U525 ( .A1(n489), .A2(n565), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n581), .A2(n292), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n465), .A2(n578), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n578), .A2(n544), .ZN(n466) );
  XOR2_X1 U529 ( .A(KEYINPUT112), .B(n466), .Z(n467) );
  XNOR2_X1 U530 ( .A(KEYINPUT46), .B(n467), .ZN(n468) );
  NAND2_X1 U531 ( .A1(n468), .A2(n570), .ZN(n469) );
  NOR2_X1 U532 ( .A1(n584), .A2(n469), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n470), .B(KEYINPUT47), .ZN(n471) );
  NAND2_X1 U534 ( .A1(n472), .A2(n471), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(n523) );
  INV_X1 U537 ( .A(n514), .ZN(n475) );
  NOR2_X1 U538 ( .A1(n523), .A2(n475), .ZN(n477) );
  INV_X1 U539 ( .A(KEYINPUT54), .ZN(n476) );
  XNOR2_X1 U540 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U541 ( .A1(n554), .A2(n479), .ZN(n480) );
  INV_X1 U542 ( .A(n585), .ZN(n577) );
  NOR2_X1 U543 ( .A1(n489), .A2(n577), .ZN(n483) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n512), .A2(n487), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n514), .A2(n487), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(G8GAT), .ZN(G1325GAT) );
  NAND2_X1 U549 ( .A1(n487), .A2(n525), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  OR2_X1 U551 ( .A1(n489), .A2(n584), .ZN(n490) );
  NOR2_X1 U552 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT37), .ZN(n511) );
  NOR2_X1 U554 ( .A1(n511), .A2(n493), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(KEYINPUT38), .ZN(n502) );
  NAND2_X1 U556 ( .A1(n512), .A2(n502), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT39), .B(KEYINPUT104), .Z(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U560 ( .A1(n514), .A2(n502), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n568), .A2(n502), .ZN(n500) );
  XOR2_X1 U563 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(G43GAT), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n525), .A2(n502), .ZN(n503) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n503), .ZN(G1331GAT) );
  NAND2_X1 U568 ( .A1(n512), .A2(n508), .ZN(n504) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n504), .ZN(n505) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n514), .A2(n508), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(KEYINPUT108), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n508), .A2(n568), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  NOR2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n512), .A2(n519), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n519), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  XOR2_X1 U582 ( .A(G99GAT), .B(KEYINPUT111), .Z(n518) );
  NAND2_X1 U583 ( .A1(n519), .A2(n568), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1338GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n525), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(KEYINPUT44), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n529) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(KEYINPUT113), .B(n524), .ZN(n540) );
  NOR2_X1 U591 ( .A1(n525), .A2(n540), .ZN(n526) );
  NAND2_X1 U592 ( .A1(n568), .A2(n526), .ZN(n527) );
  XNOR2_X1 U593 ( .A(KEYINPUT114), .B(n527), .ZN(n536) );
  NOR2_X1 U594 ( .A1(n578), .A2(n536), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n531) );
  NOR2_X1 U597 ( .A1(n559), .A2(n536), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n533) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n536), .A2(n565), .ZN(n534) );
  XOR2_X1 U603 ( .A(n535), .B(n534), .Z(G1342GAT) );
  XNOR2_X1 U604 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n538) );
  NOR2_X1 U605 ( .A1(n570), .A2(n536), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n549), .A2(n542), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  INV_X1 U611 ( .A(n549), .ZN(n551) );
  NOR2_X1 U612 ( .A1(n551), .A2(n544), .ZN(n548) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n549), .A2(n584), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n570), .A2(n551), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT120), .B(n552), .Z(n553) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT55), .B(n556), .ZN(n571) );
  NAND2_X1 U624 ( .A1(n571), .A2(n568), .ZN(n564) );
  NOR2_X1 U625 ( .A1(n578), .A2(n564), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  XNOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n563) );
  NOR2_X1 U629 ( .A1(n559), .A2(n564), .ZN(n561) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n560) );
  XNOR2_X1 U631 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U632 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  INV_X1 U636 ( .A(n568), .ZN(n569) );
  AND2_X1 U637 ( .A1(n571), .A2(n291), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G190GAT), .B(n574), .Z(G1351GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(n580), .B(n579), .Z(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(G1354GAT) );
endmodule

