//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n212), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n230), .B(new_n231), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G41), .ZN(new_n244));
  INV_X1    g0044(.A(G45), .ZN(new_n245));
  AOI21_X1  g0045(.A(G1), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n246), .A2(new_n248), .A3(G274), .ZN(new_n249));
  INV_X1    g0049(.A(G226), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n249), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1698), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n256), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G223), .A3(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n258), .B(new_n260), .C1(new_n261), .C2(new_n259), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n254), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G169), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT67), .ZN(new_n268));
  INV_X1    g0068(.A(G58), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(KEYINPUT8), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(new_n269), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT8), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n268), .B(G58), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n214), .A2(G33), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n267), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n213), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n279), .A2(new_n281), .B1(new_n202), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n281), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n251), .A2(G20), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT68), .B1(new_n283), .B2(new_n281), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G50), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n265), .B(new_n293), .C1(new_n294), .C2(new_n264), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n292), .B(KEYINPUT9), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n264), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G190), .B2(new_n264), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n295), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT7), .B1(new_n307), .B2(new_n214), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT7), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n305), .A2(new_n306), .A3(new_n309), .A4(G20), .ZN(new_n310));
  OAI21_X1  g0110(.A(G68), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(G58), .A2(G68), .ZN(new_n312));
  OAI21_X1  g0112(.A(G20), .B1(new_n312), .B2(new_n201), .ZN(new_n313));
  INV_X1    g0113(.A(G159), .ZN(new_n314));
  NOR4_X1   g0114(.A1(new_n314), .A2(KEYINPUT73), .A3(G20), .A4(G33), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT73), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n266), .B2(G159), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n313), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT74), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT74), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n313), .C1(new_n315), .C2(new_n317), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n311), .A2(new_n319), .A3(KEYINPUT16), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT16), .ZN(new_n323));
  INV_X1    g0123(.A(G68), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n255), .A2(new_n214), .A3(new_n256), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n309), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n256), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n323), .B1(new_n328), .B2(new_n318), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n322), .A2(new_n329), .A3(new_n281), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n282), .B1(new_n272), .B2(new_n276), .ZN(new_n331));
  INV_X1    g0131(.A(new_n277), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n290), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT75), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n330), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n250), .A2(G1698), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n338), .B1(G223), .B2(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G87), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n263), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n248), .A2(G232), .A3(new_n252), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n249), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G169), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n294), .B2(new_n346), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n335), .A2(new_n337), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT18), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n335), .A2(new_n351), .A3(new_n337), .A4(new_n348), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n342), .A2(new_n353), .A3(new_n345), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n248), .B1(new_n339), .B2(new_n340), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n297), .B1(new_n355), .B2(new_n344), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n330), .A2(new_n333), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT17), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n330), .A2(new_n333), .A3(new_n357), .A4(KEYINPUT17), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n350), .A2(new_n352), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n282), .A2(G68), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT12), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n366), .B(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n324), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n261), .B2(new_n278), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT11), .A3(new_n281), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n285), .A2(G68), .A3(new_n288), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT11), .B1(new_n370), .B2(new_n281), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n250), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G232), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G1698), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n378), .B(new_n380), .C1(new_n305), .C2(new_n306), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G97), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n263), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n248), .A2(G238), .A3(new_n252), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n249), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT70), .ZN(new_n389));
  INV_X1    g0189(.A(new_n387), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n248), .B1(new_n381), .B2(new_n382), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n249), .A2(new_n385), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT70), .B(new_n390), .C1(new_n391), .C2(new_n392), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(G169), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n391), .A2(new_n392), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n388), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n396), .A2(KEYINPUT14), .B1(new_n294), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n396), .A2(KEYINPUT14), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n376), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n394), .A2(G200), .A3(new_n395), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT71), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n394), .A2(KEYINPUT71), .A3(G200), .A4(new_n395), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n375), .B1(new_n399), .B2(new_n353), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT72), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT72), .ZN(new_n411));
  AOI211_X1 g0211(.A(new_n411), .B(new_n408), .C1(new_n405), .C2(new_n406), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n402), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(G232), .A2(G1698), .ZN(new_n415));
  INV_X1    g0215(.A(G238), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(G1698), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n307), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n263), .B1(new_n259), .B2(G107), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G244), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n249), .B1(new_n421), .B2(new_n253), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G169), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT8), .B(G58), .ZN(new_n426));
  INV_X1    g0226(.A(new_n266), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n426), .A2(new_n427), .B1(new_n214), .B2(new_n261), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n278), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n281), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n261), .B1(new_n251), .B2(G20), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n285), .A2(new_n432), .B1(new_n261), .B2(new_n283), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n420), .A2(new_n422), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n294), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n425), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n434), .B1(new_n435), .B2(G190), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n423), .A2(G200), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n304), .A2(new_n365), .A3(new_n414), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT77), .ZN(new_n444));
  OAI211_X1 g0244(.A(G250), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT76), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT76), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n259), .A2(new_n447), .A3(G250), .A4(G1698), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(G244), .B(new_n377), .C1(new_n305), .C2(new_n306), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n421), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n257), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n444), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n446), .A2(new_n448), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n257), .A2(new_n453), .B1(G33), .B2(G283), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(KEYINPUT77), .A3(new_n452), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n263), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n251), .A2(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n263), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G257), .ZN(new_n467));
  INV_X1    g0267(.A(G274), .ZN(new_n468));
  AND2_X1   g0268(.A1(G1), .A2(G13), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n247), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G41), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT78), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT78), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n464), .A2(new_n470), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n461), .A2(new_n294), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n283), .A2(new_n205), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n251), .A2(G33), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n282), .A2(new_n480), .A3(new_n213), .A4(new_n280), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(new_n205), .ZN(new_n482));
  XNOR2_X1  g0282(.A(G97), .B(G107), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT6), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n308), .A2(new_n310), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n206), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n482), .B1(new_n490), .B2(new_n281), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n477), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n458), .A2(new_n452), .A3(new_n459), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n248), .B1(new_n494), .B2(new_n444), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(new_n460), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n478), .B(new_n492), .C1(new_n496), .C2(G169), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n461), .A2(G190), .A3(new_n477), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n491), .C1(new_n496), .C2(new_n297), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT23), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n214), .B2(G107), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n214), .B(G87), .C1(new_n305), .C2(new_n306), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT22), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT22), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n259), .A2(new_n509), .A3(new_n214), .A4(G87), .ZN(new_n510));
  AOI211_X1 g0310(.A(KEYINPUT24), .B(new_n506), .C1(new_n508), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n510), .ZN(new_n513));
  INV_X1    g0313(.A(new_n506), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n281), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n481), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n283), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT25), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n282), .B2(G107), .ZN(new_n520));
  AOI22_X1  g0320(.A1(G107), .A2(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n522));
  OAI211_X1 g0322(.A(G250), .B(new_n377), .C1(new_n305), .C2(new_n306), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G294), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n263), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n466), .A2(G264), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(new_n476), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G190), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n263), .A2(new_n525), .B1(new_n466), .B2(G264), .ZN(new_n530));
  AOI21_X1  g0330(.A(G200), .B1(new_n530), .B2(new_n476), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n516), .B(new_n521), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n416), .A2(new_n377), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n421), .A2(G1698), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n305), .C2(new_n306), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT79), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n248), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(KEYINPUT79), .A3(new_n536), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n251), .A2(new_n468), .A3(G45), .ZN(new_n541));
  INV_X1    g0341(.A(G250), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n263), .B1(new_n542), .B2(new_n463), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n294), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n259), .A2(new_n214), .A3(G68), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n214), .B1(new_n382), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G87), .B2(new_n207), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n278), .B2(new_n205), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n281), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n429), .A2(new_n283), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT80), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n481), .B2(new_n429), .ZN(new_n555));
  INV_X1    g0355(.A(new_n429), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n517), .A2(KEYINPUT80), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n552), .A2(new_n553), .A3(new_n555), .A4(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n545), .B(new_n558), .C1(G169), .C2(new_n544), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n544), .A2(G190), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n517), .A2(G87), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n552), .A2(new_n553), .A3(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(new_n562), .C1(new_n297), .C2(new_n544), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n532), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n251), .B(G45), .C1(new_n244), .C2(KEYINPUT5), .ZN(new_n567));
  OAI211_X1 g0367(.A(G270), .B(new_n248), .C1(new_n567), .C2(new_n472), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n476), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G264), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n570));
  OAI211_X1 g0370(.A(G257), .B(new_n377), .C1(new_n305), .C2(new_n306), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n255), .A2(G303), .A3(new_n256), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n248), .B1(new_n573), .B2(KEYINPUT81), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT81), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n570), .A2(new_n571), .A3(new_n575), .A4(new_n572), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n569), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(G116), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n280), .A2(new_n213), .B1(G20), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n455), .B(new_n214), .C1(G33), .C2(new_n205), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(KEYINPUT20), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT20), .B1(new_n579), .B2(new_n580), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n283), .A2(new_n578), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n481), .B2(new_n578), .ZN(new_n585));
  OAI21_X1  g0385(.A(G169), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(KEYINPUT82), .B(new_n566), .C1(new_n577), .C2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT82), .B1(new_n577), .B2(new_n586), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n583), .A2(new_n585), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n294), .B(new_n569), .C1(new_n574), .C2(new_n576), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n588), .A2(KEYINPUT21), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n516), .A2(new_n521), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n530), .A2(KEYINPUT83), .A3(G179), .A4(new_n476), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n528), .A2(G169), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n530), .A2(G179), .A3(new_n476), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT83), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n577), .A2(G190), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(new_n589), .C1(new_n297), .C2(new_n577), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n587), .A2(new_n592), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n443), .A2(new_n500), .A3(new_n565), .A4(new_n602), .ZN(G372));
  NAND2_X1  g0403(.A1(new_n334), .A2(new_n348), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT18), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n334), .A2(new_n351), .A3(new_n348), .ZN(new_n606));
  INV_X1    g0406(.A(new_n402), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n410), .A2(new_n412), .ZN(new_n608));
  INV_X1    g0408(.A(new_n437), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n605), .B(new_n606), .C1(new_n610), .C2(new_n362), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n301), .A2(new_n303), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n295), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT84), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n497), .A2(new_n499), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n564), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n592), .A2(new_n599), .A3(new_n587), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n565), .A2(KEYINPUT84), .A3(new_n497), .A4(new_n499), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n559), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n559), .A2(new_n563), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n461), .A2(new_n477), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n491), .B1(new_n623), .B2(new_n424), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n622), .A2(KEYINPUT26), .A3(new_n478), .A4(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n497), .B2(new_n621), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n620), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n619), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n443), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n613), .A2(new_n630), .ZN(G369));
  NAND2_X1  g0431(.A1(new_n592), .A2(new_n587), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n251), .A2(new_n214), .A3(G13), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n589), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n632), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(G330), .A3(new_n601), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n593), .A2(new_n638), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n599), .A2(new_n532), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n599), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n638), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n638), .B1(new_n592), .B2(new_n587), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n638), .B(KEYINPUT85), .Z(new_n650));
  AOI22_X1  g0450(.A1(new_n645), .A2(new_n649), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT86), .ZN(G399));
  INV_X1    g0453(.A(new_n210), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G1), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n217), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT31), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n537), .A2(new_n538), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n263), .A3(new_n540), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n543), .A2(new_n541), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(new_n294), .A3(new_n528), .ZN(new_n666));
  INV_X1    g0466(.A(new_n577), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n623), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n663), .A2(new_n530), .A3(new_n664), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT87), .B1(new_n544), .B2(new_n530), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT30), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n496), .A4(new_n591), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n530), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n591), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT30), .B1(new_n679), .B2(new_n623), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n669), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n661), .B1(new_n681), .B2(new_n639), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n500), .A2(new_n602), .A3(new_n565), .A4(new_n650), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n677), .A2(new_n591), .A3(new_n678), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n675), .B1(new_n684), .B2(new_n496), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n679), .A2(KEYINPUT30), .A3(new_n623), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n668), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n650), .A2(new_n661), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n682), .A2(new_n683), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT88), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(KEYINPUT88), .A3(G330), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n500), .A2(new_n565), .A3(new_n617), .ZN(new_n697));
  AOI211_X1 g0497(.A(new_n696), .B(new_n638), .C1(new_n628), .C2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT29), .B1(new_n629), .B2(new_n650), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(KEYINPUT89), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT89), .ZN(new_n701));
  INV_X1    g0501(.A(new_n650), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n619), .B2(new_n628), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n703), .B2(KEYINPUT29), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n695), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n660), .B1(new_n705), .B2(G1), .ZN(G364));
  AND2_X1   g0506(.A1(new_n214), .A2(G13), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n251), .B1(new_n707), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n655), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n259), .A2(new_n210), .ZN(new_n711));
  INV_X1    g0511(.A(G355), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n711), .A2(new_n712), .B1(G116), .B2(new_n210), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n307), .A2(new_n210), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT90), .Z(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n217), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n245), .B2(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n239), .A2(new_n245), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n213), .B1(G20), .B2(new_n424), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n710), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n214), .A2(new_n294), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G190), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n259), .B1(new_n731), .B2(G311), .ZN(new_n732));
  INV_X1    g0532(.A(G294), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n353), .A2(G179), .A3(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n214), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n728), .A2(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n353), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT93), .B(G326), .ZN(new_n739));
  OAI221_X1 g0539(.A(new_n732), .B1(new_n733), .B2(new_n735), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NOR4_X1   g0540(.A1(new_n214), .A2(new_n353), .A3(new_n297), .A4(G179), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT94), .Z(new_n742));
  AOI21_X1  g0542(.A(new_n740), .B1(G303), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n736), .A2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(KEYINPUT33), .B(G317), .Z(new_n746));
  NAND3_X1  g0546(.A1(new_n728), .A2(G190), .A3(new_n297), .ZN(new_n747));
  INV_X1    g0547(.A(G322), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n745), .A2(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT95), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n353), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(G179), .B1(new_n751), .B2(KEYINPUT91), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(KEYINPUT91), .B2(new_n751), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n297), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(G200), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G283), .A2(new_n754), .B1(new_n755), .B2(G329), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n743), .A2(new_n750), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n754), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n206), .ZN(new_n759));
  INV_X1    g0559(.A(new_n735), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G97), .A2(new_n760), .B1(new_n744), .B2(G68), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n202), .B2(new_n738), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G77), .A2(new_n731), .B1(new_n741), .B2(G87), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n763), .B(new_n259), .C1(new_n269), .C2(new_n747), .ZN(new_n764));
  OR3_X1    g0564(.A1(new_n759), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n755), .A2(G159), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT92), .B(KEYINPUT32), .Z(new_n767));
  XNOR2_X1  g0567(.A(new_n766), .B(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n757), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n727), .B1(new_n769), .B2(new_n724), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n641), .A2(new_n601), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n723), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n772), .A2(G330), .ZN(new_n775));
  INV_X1    g0575(.A(new_n710), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n642), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(G396));
  NAND2_X1  g0578(.A1(new_n629), .A2(new_n650), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT96), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n437), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n425), .A2(new_n434), .A3(KEYINPUT96), .A4(new_n436), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n438), .A2(new_n439), .B1(new_n434), .B2(new_n638), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n609), .A2(new_n638), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n779), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT97), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n784), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n786), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n703), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g0594(.A1(new_n690), .A2(KEYINPUT88), .A3(G330), .ZN(new_n795));
  AOI21_X1  g0595(.A(KEYINPUT88), .B1(new_n690), .B2(G330), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n710), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n797), .B2(new_n794), .ZN(new_n799));
  INV_X1    g0599(.A(new_n724), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n722), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n710), .B1(G77), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n747), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(G143), .B1(new_n731), .B2(G159), .ZN(new_n804));
  INV_X1    g0604(.A(G150), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n745), .B2(new_n805), .C1(new_n806), .C2(new_n738), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT34), .Z(new_n808));
  OAI21_X1  g0608(.A(new_n259), .B1(new_n735), .B2(new_n269), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n742), .B2(G50), .ZN(new_n810));
  INV_X1    g0610(.A(G132), .ZN(new_n811));
  INV_X1    g0611(.A(new_n755), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n324), .B2(new_n758), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n742), .A2(G107), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n744), .A2(G283), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G97), .A2(new_n760), .B1(new_n737), .B2(G303), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n307), .B1(new_n747), .B2(new_n733), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G116), .B2(new_n731), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n754), .A2(G87), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n812), .B2(new_n821), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n808), .A2(new_n813), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n802), .B1(new_n823), .B2(new_n724), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n792), .B2(new_n722), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n799), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  NOR2_X1   g0627(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n828), .A2(new_n578), .A3(new_n216), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(KEYINPUT98), .B1(KEYINPUT35), .B2(new_n487), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(KEYINPUT98), .B2(new_n830), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT36), .Z(new_n833));
  OAI211_X1 g0633(.A(new_n717), .B(G77), .C1(new_n269), .C2(new_n324), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n202), .A2(G68), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n251), .B(G13), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G330), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT40), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT99), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n355), .A2(new_n344), .A3(new_n294), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G169), .B2(new_n346), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n311), .A2(new_n319), .A3(new_n321), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n323), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n281), .A3(new_n322), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n843), .B1(new_n846), .B2(new_n333), .ZN(new_n847));
  INV_X1    g0647(.A(new_n358), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n841), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n331), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n277), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n322), .A2(new_n281), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n845), .ZN(new_n854));
  OAI211_X1 g0654(.A(KEYINPUT99), .B(new_n358), .C1(new_n854), .C2(new_n843), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n854), .A2(new_n636), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n849), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n358), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n337), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n336), .B1(new_n330), .B2(new_n333), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(new_n862), .B2(new_n348), .ZN(new_n863));
  INV_X1    g0663(.A(new_n636), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n335), .A2(new_n337), .A3(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n857), .A2(KEYINPUT37), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n362), .B1(KEYINPUT18), .B2(new_n349), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n856), .B1(new_n867), .B2(new_n352), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n840), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n854), .A2(new_n636), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n364), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n847), .A2(new_n848), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n872), .B2(KEYINPUT99), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n858), .B1(new_n873), .B2(new_n849), .ZN(new_n874));
  INV_X1    g0674(.A(new_n859), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n349), .A2(new_n865), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT38), .B(new_n871), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n687), .A2(KEYINPUT31), .A3(new_n638), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n682), .A3(new_n683), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n375), .A2(new_n639), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n413), .A2(new_n881), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n402), .B1(new_n375), .B2(new_n639), .C1(new_n410), .C2(new_n412), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n884), .A3(new_n792), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n839), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n880), .A2(new_n884), .A3(new_n792), .ZN(new_n887));
  INV_X1    g0687(.A(new_n865), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n605), .A2(new_n606), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n362), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n604), .A2(new_n358), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n858), .B1(new_n891), .B2(new_n865), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n876), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT100), .B1(new_n893), .B2(new_n840), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n877), .ZN(new_n895));
  INV_X1    g0695(.A(new_n866), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n896), .A2(KEYINPUT100), .A3(KEYINPUT38), .A4(new_n871), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n443), .A2(new_n880), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT101), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n838), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n900), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n402), .A2(new_n638), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n869), .A2(new_n877), .A3(KEYINPUT39), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n895), .A2(new_n897), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n905), .B(new_n906), .C1(new_n907), .C2(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n889), .A2(new_n636), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n781), .A2(new_n782), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n638), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n793), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n869), .A2(new_n877), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n915), .A3(new_n884), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n909), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n779), .A2(KEYINPUT89), .A3(new_n696), .ZN(new_n918));
  INV_X1    g0718(.A(new_n698), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n704), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n613), .B1(new_n920), .B2(new_n442), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n917), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n904), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n251), .B2(new_n707), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n904), .A2(new_n922), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n837), .B1(new_n924), .B2(new_n925), .ZN(G367));
  OAI21_X1  g0726(.A(new_n725), .B1(new_n210), .B2(new_n429), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n715), .B2(new_n235), .ZN(new_n928));
  AOI22_X1  g0728(.A1(G68), .A2(new_n760), .B1(new_n737), .B2(G143), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n314), .B2(new_n745), .ZN(new_n930));
  INV_X1    g0730(.A(new_n741), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n259), .B1(new_n931), .B2(new_n269), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n747), .A2(new_n805), .B1(new_n730), .B2(new_n202), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n934), .B1(new_n261), .B2(new_n758), .C1(new_n806), .C2(new_n812), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n742), .A2(KEYINPUT46), .A3(G116), .ZN(new_n936));
  AOI22_X1  g0736(.A1(G107), .A2(new_n760), .B1(new_n737), .B2(G311), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n741), .A2(G116), .ZN(new_n938));
  XOR2_X1   g0738(.A(KEYINPUT106), .B(KEYINPUT46), .Z(new_n939));
  AOI22_X1  g0739(.A1(new_n938), .A2(new_n939), .B1(new_n744), .B2(G294), .ZN(new_n940));
  INV_X1    g0740(.A(G283), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n307), .B1(new_n730), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G303), .B2(new_n803), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n936), .A2(new_n937), .A3(new_n940), .A4(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(G317), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n205), .A2(new_n758), .B1(new_n812), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n935), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT47), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n776), .B(new_n928), .C1(new_n948), .C2(new_n724), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n562), .A2(new_n639), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n622), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n559), .A2(new_n950), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n723), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT105), .ZN(new_n955));
  INV_X1    g0755(.A(new_n649), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n647), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n645), .A2(new_n649), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(new_n642), .Z(new_n960));
  NAND3_X1  g0760(.A1(new_n705), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT45), .ZN(new_n962));
  INV_X1    g0762(.A(new_n651), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n497), .B(new_n499), .C1(new_n491), .C2(new_n650), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n624), .A2(new_n478), .A3(new_n702), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n962), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n651), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(new_n967), .A3(KEYINPUT44), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n651), .B2(new_n966), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n648), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT104), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n648), .A3(new_n974), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI211_X1 g0778(.A(KEYINPUT104), .B(new_n648), .C1(new_n970), .C2(new_n974), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n920), .A2(new_n960), .A3(new_n797), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT105), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n961), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n705), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n985));
  XNOR2_X1  g0785(.A(new_n655), .B(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n709), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n966), .A2(new_n645), .A3(new_n649), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT42), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n497), .B1(new_n964), .B2(new_n599), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n650), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n951), .A2(new_n952), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT102), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n993), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(KEYINPUT102), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n648), .A2(new_n967), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n997), .A2(new_n1002), .A3(new_n999), .A4(new_n1000), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n954), .B1(new_n987), .B2(new_n1006), .ZN(G387));
  AOI21_X1  g0807(.A(new_n955), .B1(new_n705), .B2(new_n960), .ZN(new_n1008));
  AND4_X1   g0808(.A1(new_n955), .A2(new_n920), .A3(new_n797), .A4(new_n960), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n655), .B1(new_n705), .B2(new_n960), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n647), .A2(new_n723), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n232), .A2(G45), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n426), .A2(G50), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT50), .Z(new_n1014));
  OAI211_X1 g0814(.A(new_n657), .B(new_n245), .C1(new_n324), .C2(new_n261), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1012), .B(new_n715), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(G107), .B2(new_n210), .C1(new_n657), .C2(new_n711), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n776), .B(new_n1011), .C1(new_n725), .C2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n307), .B1(new_n741), .B2(G77), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n758), .B2(new_n205), .C1(new_n805), .C2(new_n812), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT107), .Z(new_n1021));
  AOI22_X1  g0821(.A1(new_n803), .A2(G50), .B1(new_n731), .B2(G68), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n429), .B2(new_n735), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G159), .B2(new_n737), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(new_n277), .C2(new_n745), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n259), .B1(new_n754), .B2(G116), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n803), .A2(G317), .B1(new_n731), .B2(G303), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n745), .B2(new_n821), .C1(new_n748), .C2(new_n738), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n760), .A2(G283), .B1(G294), .B2(new_n741), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT108), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT108), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1026), .B1(new_n739), .B2(new_n812), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1025), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n800), .B1(new_n1039), .B2(KEYINPUT109), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(KEYINPUT109), .B2(new_n1039), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n960), .A2(new_n709), .B1(new_n1018), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1010), .A2(new_n1042), .ZN(G393));
  INV_X1    g0843(.A(new_n975), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n977), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n967), .A2(new_n723), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n725), .B1(new_n205), .B2(new_n210), .C1(new_n716), .C2(new_n242), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n710), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n259), .B1(new_n730), .B2(new_n426), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n745), .A2(new_n202), .B1(new_n261), .B2(new_n735), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(G68), .C2(new_n741), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n738), .A2(new_n805), .B1(new_n314), .B2(new_n747), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n755), .A2(G143), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n820), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT110), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n307), .B1(new_n730), .B2(new_n733), .ZN(new_n1059));
  INV_X1    g0859(.A(G303), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n745), .A2(new_n1060), .B1(new_n578), .B2(new_n735), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1059), .B(new_n1061), .C1(G283), .C2(new_n741), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n759), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n738), .A2(new_n945), .B1(new_n821), .B2(new_n747), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n755), .A2(G322), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1058), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1049), .B1(new_n1069), .B2(new_n724), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1046), .A2(new_n709), .B1(new_n1047), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(KEYINPUT111), .B(new_n1045), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n655), .A3(new_n983), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n961), .A2(new_n982), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT111), .B1(new_n1074), .B2(new_n1045), .ZN(new_n1075));
  OAI211_X1 g0875(.A(KEYINPUT112), .B(new_n1071), .C1(new_n1073), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1045), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT111), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1080), .A2(new_n655), .A3(new_n983), .A4(new_n1072), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT112), .B1(new_n1081), .B2(new_n1071), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n880), .A2(G330), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n884), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n788), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n1087), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n912), .B1(new_n703), .B2(new_n792), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n884), .B1(new_n695), .B2(new_n792), .ZN(new_n1093));
  OAI211_X1 g0893(.A(KEYINPUT113), .B(new_n914), .C1(new_n1093), .C2(new_n1088), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n695), .A2(new_n792), .A3(new_n884), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n638), .B1(new_n628), .B2(new_n697), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n791), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n912), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1087), .B1(new_n1086), .B2(new_n788), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1096), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1095), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n906), .B1(new_n907), .B2(KEYINPUT39), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n905), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n1091), .B2(new_n1087), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n895), .A2(new_n1105), .A3(new_n897), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1099), .A2(new_n1087), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1107), .A2(new_n1111), .A3(new_n1096), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1088), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1086), .A2(new_n442), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n921), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1103), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1107), .A2(new_n1111), .A3(new_n1096), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1104), .A2(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n1113), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1101), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1117), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1118), .A2(new_n655), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT114), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1118), .A2(new_n1124), .A3(KEYINPUT114), .A4(new_n655), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1115), .A2(new_n709), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1104), .A2(new_n721), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n710), .B1(new_n332), .B2(new_n801), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n745), .A2(new_n806), .B1(new_n738), .B2(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n259), .B1(new_n747), .B2(new_n811), .C1(new_n314), .C2(new_n735), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n741), .A2(G150), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT53), .Z(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT115), .Z(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1136), .B(new_n1138), .C1(new_n730), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n755), .A2(G125), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n758), .B2(new_n202), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n742), .A2(G87), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n737), .A2(G283), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G77), .A2(new_n760), .B1(new_n744), .B2(G107), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n307), .B1(new_n730), .B2(new_n205), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G116), .B2(new_n803), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n324), .A2(new_n758), .B1(new_n812), .B2(new_n733), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1142), .A2(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1132), .B1(new_n1152), .B2(new_n724), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1131), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1130), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1129), .A2(new_n1156), .ZN(G378));
  AND3_X1   g0957(.A1(new_n908), .A2(new_n909), .A3(new_n916), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n886), .A2(new_n898), .A3(G330), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n292), .A2(new_n864), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT118), .Z(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n304), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n304), .A2(new_n1164), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1162), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n1161), .A3(new_n1165), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1159), .A2(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n788), .B1(new_n883), .B2(new_n882), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n915), .A2(new_n1174), .A3(new_n880), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n838), .B1(new_n1175), .B2(new_n839), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1173), .B1(new_n1176), .B2(new_n898), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1158), .B1(new_n1172), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1159), .A2(new_n1171), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n898), .A3(new_n1173), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n917), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n708), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1173), .A2(new_n721), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n710), .B1(G50), .B2(new_n801), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n269), .A2(new_n758), .B1(new_n812), .B2(new_n941), .ZN(new_n1185));
  OR3_X1    g0985(.A1(new_n747), .A2(KEYINPUT116), .A3(new_n206), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT116), .B1(new_n747), .B2(new_n206), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n578), .C2(new_n738), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n259), .A2(G41), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n429), .B2(new_n730), .C1(new_n931), .C2(new_n261), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n745), .A2(new_n205), .B1(new_n324), .B2(new_n735), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1185), .A2(new_n1188), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT58), .Z(new_n1193));
  OAI22_X1  g0993(.A1(new_n747), .A2(new_n1133), .B1(new_n730), .B2(new_n806), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G132), .B2(new_n744), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G150), .A2(new_n760), .B1(new_n737), .B2(G125), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n1141), .C2(new_n931), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n755), .A2(G124), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n754), .C2(G159), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1193), .B1(new_n1198), .B2(new_n1202), .C1(new_n1189), .C2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT117), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n800), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1184), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1183), .A2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT119), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1182), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT120), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n917), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT120), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1117), .B1(new_n1122), .B2(new_n1121), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n655), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1211), .B1(new_n1219), .B2(new_n1221), .ZN(G375));
  OAI21_X1  g1022(.A(new_n710), .B1(G68), .B2(new_n801), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n742), .A2(G97), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n744), .A2(G116), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n556), .A2(new_n760), .B1(new_n737), .B2(G294), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n307), .B1(new_n747), .B2(new_n941), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G107), .B2(new_n731), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1228), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n261), .A2(new_n758), .B1(new_n812), .B2(new_n1060), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n742), .A2(G159), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n259), .B1(new_n747), .B2(new_n806), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G150), .B2(new_n731), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G50), .A2(new_n760), .B1(new_n737), .B2(G132), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1140), .A2(new_n744), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n269), .A2(new_n758), .B1(new_n812), .B2(new_n1133), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n1229), .A2(new_n1230), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1223), .B1(new_n1238), .B2(new_n724), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n884), .B2(new_n722), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1122), .B2(new_n708), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT121), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT121), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1240), .C1(new_n1122), .C2(new_n708), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n986), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1245), .A2(new_n1249), .ZN(G381));
  INV_X1    g1050(.A(new_n1211), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT57), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1179), .A2(new_n917), .A3(new_n1180), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT120), .B1(new_n1253), .B2(new_n1214), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1178), .A2(new_n1212), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1252), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n656), .B1(new_n1256), .B2(new_n1217), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1221), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1251), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1125), .A2(new_n1156), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G381), .A2(new_n1260), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(G387), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .A4(new_n1083), .ZN(G407));
  INV_X1    g1063(.A(new_n1260), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1259), .A2(new_n637), .A3(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G407), .A2(G213), .A3(new_n1265), .ZN(G409));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1155), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(G375), .A2(new_n1270), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1217), .A2(new_n986), .A3(new_n1220), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1209), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1273), .B1(new_n1274), .B2(new_n709), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT122), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1272), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n708), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT122), .B1(new_n1278), .B2(new_n1273), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1260), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1269), .B1(new_n1271), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1268), .A2(G2897), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1122), .A2(KEYINPUT60), .A3(new_n1123), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1283), .A2(new_n655), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT60), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1248), .B1(new_n1246), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1287), .A2(new_n1245), .A3(G384), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1287), .B2(new_n1245), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1282), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1245), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n826), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1287), .A2(new_n1245), .A3(G384), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1282), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1281), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G378), .A2(new_n1259), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1272), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n709), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1276), .A3(new_n1209), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1279), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1264), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1269), .A4(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1269), .B(new_n1306), .C1(new_n1271), .C2(new_n1280), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1297), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1310));
  XOR2_X1   g1110(.A(G393), .B(G396), .Z(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n984), .A2(new_n986), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n708), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1315));
  AOI22_X1  g1115(.A1(new_n1314), .A2(new_n1315), .B1(new_n953), .B2(new_n949), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1071), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT112), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(G387), .A3(new_n1076), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1312), .B1(new_n1317), .B2(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1320), .A2(KEYINPUT124), .A3(G387), .A4(new_n1076), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G387), .B1(new_n1320), .B2(new_n1076), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1323), .B1(new_n1324), .B2(KEYINPUT125), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1326), .B(G387), .C1(new_n1320), .C2(new_n1076), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT124), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1311), .B1(new_n1321), .B2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1322), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1310), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT123), .ZN(new_n1333));
  AOI22_X1  g1133(.A1(G378), .A2(new_n1259), .B1(new_n1302), .B2(new_n1264), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1333), .B1(new_n1334), .B2(new_n1268), .ZN(new_n1335));
  OAI211_X1 g1135(.A(KEYINPUT123), .B(new_n1269), .C1(new_n1271), .C2(new_n1280), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1335), .A2(new_n1296), .A3(new_n1336), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1334), .A2(new_n1268), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT63), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT61), .B1(new_n1338), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1317), .A2(new_n1326), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1324), .A2(KEYINPUT125), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1330), .A2(new_n1343), .A3(new_n1344), .A4(new_n1323), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1322), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1308), .A2(new_n1340), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1337), .A2(new_n1342), .A3(new_n1347), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1332), .A2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1260), .B1(new_n1351), .B2(new_n1211), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1306), .B1(new_n1271), .B2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(G375), .A2(new_n1264), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1298), .A2(new_n1339), .A3(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1347), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT127), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1356), .A2(new_n1347), .A3(KEYINPUT127), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT126), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1331), .A2(new_n1361), .A3(new_n1353), .A4(new_n1355), .ZN(new_n1362));
  OAI21_X1  g1162(.A(KEYINPUT126), .B1(new_n1356), .B2(new_n1347), .ZN(new_n1363));
  AOI22_X1  g1163(.A1(new_n1359), .A2(new_n1360), .B1(new_n1362), .B2(new_n1363), .ZN(G402));
endmodule


