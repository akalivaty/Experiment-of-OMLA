//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT64), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G101), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT71), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n465), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n478), .A2(new_n480), .A3(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(G113), .A3(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n478), .A2(new_n480), .A3(G125), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n483), .A3(new_n485), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n477), .B1(new_n489), .B2(new_n492), .ZN(G160));
  INV_X1    g068(.A(new_n476), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n475), .A2(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G124), .ZN(new_n497));
  OR2_X1    g072(.A1(G100), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G162));
  NAND4_X1  g076(.A1(new_n478), .A2(new_n480), .A3(G138), .A4(new_n465), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n475), .A2(KEYINPUT4), .A3(G138), .A4(new_n465), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n478), .A2(new_n480), .A3(G126), .A4(G2105), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n507), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT72), .B1(new_n512), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n511), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(G50), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G166));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT6), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n527), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n539), .A2(new_n541), .A3(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G51), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n527), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n520), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n543), .A2(new_n545), .A3(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  AOI21_X1  g125(.A(new_n518), .B1(new_n513), .B2(new_n516), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n534), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n542), .A2(G52), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n520), .A2(new_n538), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G90), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n520), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(G43), .A2(new_n542), .B1(new_n555), .B2(G81), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n561), .A2(KEYINPUT76), .A3(G651), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND3_X1  g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G188));
  NAND3_X1  g149(.A1(new_n551), .A2(G91), .A3(new_n527), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT78), .Z(new_n576));
  AND2_X1   g151(.A1(KEYINPUT77), .A2(G53), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n539), .A2(new_n541), .A3(G543), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n551), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(G65), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n576), .B(new_n579), .C1(new_n585), .C2(new_n534), .ZN(G299));
  INV_X1    g161(.A(G166), .ZN(G303));
  NAND2_X1  g162(.A1(new_n542), .A2(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n551), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n555), .A2(G87), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G288));
  NAND3_X1  g167(.A1(new_n517), .A2(G61), .A3(new_n519), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  AOI211_X1 g172(.A(new_n597), .B(new_n518), .C1(new_n513), .C2(new_n516), .ZN(new_n598));
  NAND2_X1  g173(.A1(G48), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n527), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n596), .A2(new_n601), .ZN(G305));
  INV_X1    g177(.A(new_n555), .ZN(new_n603));
  XNOR2_X1  g178(.A(KEYINPUT81), .B(G85), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n539), .A2(new_n541), .A3(G543), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT80), .B(G47), .Z(new_n606));
  OAI22_X1  g181(.A1(new_n603), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n551), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n534), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(G54), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n551), .B(KEYINPUT79), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n618), .B2(new_n534), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n555), .A2(G92), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT10), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n612), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n612), .B1(new_n622), .B2(G868), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  INV_X1    g200(.A(G299), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n475), .A2(new_n470), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n494), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n496), .A2(G123), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT84), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT83), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT86), .Z(new_n669));
  INV_X1    g244(.A(new_n666), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n667), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n665), .C2(new_n667), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n670), .A2(new_n664), .A3(new_n667), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n669), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT87), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(KEYINPUT87), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n678), .A2(new_n680), .ZN(new_n691));
  AOI22_X1  g266(.A1(new_n689), .A2(new_n690), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  OR3_X1    g267(.A1(new_n687), .A2(new_n682), .A3(new_n691), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n692), .B(new_n693), .C1(new_n690), .C2(new_n689), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  INV_X1    g272(.A(G1981), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n696), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G23), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n591), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT33), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1976), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G6), .B(G305), .S(G16), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT32), .B(G1981), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n706), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n702), .A2(G24), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n610), .B2(new_n702), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G1986), .Z(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n706), .A2(new_n719), .A3(new_n710), .A4(new_n713), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n494), .A2(KEYINPUT88), .A3(G131), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n722));
  INV_X1    g297(.A(G131), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n476), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n496), .A2(G119), .ZN(new_n725));
  OR2_X1    g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n721), .A2(new_n724), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT89), .ZN(new_n729));
  MUX2_X1   g304(.A(G25), .B(new_n729), .S(G29), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT35), .B(G1991), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n730), .B(new_n731), .Z(new_n732));
  NAND4_X1  g307(.A1(new_n715), .A2(new_n718), .A3(new_n720), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(KEYINPUT36), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT91), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(KEYINPUT36), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT90), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n470), .A2(G103), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n494), .A2(G139), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n739), .B(new_n740), .C1(new_n465), .C2(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G33), .B(new_n742), .S(G29), .Z(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G2072), .Z(new_n744));
  OR2_X1    g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G160), .B2(new_n746), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G2084), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n494), .A2(G141), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n496), .A2(G129), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n470), .A2(G105), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT26), .Z(new_n755));
  NAND4_X1  g330(.A1(new_n751), .A2(new_n752), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G29), .B2(G32), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n744), .A2(new_n750), .A3(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT95), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n643), .A2(new_n746), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n762), .B2(KEYINPUT95), .ZN(new_n765));
  NOR2_X1   g340(.A1(G4), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n622), .B2(G16), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT92), .B(G1348), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(G11), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n772));
  INV_X1    g347(.A(G26), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G29), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G140), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n476), .A2(KEYINPUT94), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(KEYINPUT94), .B1(new_n476), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n496), .A2(G128), .ZN(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(G29), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n772), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n771), .B1(new_n784), .B2(G2067), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G2067), .B2(new_n784), .ZN(new_n786));
  INV_X1    g361(.A(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(KEYINPUT97), .B1(new_n787), .B2(G29), .ZN(new_n788));
  OR3_X1    g363(.A1(new_n787), .A2(KEYINPUT97), .A3(G29), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n788), .B(new_n789), .C1(G164), .C2(new_n746), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT30), .B(G28), .Z(new_n793));
  OAI221_X1 g368(.A(new_n792), .B1(G29), .B2(new_n793), .C1(new_n759), .C2(new_n760), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G1961), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n786), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n763), .A2(new_n765), .A3(new_n769), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n770), .B2(G11), .ZN(new_n800));
  NOR2_X1   g375(.A1(G29), .A2(G35), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G162), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT29), .ZN(new_n803));
  INV_X1    g378(.A(G2090), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n807));
  INV_X1    g382(.A(G20), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G16), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n806), .B(new_n809), .C1(new_n626), .C2(new_n702), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1956), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n702), .A2(G21), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G168), .B2(new_n702), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n796), .A2(G1961), .B1(G1966), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G1966), .B2(new_n813), .ZN(new_n815));
  INV_X1    g390(.A(G19), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT93), .B1(new_n816), .B2(G16), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n816), .A2(KEYINPUT93), .A3(G16), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n817), .B(new_n818), .C1(new_n567), .C2(new_n702), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1341), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n749), .A2(G2084), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT96), .Z(new_n822));
  NOR4_X1   g397(.A1(new_n811), .A2(new_n815), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n800), .A2(new_n805), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n735), .A2(new_n737), .B1(new_n826), .B2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n735), .A2(new_n737), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(G150));
  NAND2_X1  g406(.A1(new_n555), .A2(G93), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n605), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n551), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n534), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT100), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT99), .B(KEYINPUT37), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n622), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n837), .A2(new_n567), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n834), .A2(new_n836), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT39), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n843), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n841), .B1(new_n850), .B2(G860), .ZN(G145));
  XOR2_X1   g426(.A(new_n500), .B(KEYINPUT101), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n643), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G160), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n742), .B(new_n756), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n729), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n509), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n508), .A2(new_n506), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n860), .A2(KEYINPUT102), .A3(new_n504), .A4(new_n505), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n863), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n864));
  INV_X1    g439(.A(G142), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n476), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G130), .B2(new_n496), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n862), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n636), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n782), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n857), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n857), .A2(new_n870), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g450(.A(G166), .B(G305), .ZN(new_n876));
  XNOR2_X1  g451(.A(G288), .B(new_n610), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n631), .B(new_n848), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n620), .B(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(new_n616), .C1(new_n534), .C2(new_n618), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n626), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n622), .A2(G299), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT41), .B1(new_n885), .B2(new_n886), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n881), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n885), .A2(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(new_n881), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n880), .B(new_n893), .ZN(new_n894));
  MUX2_X1   g469(.A(new_n837), .B(new_n894), .S(G868), .Z(G295));
  MUX2_X1   g470(.A(new_n837), .B(new_n894), .S(G868), .Z(G331));
  XNOR2_X1  g471(.A(G168), .B(G301), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n848), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n889), .B2(new_n890), .ZN(new_n899));
  XNOR2_X1  g474(.A(G301), .B(G286), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n848), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n887), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n899), .A2(new_n878), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n878), .B1(new_n899), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n872), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n907));
  INV_X1    g482(.A(new_n878), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n909));
  INV_X1    g484(.A(new_n890), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n901), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n898), .A2(new_n892), .ZN(new_n912));
  OAI211_X1 g487(.A(KEYINPUT104), .B(new_n908), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n899), .B(new_n902), .C1(new_n914), .C2(new_n878), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n872), .A3(new_n915), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n907), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n905), .A2(new_n918), .A3(new_n919), .A4(new_n872), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n899), .A2(new_n878), .A3(new_n902), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n922), .A2(new_n919), .A3(new_n872), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT105), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n920), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n917), .B1(new_n929), .B2(new_n930), .ZN(G397));
  AOI21_X1  g506(.A(G1384), .B1(new_n859), .B2(new_n861), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n494), .A2(G137), .B1(new_n468), .B2(new_n472), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n483), .A2(new_n485), .ZN(new_n934));
  AOI211_X1 g509(.A(new_n488), .B(new_n465), .C1(new_n934), .C2(new_n490), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT70), .B1(new_n491), .B2(G2105), .ZN(new_n936));
  OAI211_X1 g511(.A(G40), .B(new_n933), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  OR3_X1    g512(.A1(new_n932), .A2(KEYINPUT45), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT107), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(G1996), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n757), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n729), .A2(new_n731), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n939), .B(KEYINPUT109), .ZN(new_n945));
  INV_X1    g520(.A(G2067), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n782), .B(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(new_n757), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(new_n944), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G2067), .B2(new_n782), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n945), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n947), .A2(new_n757), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n945), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n940), .A2(KEYINPUT46), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n940), .A2(KEYINPUT46), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n959));
  XNOR2_X1  g534(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n729), .A2(new_n731), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n945), .B1(new_n944), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n939), .ZN(new_n963));
  NOR2_X1   g538(.A1(G290), .A2(G1986), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT48), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n943), .A2(new_n962), .A3(new_n950), .A4(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n953), .A2(new_n960), .A3(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT111), .B(G8), .Z(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n509), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n937), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n596), .A2(new_n601), .A3(new_n698), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n534), .B1(new_n593), .B2(new_n594), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n514), .B1(KEYINPUT5), .B2(new_n515), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n512), .A2(KEYINPUT72), .A3(G543), .ZN(new_n976));
  OAI211_X1 g551(.A(G86), .B(new_n519), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n538), .B1(new_n977), .B2(new_n599), .ZN(new_n978));
  OAI21_X1  g553(.A(G1981), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n973), .A2(KEYINPUT49), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n972), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n698), .B1(new_n596), .B2(new_n601), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n974), .A2(new_n978), .A3(G1981), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT112), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n973), .A2(new_n979), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n982), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n981), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n987), .B2(new_n982), .ZN(new_n993));
  AOI211_X1 g568(.A(KEYINPUT112), .B(KEYINPUT49), .C1(new_n973), .C2(new_n979), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(KEYINPUT113), .A3(new_n981), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n591), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n972), .B1(new_n999), .B2(new_n973), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n1002));
  INV_X1    g577(.A(new_n969), .ZN(new_n1003));
  NOR2_X1   g578(.A1(G168), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n509), .A2(new_n970), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n509), .B2(new_n970), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n937), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G2084), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n971), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(G160), .A3(G40), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1966), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1011), .A2(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1005), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1021));
  INV_X1    g596(.A(new_n937), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1010), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n509), .A2(new_n970), .A3(new_n1007), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1022), .A2(new_n1012), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n969), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1004), .A2(KEYINPUT51), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1020), .A2(KEYINPUT51), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1018), .A2(new_n1005), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1002), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1019), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT51), .B1(new_n1032), .B2(new_n1004), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1028), .B1(new_n1018), .B2(new_n1003), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1030), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(KEYINPUT119), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1001), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n937), .B1(new_n1013), .B2(new_n971), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n932), .A2(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n709), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1011), .A2(new_n804), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(G166), .B2(new_n1019), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n531), .A2(KEYINPUT55), .A3(G8), .A4(new_n532), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n971), .A2(new_n1006), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n509), .A2(new_n1009), .A3(new_n970), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1050), .A2(G160), .A3(G40), .A4(new_n1051), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1052), .A2(G2090), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1003), .B1(new_n1042), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1049), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n588), .A2(new_n590), .A3(G1976), .A4(new_n589), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n969), .C1(new_n937), .C2(new_n971), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n591), .B2(G1976), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1060), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1057), .B1(new_n997), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT115), .B(new_n1063), .C1(new_n992), .C2(new_n996), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1056), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1038), .A2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1041), .B2(G2078), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1071));
  INV_X1    g646(.A(G1961), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1070), .B(new_n1073), .C1(new_n1016), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G171), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT119), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1002), .B(new_n1030), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1079), .B2(new_n1001), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1000), .B1(new_n1068), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT113), .B1(new_n995), .B2(new_n981), .ZN(new_n1082));
  AND4_X1   g657(.A1(KEYINPUT113), .A2(new_n981), .A3(new_n986), .A4(new_n989), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1064), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1049), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n997), .A2(KEYINPUT114), .A3(new_n1064), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1073), .B(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n933), .A2(G40), .A3(new_n487), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1092), .B(new_n1093), .C1(new_n932), .C2(KEYINPUT45), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1094), .A2(new_n1040), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1093), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1074), .B1(new_n1097), .B2(KEYINPUT122), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1070), .B(new_n1091), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G171), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1075), .A2(G171), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1101), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1076), .B1(new_n1101), .B2(G171), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1110), .A2(new_n1106), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n937), .A2(new_n971), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT58), .B(G1341), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1041), .A2(G1996), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n567), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT59), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1117), .A3(new_n567), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G1348), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1071), .A2(new_n1120), .B1(new_n946), .B2(new_n1112), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n884), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n884), .B1(new_n1121), .B2(KEYINPUT60), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n1122), .A2(new_n1123), .B1(KEYINPUT60), .B2(new_n1121), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1039), .A2(new_n1040), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1052), .A2(KEYINPUT118), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT118), .B1(new_n1052), .B2(new_n1127), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n1131));
  NAND2_X1  g706(.A1(G299), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT9), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n578), .B(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n534), .B1(new_n583), .B2(new_n584), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(KEYINPUT57), .A3(new_n576), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1130), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1138), .B(new_n1126), .C1(new_n1129), .C2(new_n1128), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1119), .B(new_n1124), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1142), .A2(new_n622), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1121), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1146), .A2(new_n1147), .B1(new_n1139), .B2(new_n1130), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1067), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1109), .A2(new_n1111), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1081), .A2(new_n1089), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1044), .A2(G8), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1086), .A2(new_n1088), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1086), .A2(KEYINPUT116), .A3(new_n1088), .A4(new_n1155), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1027), .A2(G286), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1049), .A2(KEYINPUT63), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1153), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  AOI211_X1 g739(.A(KEYINPUT117), .B(new_n1162), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1067), .A2(G286), .A3(new_n1027), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1167), .A2(KEYINPUT63), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1152), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n963), .B1(new_n964), .B2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n943), .A2(new_n962), .A3(new_n950), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n968), .B1(new_n1169), .B2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g748(.A1(G227), .A2(new_n463), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n1175), .A2(KEYINPUT126), .ZN(new_n1176));
  AND2_X1   g750(.A1(new_n874), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g751(.A(G229), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n1175), .A2(KEYINPUT126), .ZN(new_n1179));
  AOI21_X1  g753(.A(new_n1179), .B1(new_n660), .B2(new_n662), .ZN(new_n1180));
  NAND4_X1  g754(.A1(new_n1177), .A2(new_n1178), .A3(new_n926), .A4(new_n1180), .ZN(G225));
  INV_X1    g755(.A(G225), .ZN(G308));
endmodule


