

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n766), .A2(n765), .ZN(n769) );
  NOR2_X1 U553 ( .A1(G299), .A2(n642), .ZN(n638) );
  INV_X1 U554 ( .A(KEYINPUT29), .ZN(n646) );
  XNOR2_X1 U555 ( .A(n646), .B(KEYINPUT103), .ZN(n647) );
  AND2_X1 U556 ( .A1(n707), .A2(n596), .ZN(n624) );
  NAND2_X1 U557 ( .A1(n664), .A2(n663), .ZN(n676) );
  XNOR2_X1 U558 ( .A(n534), .B(KEYINPUT65), .ZN(n999) );
  INV_X1 U559 ( .A(KEYINPUT108), .ZN(n767) );
  NOR2_X1 U560 ( .A1(G651), .A2(n579), .ZN(n807) );
  XNOR2_X1 U561 ( .A(n767), .B(KEYINPUT40), .ZN(n768) );
  XNOR2_X1 U562 ( .A(n769), .B(n768), .ZN(G329) );
  NOR2_X1 U563 ( .A1(n545), .A2(n544), .ZN(G160) );
  NOR2_X1 U564 ( .A1(G543), .A2(G651), .ZN(n803) );
  NAND2_X1 U565 ( .A1(G89), .A2(n803), .ZN(n519) );
  XNOR2_X1 U566 ( .A(n519), .B(KEYINPUT72), .ZN(n520) );
  XNOR2_X1 U567 ( .A(n520), .B(KEYINPUT4), .ZN(n522) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n579) );
  INV_X1 U569 ( .A(G651), .ZN(n524) );
  NOR2_X1 U570 ( .A1(n579), .A2(n524), .ZN(n804) );
  NAND2_X1 U571 ( .A1(G76), .A2(n804), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n523), .B(KEYINPUT5), .ZN(n531) );
  NAND2_X1 U574 ( .A1(G51), .A2(n807), .ZN(n528) );
  NOR2_X1 U575 ( .A1(G543), .A2(n524), .ZN(n526) );
  XNOR2_X1 U576 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n525) );
  XNOR2_X1 U577 ( .A(n526), .B(n525), .ZN(n808) );
  NAND2_X1 U578 ( .A1(G63), .A2(n808), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U582 ( .A(n532), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n533), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  NAND2_X1 U586 ( .A1(G113), .A2(n999), .ZN(n537) );
  NOR2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  XOR2_X1 U588 ( .A(KEYINPUT17), .B(n535), .Z(n691) );
  NAND2_X1 U589 ( .A1(G137), .A2(n691), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U591 ( .A(n538), .B(KEYINPUT66), .ZN(n545) );
  INV_X1 U592 ( .A(G2104), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G2105), .A2(n541), .ZN(n553) );
  NAND2_X1 U594 ( .A1(G101), .A2(n553), .ZN(n539) );
  XOR2_X1 U595 ( .A(KEYINPUT23), .B(n539), .Z(n540) );
  XNOR2_X1 U596 ( .A(n540), .B(KEYINPUT64), .ZN(n543) );
  AND2_X1 U597 ( .A1(n541), .A2(G2105), .ZN(n1000) );
  NAND2_X1 U598 ( .A1(G125), .A2(n1000), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U600 ( .A1(G78), .A2(n804), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G65), .A2(n808), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G91), .A2(n803), .ZN(n548) );
  XNOR2_X1 U604 ( .A(KEYINPUT69), .B(n548), .ZN(n549) );
  NOR2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n807), .A2(G53), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(G299) );
  INV_X1 U608 ( .A(n553), .ZN(n554) );
  INV_X1 U609 ( .A(n554), .ZN(n1003) );
  NAND2_X1 U610 ( .A1(G102), .A2(n1003), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G138), .A2(n691), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U613 ( .A1(G114), .A2(n999), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G126), .A2(n1000), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U616 ( .A1(n560), .A2(n559), .ZN(G164) );
  NAND2_X1 U617 ( .A1(G52), .A2(n807), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G64), .A2(n808), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U620 ( .A(KEYINPUT68), .B(n563), .ZN(n568) );
  NAND2_X1 U621 ( .A1(G90), .A2(n803), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G77), .A2(n804), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n566), .Z(n567) );
  NOR2_X1 U625 ( .A1(n568), .A2(n567), .ZN(G171) );
  NAND2_X1 U626 ( .A1(G50), .A2(n807), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G88), .A2(n803), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U629 ( .A1(G75), .A2(n804), .ZN(n571) );
  XNOR2_X1 U630 ( .A(KEYINPUT79), .B(n571), .ZN(n572) );
  NOR2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n808), .A2(G62), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n575), .A2(n574), .ZN(G303) );
  NAND2_X1 U634 ( .A1(G49), .A2(n807), .ZN(n577) );
  NAND2_X1 U635 ( .A1(G74), .A2(G651), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U637 ( .A1(n808), .A2(n578), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n579), .A2(G87), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n581), .A2(n580), .ZN(G288) );
  NAND2_X1 U640 ( .A1(G61), .A2(n808), .ZN(n588) );
  NAND2_X1 U641 ( .A1(G48), .A2(n807), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G86), .A2(n803), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n804), .A2(G73), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT2), .B(n584), .Z(n585) );
  NOR2_X1 U646 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U648 ( .A(n589), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U649 ( .A1(G85), .A2(n803), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G72), .A2(n804), .ZN(n590) );
  NAND2_X1 U651 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U652 ( .A1(G47), .A2(n807), .ZN(n593) );
  NAND2_X1 U653 ( .A1(G60), .A2(n808), .ZN(n592) );
  NAND2_X1 U654 ( .A1(n593), .A2(n592), .ZN(n594) );
  OR2_X1 U655 ( .A1(n595), .A2(n594), .ZN(G290) );
  INV_X1 U656 ( .A(KEYINPUT26), .ZN(n611) );
  NOR2_X1 U657 ( .A1(G164), .A2(G1384), .ZN(n707) );
  NAND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n706) );
  INV_X1 U659 ( .A(n706), .ZN(n596) );
  NAND2_X1 U660 ( .A1(G1996), .A2(n624), .ZN(n597) );
  XOR2_X1 U661 ( .A(n611), .B(n597), .Z(n598) );
  INV_X1 U662 ( .A(n624), .ZN(n666) );
  NAND2_X1 U663 ( .A1(n666), .A2(G1341), .ZN(n610) );
  NAND2_X1 U664 ( .A1(n598), .A2(n610), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n599), .A2(KEYINPUT98), .ZN(n609) );
  NAND2_X1 U666 ( .A1(n803), .A2(G81), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n600), .B(KEYINPUT12), .ZN(n602) );
  NAND2_X1 U668 ( .A1(G68), .A2(n804), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n603), .B(KEYINPUT13), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G43), .A2(n807), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U673 ( .A1(n808), .A2(G56), .ZN(n606) );
  XOR2_X1 U674 ( .A(KEYINPUT14), .B(n606), .Z(n607) );
  NOR2_X1 U675 ( .A1(n608), .A2(n607), .ZN(n967) );
  NAND2_X1 U676 ( .A1(n609), .A2(n967), .ZN(n614) );
  NOR2_X1 U677 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U678 ( .A1(KEYINPUT98), .A2(n612), .ZN(n613) );
  NOR2_X1 U679 ( .A1(n614), .A2(n613), .ZN(n631) );
  NAND2_X1 U680 ( .A1(n803), .A2(G92), .ZN(n621) );
  NAND2_X1 U681 ( .A1(G79), .A2(n804), .ZN(n616) );
  NAND2_X1 U682 ( .A1(G66), .A2(n808), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U684 ( .A1(G54), .A2(n807), .ZN(n617) );
  XNOR2_X1 U685 ( .A(KEYINPUT71), .B(n617), .ZN(n618) );
  NOR2_X1 U686 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U688 ( .A(n622), .B(KEYINPUT15), .ZN(n971) );
  NAND2_X1 U689 ( .A1(n631), .A2(n971), .ZN(n629) );
  NAND2_X1 U690 ( .A1(G1348), .A2(n666), .ZN(n623) );
  XOR2_X1 U691 ( .A(KEYINPUT99), .B(n623), .Z(n627) );
  INV_X1 U692 ( .A(KEYINPUT96), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n625), .B(n624), .ZN(n649) );
  INV_X1 U694 ( .A(n649), .ZN(n634) );
  NAND2_X1 U695 ( .A1(G2067), .A2(n634), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n630), .B(KEYINPUT100), .ZN(n633) );
  OR2_X1 U699 ( .A1(n971), .A2(n631), .ZN(n632) );
  AND2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n640) );
  NAND2_X1 U701 ( .A1(G2072), .A2(n634), .ZN(n635) );
  XOR2_X1 U702 ( .A(KEYINPUT27), .B(n635), .Z(n637) );
  NAND2_X1 U703 ( .A1(n649), .A2(G1956), .ZN(n636) );
  NAND2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n642) );
  XOR2_X1 U705 ( .A(KEYINPUT101), .B(n638), .Z(n639) );
  NOR2_X1 U706 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U707 ( .A(KEYINPUT102), .B(n641), .ZN(n645) );
  NAND2_X1 U708 ( .A1(G299), .A2(n642), .ZN(n643) );
  XOR2_X1 U709 ( .A(n643), .B(KEYINPUT28), .Z(n644) );
  NOR2_X1 U710 ( .A1(n645), .A2(n644), .ZN(n648) );
  XNOR2_X1 U711 ( .A(n648), .B(n647), .ZN(n654) );
  XOR2_X1 U712 ( .A(G2078), .B(KEYINPUT25), .Z(n856) );
  NOR2_X1 U713 ( .A1(n649), .A2(n856), .ZN(n650) );
  XNOR2_X1 U714 ( .A(n650), .B(KEYINPUT97), .ZN(n652) );
  XNOR2_X1 U715 ( .A(G1961), .B(KEYINPUT95), .ZN(n885) );
  NAND2_X1 U716 ( .A1(n885), .A2(n666), .ZN(n651) );
  NAND2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n659) );
  NAND2_X1 U718 ( .A1(G171), .A2(n659), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n664) );
  NAND2_X1 U720 ( .A1(G8), .A2(n666), .ZN(n757) );
  NOR2_X1 U721 ( .A1(G1966), .A2(n757), .ZN(n678) );
  NOR2_X1 U722 ( .A1(G2084), .A2(n666), .ZN(n674) );
  NOR2_X1 U723 ( .A1(n678), .A2(n674), .ZN(n655) );
  XNOR2_X1 U724 ( .A(KEYINPUT104), .B(n655), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n656), .A2(G8), .ZN(n657) );
  XNOR2_X1 U726 ( .A(KEYINPUT30), .B(n657), .ZN(n658) );
  NOR2_X1 U727 ( .A1(G168), .A2(n658), .ZN(n661) );
  NOR2_X1 U728 ( .A1(G171), .A2(n659), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT31), .B(n662), .Z(n663) );
  NAND2_X1 U731 ( .A1(n676), .A2(G286), .ZN(n665) );
  XNOR2_X1 U732 ( .A(KEYINPUT106), .B(n665), .ZN(n671) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n757), .ZN(n668) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n666), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U736 ( .A1(G303), .A2(n669), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n672), .A2(G8), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n673), .B(KEYINPUT32), .ZN(n681) );
  NAND2_X1 U740 ( .A1(G8), .A2(n674), .ZN(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U743 ( .A(KEYINPUT105), .B(n679), .ZN(n680) );
  NAND2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n756) );
  NOR2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NOR2_X1 U746 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n687), .A2(n682), .ZN(n955) );
  INV_X1 U748 ( .A(KEYINPUT33), .ZN(n683) );
  AND2_X1 U749 ( .A1(n955), .A2(n683), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n756), .A2(n684), .ZN(n735) );
  INV_X1 U751 ( .A(n757), .ZN(n685) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n950) );
  AND2_X1 U753 ( .A1(n685), .A2(n950), .ZN(n686) );
  OR2_X1 U754 ( .A1(KEYINPUT33), .A2(n686), .ZN(n690) );
  NAND2_X1 U755 ( .A1(n687), .A2(KEYINPUT33), .ZN(n688) );
  OR2_X1 U756 ( .A1(n757), .A2(n688), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n733) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n942) );
  XOR2_X1 U759 ( .A(G1986), .B(G290), .Z(n952) );
  XOR2_X1 U760 ( .A(G2067), .B(KEYINPUT37), .Z(n741) );
  XNOR2_X1 U761 ( .A(KEYINPUT34), .B(KEYINPUT88), .ZN(n696) );
  NAND2_X1 U762 ( .A1(G104), .A2(n1003), .ZN(n694) );
  INV_X1 U763 ( .A(n691), .ZN(n692) );
  INV_X1 U764 ( .A(n692), .ZN(n1004) );
  NAND2_X1 U765 ( .A1(G140), .A2(n1004), .ZN(n693) );
  NAND2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U767 ( .A(n696), .B(n695), .ZN(n701) );
  NAND2_X1 U768 ( .A1(G116), .A2(n999), .ZN(n698) );
  NAND2_X1 U769 ( .A1(G128), .A2(n1000), .ZN(n697) );
  NAND2_X1 U770 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U771 ( .A(KEYINPUT35), .B(n699), .Z(n700) );
  NOR2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U773 ( .A(n702), .B(KEYINPUT36), .ZN(n703) );
  XNOR2_X1 U774 ( .A(n703), .B(KEYINPUT89), .ZN(n1014) );
  NAND2_X1 U775 ( .A1(n741), .A2(n1014), .ZN(n704) );
  XOR2_X1 U776 ( .A(n704), .B(KEYINPUT90), .Z(n932) );
  INV_X1 U777 ( .A(n932), .ZN(n705) );
  NAND2_X1 U778 ( .A1(n952), .A2(n705), .ZN(n709) );
  NOR2_X1 U779 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U780 ( .A(KEYINPUT87), .B(n708), .ZN(n751) );
  INV_X1 U781 ( .A(n751), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n709), .A2(n729), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n1004), .A2(G141), .ZN(n710) );
  XNOR2_X1 U784 ( .A(n710), .B(KEYINPUT94), .ZN(n717) );
  NAND2_X1 U785 ( .A1(G117), .A2(n999), .ZN(n712) );
  NAND2_X1 U786 ( .A1(G129), .A2(n1000), .ZN(n711) );
  NAND2_X1 U787 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U788 ( .A1(G105), .A2(n1003), .ZN(n713) );
  XOR2_X1 U789 ( .A(KEYINPUT38), .B(n713), .Z(n714) );
  NOR2_X1 U790 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U791 ( .A1(n717), .A2(n716), .ZN(n1020) );
  NAND2_X1 U792 ( .A1(G1996), .A2(n1020), .ZN(n728) );
  NAND2_X1 U793 ( .A1(G107), .A2(n999), .ZN(n718) );
  XNOR2_X1 U794 ( .A(n718), .B(KEYINPUT92), .ZN(n725) );
  NAND2_X1 U795 ( .A1(G95), .A2(n1003), .ZN(n720) );
  NAND2_X1 U796 ( .A1(G131), .A2(n1004), .ZN(n719) );
  NAND2_X1 U797 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U798 ( .A1(G119), .A2(n1000), .ZN(n721) );
  XNOR2_X1 U799 ( .A(KEYINPUT91), .B(n721), .ZN(n722) );
  NOR2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U801 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U802 ( .A(KEYINPUT93), .B(n726), .Z(n1021) );
  NAND2_X1 U803 ( .A1(G1991), .A2(n1021), .ZN(n727) );
  NAND2_X1 U804 ( .A1(n728), .A2(n727), .ZN(n907) );
  NAND2_X1 U805 ( .A1(n729), .A2(n907), .ZN(n742) );
  NAND2_X1 U806 ( .A1(n730), .A2(n742), .ZN(n759) );
  INV_X1 U807 ( .A(n759), .ZN(n731) );
  NAND2_X1 U808 ( .A1(n942), .A2(n731), .ZN(n732) );
  NOR2_X1 U809 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n766) );
  NOR2_X1 U811 ( .A1(G2090), .A2(G303), .ZN(n736) );
  NAND2_X1 U812 ( .A1(G8), .A2(n736), .ZN(n740) );
  NOR2_X1 U813 ( .A1(G1981), .A2(G305), .ZN(n737) );
  XOR2_X1 U814 ( .A(n737), .B(KEYINPUT24), .Z(n738) );
  NOR2_X1 U815 ( .A1(n757), .A2(n738), .ZN(n758) );
  INV_X1 U816 ( .A(n758), .ZN(n739) );
  AND2_X1 U817 ( .A1(n740), .A2(n739), .ZN(n754) );
  NOR2_X1 U818 ( .A1(n1014), .A2(n741), .ZN(n912) );
  NOR2_X1 U819 ( .A1(G1996), .A2(n1020), .ZN(n909) );
  INV_X1 U820 ( .A(n742), .ZN(n745) );
  NOR2_X1 U821 ( .A1(G1986), .A2(G290), .ZN(n743) );
  NOR2_X1 U822 ( .A1(G1991), .A2(n1021), .ZN(n911) );
  NOR2_X1 U823 ( .A1(n743), .A2(n911), .ZN(n744) );
  NOR2_X1 U824 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U825 ( .A1(n909), .A2(n746), .ZN(n747) );
  XOR2_X1 U826 ( .A(KEYINPUT39), .B(n747), .Z(n748) );
  NOR2_X1 U827 ( .A1(n932), .A2(n748), .ZN(n749) );
  NOR2_X1 U828 ( .A1(n912), .A2(n749), .ZN(n750) );
  NOR2_X1 U829 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U830 ( .A(KEYINPUT107), .B(n752), .Z(n762) );
  INV_X1 U831 ( .A(n762), .ZN(n753) );
  AND2_X1 U832 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U833 ( .A1(n756), .A2(n755), .ZN(n764) );
  NOR2_X1 U834 ( .A1(n758), .A2(n757), .ZN(n760) );
  NOR2_X1 U835 ( .A1(n760), .A2(n759), .ZN(n761) );
  OR2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U838 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U839 ( .A(G2443), .B(G2446), .Z(n771) );
  XNOR2_X1 U840 ( .A(G2427), .B(G2451), .ZN(n770) );
  XNOR2_X1 U841 ( .A(n771), .B(n770), .ZN(n777) );
  XOR2_X1 U842 ( .A(G2430), .B(G2454), .Z(n773) );
  XNOR2_X1 U843 ( .A(G1348), .B(G1341), .ZN(n772) );
  XNOR2_X1 U844 ( .A(n773), .B(n772), .ZN(n775) );
  XOR2_X1 U845 ( .A(G2435), .B(G2438), .Z(n774) );
  XNOR2_X1 U846 ( .A(n775), .B(n774), .ZN(n776) );
  XOR2_X1 U847 ( .A(n777), .B(n776), .Z(n778) );
  AND2_X1 U848 ( .A1(G14), .A2(n778), .ZN(G401) );
  AND2_X1 U849 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U850 ( .A1(n1003), .A2(G99), .ZN(n779) );
  XOR2_X1 U851 ( .A(KEYINPUT75), .B(n779), .Z(n781) );
  NAND2_X1 U852 ( .A1(n999), .A2(G111), .ZN(n780) );
  NAND2_X1 U853 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U854 ( .A(KEYINPUT76), .B(n782), .ZN(n785) );
  NAND2_X1 U855 ( .A1(n1000), .A2(G123), .ZN(n783) );
  XOR2_X1 U856 ( .A(KEYINPUT18), .B(n783), .Z(n784) );
  NOR2_X1 U857 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U858 ( .A1(n1004), .A2(G135), .ZN(n786) );
  NAND2_X1 U859 ( .A1(n787), .A2(n786), .ZN(n1019) );
  XNOR2_X1 U860 ( .A(G2096), .B(n1019), .ZN(n788) );
  OR2_X1 U861 ( .A1(G2100), .A2(n788), .ZN(G156) );
  INV_X1 U862 ( .A(G171), .ZN(G301) );
  INV_X1 U863 ( .A(G132), .ZN(G219) );
  INV_X1 U864 ( .A(G57), .ZN(G237) );
  INV_X1 U865 ( .A(G120), .ZN(G236) );
  NAND2_X1 U866 ( .A1(G7), .A2(G661), .ZN(n789) );
  XOR2_X1 U867 ( .A(n789), .B(KEYINPUT10), .Z(n1033) );
  NAND2_X1 U868 ( .A1(n1033), .A2(G567), .ZN(n790) );
  XOR2_X1 U869 ( .A(KEYINPUT11), .B(n790), .Z(G234) );
  NAND2_X1 U870 ( .A1(n967), .A2(G860), .ZN(G153) );
  NAND2_X1 U871 ( .A1(G868), .A2(G301), .ZN(n792) );
  OR2_X1 U872 ( .A1(n971), .A2(G868), .ZN(n791) );
  NAND2_X1 U873 ( .A1(n792), .A2(n791), .ZN(G284) );
  NOR2_X1 U874 ( .A1(G868), .A2(G299), .ZN(n793) );
  XNOR2_X1 U875 ( .A(n793), .B(KEYINPUT74), .ZN(n795) );
  INV_X1 U876 ( .A(G868), .ZN(n821) );
  NOR2_X1 U877 ( .A1(n821), .A2(G286), .ZN(n794) );
  NOR2_X1 U878 ( .A1(n795), .A2(n794), .ZN(G297) );
  INV_X1 U879 ( .A(G860), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n796), .A2(G559), .ZN(n797) );
  NAND2_X1 U881 ( .A1(n797), .A2(n971), .ZN(n798) );
  XNOR2_X1 U882 ( .A(n798), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U883 ( .A1(n971), .A2(G868), .ZN(n799) );
  NOR2_X1 U884 ( .A1(G559), .A2(n799), .ZN(n801) );
  AND2_X1 U885 ( .A1(n821), .A2(n967), .ZN(n800) );
  NOR2_X1 U886 ( .A1(n801), .A2(n800), .ZN(G282) );
  XOR2_X1 U887 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n802) );
  XNOR2_X1 U888 ( .A(G288), .B(n802), .ZN(n814) );
  NAND2_X1 U889 ( .A1(G93), .A2(n803), .ZN(n806) );
  NAND2_X1 U890 ( .A1(G80), .A2(n804), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n812) );
  NAND2_X1 U892 ( .A1(G55), .A2(n807), .ZN(n810) );
  NAND2_X1 U893 ( .A1(G67), .A2(n808), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U895 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U896 ( .A(KEYINPUT77), .B(n813), .Z(n970) );
  XOR2_X1 U897 ( .A(n814), .B(n970), .Z(n816) );
  XOR2_X1 U898 ( .A(n967), .B(G303), .Z(n815) );
  XNOR2_X1 U899 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U900 ( .A(n817), .B(G299), .ZN(n818) );
  XNOR2_X1 U901 ( .A(n818), .B(G290), .ZN(n819) );
  XNOR2_X1 U902 ( .A(G305), .B(n819), .ZN(n974) );
  NAND2_X1 U903 ( .A1(n971), .A2(G559), .ZN(n966) );
  XOR2_X1 U904 ( .A(n974), .B(n966), .Z(n820) );
  NOR2_X1 U905 ( .A1(n821), .A2(n820), .ZN(n823) );
  NOR2_X1 U906 ( .A1(n970), .A2(G868), .ZN(n822) );
  NOR2_X1 U907 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U908 ( .A(KEYINPUT81), .B(n824), .ZN(G295) );
  NAND2_X1 U909 ( .A1(G2078), .A2(G2084), .ZN(n825) );
  XOR2_X1 U910 ( .A(KEYINPUT20), .B(n825), .Z(n826) );
  NAND2_X1 U911 ( .A1(G2090), .A2(n826), .ZN(n828) );
  XNOR2_X1 U912 ( .A(KEYINPUT82), .B(KEYINPUT21), .ZN(n827) );
  XNOR2_X1 U913 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U914 ( .A1(n829), .A2(G2072), .ZN(n830) );
  XOR2_X1 U915 ( .A(KEYINPUT83), .B(n830), .Z(G158) );
  XOR2_X1 U916 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U917 ( .A1(G236), .A2(G237), .ZN(n831) );
  NAND2_X1 U918 ( .A1(G69), .A2(n831), .ZN(n832) );
  XNOR2_X1 U919 ( .A(KEYINPUT85), .B(n832), .ZN(n833) );
  NAND2_X1 U920 ( .A1(n833), .A2(G108), .ZN(n964) );
  NAND2_X1 U921 ( .A1(G567), .A2(n964), .ZN(n834) );
  XOR2_X1 U922 ( .A(KEYINPUT86), .B(n834), .Z(n840) );
  NOR2_X1 U923 ( .A1(G220), .A2(G219), .ZN(n836) );
  XNOR2_X1 U924 ( .A(KEYINPUT84), .B(KEYINPUT22), .ZN(n835) );
  XNOR2_X1 U925 ( .A(n836), .B(n835), .ZN(n837) );
  NAND2_X1 U926 ( .A1(G96), .A2(n837), .ZN(n838) );
  OR2_X1 U927 ( .A1(G218), .A2(n838), .ZN(n965) );
  AND2_X1 U928 ( .A1(n965), .A2(G2106), .ZN(n839) );
  NOR2_X1 U929 ( .A1(n840), .A2(n839), .ZN(G319) );
  INV_X1 U930 ( .A(G319), .ZN(n1026) );
  NAND2_X1 U931 ( .A1(G661), .A2(G483), .ZN(n841) );
  NOR2_X1 U932 ( .A1(n1026), .A2(n841), .ZN(n846) );
  NAND2_X1 U933 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n1033), .ZN(G217) );
  NAND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n843) );
  INV_X1 U936 ( .A(G661), .ZN(n842) );
  NOR2_X1 U937 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U938 ( .A(n844), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n846), .A2(n845), .ZN(G188) );
  NAND2_X1 U942 ( .A1(G124), .A2(n1000), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n847), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U944 ( .A1(G136), .A2(n1004), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n848), .B(KEYINPUT112), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U947 ( .A1(G100), .A2(n1003), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G112), .A2(n999), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U950 ( .A1(n854), .A2(n853), .ZN(G162) );
  XNOR2_X1 U951 ( .A(G2067), .B(KEYINPUT120), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n855), .B(G26), .ZN(n861) );
  XNOR2_X1 U953 ( .A(G1996), .B(G32), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n856), .B(G27), .ZN(n857) );
  NOR2_X1 U955 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U956 ( .A(KEYINPUT121), .B(n859), .ZN(n860) );
  NOR2_X1 U957 ( .A1(n861), .A2(n860), .ZN(n866) );
  XOR2_X1 U958 ( .A(G2072), .B(G33), .Z(n862) );
  NAND2_X1 U959 ( .A1(n862), .A2(G28), .ZN(n864) );
  XNOR2_X1 U960 ( .A(G25), .B(G1991), .ZN(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U962 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U963 ( .A(n867), .B(KEYINPUT53), .ZN(n868) );
  XNOR2_X1 U964 ( .A(KEYINPUT122), .B(n868), .ZN(n874) );
  XOR2_X1 U965 ( .A(G34), .B(KEYINPUT123), .Z(n870) );
  XNOR2_X1 U966 ( .A(G2084), .B(KEYINPUT54), .ZN(n869) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(n872) );
  XNOR2_X1 U968 ( .A(G35), .B(G2090), .ZN(n871) );
  NOR2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U971 ( .A(KEYINPUT55), .B(n875), .Z(n877) );
  INV_X1 U972 ( .A(G29), .ZN(n876) );
  NAND2_X1 U973 ( .A1(n877), .A2(n876), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G11), .A2(n878), .ZN(n904) );
  XNOR2_X1 U975 ( .A(G1986), .B(G24), .ZN(n883) );
  XNOR2_X1 U976 ( .A(G1971), .B(G22), .ZN(n880) );
  XNOR2_X1 U977 ( .A(G1976), .B(G23), .ZN(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U979 ( .A(KEYINPUT125), .B(n881), .ZN(n882) );
  NOR2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U981 ( .A(KEYINPUT58), .B(n884), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n885), .B(G5), .ZN(n886) );
  NAND2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n899) );
  XOR2_X1 U984 ( .A(G1966), .B(G21), .Z(n897) );
  XOR2_X1 U985 ( .A(G19), .B(G1341), .Z(n891) );
  XNOR2_X1 U986 ( .A(G1956), .B(G20), .ZN(n889) );
  XNOR2_X1 U987 ( .A(G1981), .B(G6), .ZN(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n894) );
  XOR2_X1 U990 ( .A(KEYINPUT59), .B(G1348), .Z(n892) );
  XNOR2_X1 U991 ( .A(G4), .B(n892), .ZN(n893) );
  NOR2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n895), .B(KEYINPUT60), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  NOR2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U996 ( .A(KEYINPUT61), .B(n900), .Z(n901) );
  NOR2_X1 U997 ( .A1(G16), .A2(n901), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n902), .B(KEYINPUT126), .ZN(n903) );
  NOR2_X1 U999 ( .A1(n904), .A2(n903), .ZN(n938) );
  XNOR2_X1 U1000 ( .A(G160), .B(G2084), .ZN(n905) );
  NAND2_X1 U1001 ( .A1(n905), .A2(n1019), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n930) );
  XOR2_X1 U1003 ( .A(G2090), .B(G162), .Z(n908) );
  NOR2_X1 U1004 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1005 ( .A(KEYINPUT51), .B(n910), .Z(n914) );
  NOR2_X1 U1006 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(n914), .A2(n913), .ZN(n928) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n1004), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(KEYINPUT116), .ZN(n918) );
  NAND2_X1 U1010 ( .A1(G103), .A2(n1003), .ZN(n916) );
  XOR2_X1 U1011 ( .A(KEYINPUT115), .B(n916), .Z(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n923) );
  NAND2_X1 U1013 ( .A1(G115), .A2(n999), .ZN(n920) );
  NAND2_X1 U1014 ( .A1(G127), .A2(n1000), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1016 ( .A(KEYINPUT47), .B(n921), .Z(n922) );
  NOR2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(n996) );
  XOR2_X1 U1018 ( .A(G2072), .B(n996), .Z(n925) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1021 ( .A(KEYINPUT50), .B(n926), .Z(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(KEYINPUT52), .B(n933), .ZN(n935) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n934) );
  NAND2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1028 ( .A1(n936), .A2(G29), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n962) );
  XOR2_X1 U1030 ( .A(KEYINPUT56), .B(G16), .Z(n960) );
  XOR2_X1 U1031 ( .A(G1961), .B(G301), .Z(n939) );
  XNOR2_X1 U1032 ( .A(n939), .B(KEYINPUT124), .ZN(n948) );
  XNOR2_X1 U1033 ( .A(n967), .B(G1341), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n971), .B(G1348), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n946) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G168), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1038 ( .A(KEYINPUT57), .B(n944), .Z(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n958) );
  NAND2_X1 U1041 ( .A1(G1971), .A2(G303), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1043 ( .A(G1956), .B(G299), .Z(n951) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1045 ( .A1(n954), .A2(n953), .ZN(n956) );
  NAND2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1047 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1048 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1049 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1050 ( .A(n963), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1051 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1052 ( .A(G108), .ZN(G238) );
  NOR2_X1 U1053 ( .A1(n965), .A2(n964), .ZN(G325) );
  INV_X1 U1054 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1055 ( .A(n967), .B(n966), .Z(n968) );
  NOR2_X1 U1056 ( .A1(G860), .A2(n968), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(n970), .B(n969), .ZN(G145) );
  XOR2_X1 U1058 ( .A(KEYINPUT118), .B(G286), .Z(n973) );
  XOR2_X1 U1059 ( .A(n971), .B(G301), .Z(n972) );
  XNOR2_X1 U1060 ( .A(n973), .B(n972), .ZN(n975) );
  XNOR2_X1 U1061 ( .A(n975), .B(n974), .ZN(n976) );
  NOR2_X1 U1062 ( .A1(G37), .A2(n976), .ZN(G397) );
  XOR2_X1 U1063 ( .A(G2100), .B(G2096), .Z(n978) );
  XNOR2_X1 U1064 ( .A(G2090), .B(KEYINPUT43), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(n978), .B(n977), .ZN(n979) );
  XOR2_X1 U1066 ( .A(n979), .B(G2678), .Z(n981) );
  XNOR2_X1 U1067 ( .A(G2072), .B(KEYINPUT110), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(n981), .B(n980), .ZN(n985) );
  XOR2_X1 U1069 ( .A(KEYINPUT42), .B(G2084), .Z(n983) );
  XNOR2_X1 U1070 ( .A(G2067), .B(G2078), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(n983), .B(n982), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(n985), .B(n984), .ZN(G227) );
  XOR2_X1 U1073 ( .A(G1971), .B(G1956), .Z(n987) );
  XNOR2_X1 U1074 ( .A(G1996), .B(G1966), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(n987), .B(n986), .ZN(n991) );
  XOR2_X1 U1076 ( .A(G2474), .B(KEYINPUT111), .Z(n989) );
  XNOR2_X1 U1077 ( .A(G1961), .B(G1981), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(n989), .B(n988), .ZN(n990) );
  XOR2_X1 U1079 ( .A(n991), .B(n990), .Z(n993) );
  XNOR2_X1 U1080 ( .A(G1991), .B(G1976), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n993), .B(n992), .ZN(n995) );
  XOR2_X1 U1082 ( .A(G1986), .B(KEYINPUT41), .Z(n994) );
  XNOR2_X1 U1083 ( .A(n995), .B(n994), .ZN(G229) );
  XOR2_X1 U1084 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n998) );
  XNOR2_X1 U1085 ( .A(n996), .B(KEYINPUT117), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n998), .B(n997), .ZN(n1013) );
  NAND2_X1 U1087 ( .A1(G118), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1088 ( .A1(G130), .A2(n1000), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1011) );
  XNOR2_X1 U1090 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n1009) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(G106), .ZN(n1007) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(G142), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT113), .B(n1005), .Z(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(n1009), .B(n1008), .Z(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(n1013), .B(n1012), .Z(n1016) );
  XNOR2_X1 U1098 ( .A(G164), .B(n1014), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XOR2_X1 U1100 ( .A(G160), .B(n1017), .Z(n1018) );
  XNOR2_X1 U1101 ( .A(n1019), .B(n1018), .ZN(n1024) );
  XNOR2_X1 U1102 ( .A(G162), .B(n1020), .ZN(n1022) );
  XNOR2_X1 U1103 ( .A(n1022), .B(n1021), .ZN(n1023) );
  XNOR2_X1 U1104 ( .A(n1024), .B(n1023), .ZN(n1025) );
  NOR2_X1 U1105 ( .A1(G37), .A2(n1025), .ZN(G395) );
  NOR2_X1 U1106 ( .A1(G401), .A2(n1026), .ZN(n1030) );
  NOR2_X1 U1107 ( .A1(G227), .A2(G229), .ZN(n1027) );
  XNOR2_X1 U1108 ( .A(KEYINPUT49), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1109 ( .A1(G397), .A2(n1028), .ZN(n1029) );
  NAND2_X1 U1110 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1111 ( .A1(n1031), .A2(G395), .ZN(n1032) );
  XOR2_X1 U1112 ( .A(n1032), .B(KEYINPUT119), .Z(G308) );
  INV_X1 U1113 ( .A(G308), .ZN(G225) );
  INV_X1 U1114 ( .A(G96), .ZN(G221) );
  INV_X1 U1115 ( .A(G69), .ZN(G235) );
  INV_X1 U1116 ( .A(n1033), .ZN(G223) );
  INV_X1 U1117 ( .A(G303), .ZN(G166) );
endmodule

