

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U556 ( .A1(n793), .A2(n693), .ZN(n733) );
  BUF_X1 U557 ( .A(n893), .Z(n521) );
  NOR2_X1 U558 ( .A1(G2104), .A2(n551), .ZN(n893) );
  NOR2_X1 U559 ( .A1(n733), .A2(n815), .ZN(n695) );
  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n649) );
  XOR2_X1 U561 ( .A(G543), .B(KEYINPUT0), .Z(n522) );
  XOR2_X1 U562 ( .A(KEYINPUT72), .B(n527), .Z(n523) );
  AND2_X1 U563 ( .A1(n986), .A2(n825), .ZN(n524) );
  AND2_X1 U564 ( .A1(n795), .A2(n823), .ZN(n525) );
  INV_X1 U565 ( .A(KEYINPUT26), .ZN(n694) );
  NOR2_X1 U566 ( .A1(n978), .A2(n698), .ZN(n704) );
  NOR2_X1 U567 ( .A1(n729), .A2(n728), .ZN(n730) );
  AND2_X1 U568 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U569 ( .A1(n758), .A2(n757), .ZN(n766) );
  INV_X1 U570 ( .A(KEYINPUT12), .ZN(n574) );
  NOR2_X1 U571 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U572 ( .A(n575), .B(n574), .ZN(n576) );
  INV_X1 U573 ( .A(KEYINPUT13), .ZN(n579) );
  NOR2_X1 U574 ( .A1(G164), .A2(G1384), .ZN(n793) );
  NOR2_X1 U575 ( .A1(n812), .A2(n524), .ZN(n813) );
  NOR2_X1 U576 ( .A1(n531), .A2(n655), .ZN(n646) );
  XNOR2_X1 U577 ( .A(KEYINPUT5), .B(KEYINPUT73), .ZN(n529) );
  NOR2_X1 U578 ( .A1(G651), .A2(n655), .ZN(n660) );
  XNOR2_X1 U579 ( .A(n530), .B(n529), .ZN(n539) );
  NOR2_X1 U580 ( .A1(n553), .A2(n552), .ZN(n692) );
  XNOR2_X1 U581 ( .A(KEYINPUT7), .B(n540), .ZN(G168) );
  NAND2_X1 U582 ( .A1(n649), .A2(G89), .ZN(n526) );
  XOR2_X1 U583 ( .A(KEYINPUT4), .B(n526), .Z(n528) );
  INV_X1 U584 ( .A(G651), .ZN(n531) );
  XNOR2_X1 U585 ( .A(KEYINPUT66), .B(n522), .ZN(n655) );
  NAND2_X1 U586 ( .A1(n646), .A2(G76), .ZN(n527) );
  NOR2_X1 U587 ( .A1(n528), .A2(n523), .ZN(n530) );
  NOR2_X1 U588 ( .A1(G543), .A2(n531), .ZN(n533) );
  XNOR2_X1 U589 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n532) );
  XNOR2_X1 U590 ( .A(n533), .B(n532), .ZN(n659) );
  NAND2_X1 U591 ( .A1(G63), .A2(n659), .ZN(n535) );
  NAND2_X1 U592 ( .A1(G51), .A2(n660), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n535), .A2(n534), .ZN(n537) );
  XOR2_X1 U594 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n536) );
  XNOR2_X1 U595 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U597 ( .A1(G91), .A2(n649), .ZN(n542) );
  NAND2_X1 U598 ( .A1(G78), .A2(n646), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G65), .A2(n659), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G53), .A2(n660), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(G299) );
  NOR2_X1 U604 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  XOR2_X2 U605 ( .A(KEYINPUT17), .B(n547), .Z(n898) );
  NAND2_X1 U606 ( .A1(G137), .A2(n898), .ZN(n549) );
  INV_X1 U607 ( .A(G2104), .ZN(n554) );
  INV_X1 U608 ( .A(G2105), .ZN(n551) );
  NOR2_X1 U609 ( .A1(n554), .A2(n551), .ZN(n894) );
  NAND2_X1 U610 ( .A1(G113), .A2(n894), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n550), .B(KEYINPUT64), .ZN(n553) );
  AND2_X1 U613 ( .A1(n521), .A2(G125), .ZN(n552) );
  NOR2_X1 U614 ( .A1(G2105), .A2(n554), .ZN(n897) );
  NAND2_X1 U615 ( .A1(G101), .A2(n897), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT23), .B(n555), .Z(n690) );
  AND2_X1 U617 ( .A1(n692), .A2(n690), .ZN(G160) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G57), .ZN(G237) );
  INV_X1 U620 ( .A(G132), .ZN(G219) );
  NAND2_X1 U621 ( .A1(n893), .A2(G126), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT91), .B(n556), .Z(n558) );
  NAND2_X1 U623 ( .A1(n894), .A2(G114), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT92), .B(n559), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G102), .A2(n897), .ZN(n561) );
  NAND2_X1 U627 ( .A1(G138), .A2(n898), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(G164) );
  NAND2_X1 U630 ( .A1(G64), .A2(n659), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G52), .A2(n660), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G90), .A2(n649), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G77), .A2(n646), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(G171) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n830) );
  NAND2_X1 U642 ( .A1(n830), .A2(G567), .ZN(n572) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  NAND2_X1 U644 ( .A1(n659), .A2(G56), .ZN(n573) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n573), .Z(n582) );
  NAND2_X1 U646 ( .A1(G81), .A2(n649), .ZN(n575) );
  XNOR2_X1 U647 ( .A(n576), .B(KEYINPUT69), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G68), .A2(n646), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(n579), .ZN(n581) );
  NOR2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n583), .B(KEYINPUT70), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G43), .A2(n660), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n978) );
  INV_X1 U655 ( .A(G860), .ZN(n599) );
  OR2_X1 U656 ( .A1(n978), .A2(n599), .ZN(n586) );
  XOR2_X1 U657 ( .A(KEYINPUT71), .B(n586), .Z(G153) );
  INV_X1 U658 ( .A(G171), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G92), .A2(n649), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G79), .A2(n646), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G66), .A2(n659), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G54), .A2(n660), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U667 ( .A(KEYINPUT15), .B(n593), .Z(n989) );
  OR2_X1 U668 ( .A1(n989), .A2(G868), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(G284) );
  INV_X1 U670 ( .A(G868), .ZN(n596) );
  NOR2_X1 U671 ( .A1(G286), .A2(n596), .ZN(n598) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U673 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n600), .A2(n989), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n978), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n989), .A2(G868), .ZN(n602) );
  NOR2_X1 U679 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(G282) );
  XNOR2_X1 U681 ( .A(G2100), .B(KEYINPUT79), .ZN(n617) );
  NAND2_X1 U682 ( .A1(G123), .A2(n521), .ZN(n605) );
  XOR2_X1 U683 ( .A(KEYINPUT75), .B(n605), .Z(n606) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT18), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G135), .A2(n898), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT76), .B(n609), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G111), .A2(n894), .ZN(n611) );
  NAND2_X1 U689 ( .A1(G99), .A2(n897), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U692 ( .A(KEYINPUT77), .B(n614), .Z(n936) );
  XNOR2_X1 U693 ( .A(n936), .B(G2096), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n615), .B(KEYINPUT78), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G93), .A2(n649), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G80), .A2(n646), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G67), .A2(n659), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G55), .A2(n660), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U702 ( .A(KEYINPUT81), .B(n622), .Z(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n667) );
  XNOR2_X1 U704 ( .A(n667), .B(KEYINPUT82), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n978), .B(KEYINPUT80), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n989), .A2(G559), .ZN(n625) );
  XNOR2_X1 U707 ( .A(n626), .B(n625), .ZN(n672) );
  NOR2_X1 U708 ( .A1(n672), .A2(G860), .ZN(n627) );
  XNOR2_X1 U709 ( .A(n628), .B(n627), .ZN(G145) );
  NAND2_X1 U710 ( .A1(G73), .A2(n646), .ZN(n629) );
  XNOR2_X1 U711 ( .A(n629), .B(KEYINPUT2), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G86), .A2(n649), .ZN(n631) );
  NAND2_X1 U713 ( .A1(G48), .A2(n660), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n659), .A2(G61), .ZN(n632) );
  XOR2_X1 U716 ( .A(KEYINPUT84), .B(n632), .Z(n633) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U719 ( .A1(G62), .A2(n659), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n637), .B(KEYINPUT85), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n649), .A2(G88), .ZN(n638) );
  XNOR2_X1 U722 ( .A(n638), .B(KEYINPUT86), .ZN(n640) );
  NAND2_X1 U723 ( .A1(G75), .A2(n646), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U725 ( .A(KEYINPUT87), .B(n641), .Z(n642) );
  NOR2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n660), .A2(G50), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(G303) );
  INV_X1 U729 ( .A(G303), .ZN(G166) );
  NAND2_X1 U730 ( .A1(G72), .A2(n646), .ZN(n648) );
  NAND2_X1 U731 ( .A1(G60), .A2(n659), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G85), .A2(n649), .ZN(n650) );
  XNOR2_X1 U734 ( .A(KEYINPUT65), .B(n650), .ZN(n651) );
  NOR2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n660), .A2(G47), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n654), .A2(n653), .ZN(G290) );
  NAND2_X1 U738 ( .A1(G651), .A2(G74), .ZN(n657) );
  NAND2_X1 U739 ( .A1(G87), .A2(n655), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U741 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U742 ( .A1(G49), .A2(n660), .ZN(n661) );
  XOR2_X1 U743 ( .A(KEYINPUT83), .B(n661), .Z(n662) );
  NAND2_X1 U744 ( .A1(n663), .A2(n662), .ZN(G288) );
  NOR2_X1 U745 ( .A1(G868), .A2(n667), .ZN(n664) );
  XNOR2_X1 U746 ( .A(n664), .B(KEYINPUT89), .ZN(n675) );
  XOR2_X1 U747 ( .A(KEYINPUT88), .B(KEYINPUT19), .Z(n665) );
  XNOR2_X1 U748 ( .A(G305), .B(n665), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n667), .B(n666), .ZN(n669) );
  XNOR2_X1 U750 ( .A(G299), .B(G166), .ZN(n668) );
  XNOR2_X1 U751 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(G290), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n671), .B(G288), .ZN(n909) );
  XNOR2_X1 U754 ( .A(n909), .B(n672), .ZN(n673) );
  NAND2_X1 U755 ( .A1(G868), .A2(n673), .ZN(n674) );
  NAND2_X1 U756 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U763 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U767 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G96), .A2(n682), .ZN(n834) );
  NAND2_X1 U769 ( .A1(n834), .A2(G2106), .ZN(n686) );
  NAND2_X1 U770 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U771 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U772 ( .A1(G108), .A2(n684), .ZN(n835) );
  NAND2_X1 U773 ( .A1(n835), .A2(G567), .ZN(n685) );
  NAND2_X1 U774 ( .A1(n686), .A2(n685), .ZN(n919) );
  NOR2_X1 U775 ( .A1(n687), .A2(n919), .ZN(n688) );
  XNOR2_X1 U776 ( .A(n688), .B(KEYINPUT90), .ZN(n833) );
  NAND2_X1 U777 ( .A1(G36), .A2(n833), .ZN(G176) );
  AND2_X1 U778 ( .A1(G40), .A2(n690), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n792) );
  INV_X1 U780 ( .A(n792), .ZN(n693) );
  INV_X1 U781 ( .A(G1996), .ZN(n815) );
  XNOR2_X1 U782 ( .A(n695), .B(n694), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n733), .A2(G1341), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n704), .A2(n989), .ZN(n702) );
  INV_X1 U786 ( .A(n733), .ZN(n718) );
  NOR2_X1 U787 ( .A1(n718), .A2(G1348), .ZN(n700) );
  NOR2_X1 U788 ( .A1(G2067), .A2(n733), .ZN(n699) );
  NOR2_X1 U789 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U790 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U791 ( .A(n703), .B(KEYINPUT101), .ZN(n706) );
  NOR2_X1 U792 ( .A1(n989), .A2(n704), .ZN(n705) );
  NOR2_X1 U793 ( .A1(n706), .A2(n705), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n718), .A2(G2072), .ZN(n707) );
  XOR2_X1 U795 ( .A(KEYINPUT27), .B(n707), .Z(n709) );
  NAND2_X1 U796 ( .A1(G1956), .A2(n733), .ZN(n708) );
  NAND2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U798 ( .A1(G299), .A2(n713), .ZN(n710) );
  XNOR2_X1 U799 ( .A(n710), .B(KEYINPUT102), .ZN(n711) );
  NOR2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U801 ( .A1(G299), .A2(n713), .ZN(n714) );
  XOR2_X1 U802 ( .A(KEYINPUT28), .B(n714), .Z(n715) );
  NOR2_X1 U803 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U804 ( .A(n717), .B(KEYINPUT29), .ZN(n722) );
  NAND2_X1 U805 ( .A1(G1961), .A2(n733), .ZN(n720) );
  XOR2_X1 U806 ( .A(G2078), .B(KEYINPUT25), .Z(n951) );
  NAND2_X1 U807 ( .A1(n718), .A2(n951), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n723) );
  OR2_X1 U809 ( .A1(n723), .A2(G301), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n732) );
  NAND2_X1 U811 ( .A1(G301), .A2(n723), .ZN(n724) );
  XNOR2_X1 U812 ( .A(n724), .B(KEYINPUT103), .ZN(n729) );
  NAND2_X1 U813 ( .A1(G8), .A2(n733), .ZN(n776) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n776), .ZN(n745) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n733), .ZN(n742) );
  NOR2_X1 U816 ( .A1(n745), .A2(n742), .ZN(n725) );
  NAND2_X1 U817 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U819 ( .A1(n727), .A2(G168), .ZN(n728) );
  XOR2_X1 U820 ( .A(KEYINPUT31), .B(n730), .Z(n731) );
  NAND2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n743) );
  NAND2_X1 U822 ( .A1(n743), .A2(G286), .ZN(n740) );
  INV_X1 U823 ( .A(G8), .ZN(n738) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n776), .ZN(n735) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U829 ( .A(n741), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U830 ( .A1(G8), .A2(n742), .ZN(n747) );
  INV_X1 U831 ( .A(n743), .ZN(n744) );
  NOR2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n749), .A2(n748), .ZN(n775) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n982) );
  XNOR2_X1 U836 ( .A(KEYINPUT104), .B(n982), .ZN(n750) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n775), .A2(n751), .ZN(n755) );
  INV_X1 U839 ( .A(n776), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n752), .A2(KEYINPUT105), .ZN(n753) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n974) );
  AND2_X1 U842 ( .A1(n753), .A2(n974), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n758) );
  INV_X1 U844 ( .A(n974), .ZN(n756) );
  OR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n980) );
  OR2_X1 U846 ( .A1(n756), .A2(n980), .ZN(n757) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n984) );
  NOR2_X1 U848 ( .A1(KEYINPUT105), .A2(n776), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n984), .A2(n761), .ZN(n759) );
  INV_X1 U850 ( .A(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n759), .A2(n760), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n980), .A2(n760), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U855 ( .A(n767), .B(KEYINPUT106), .ZN(n772) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XOR2_X1 U857 ( .A(n768), .B(KEYINPUT24), .Z(n769) );
  XNOR2_X1 U858 ( .A(KEYINPUT100), .B(n769), .ZN(n770) );
  NOR2_X1 U859 ( .A1(n776), .A2(n770), .ZN(n771) );
  NOR2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n779) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n795) );
  XNOR2_X1 U866 ( .A(KEYINPUT37), .B(G2067), .ZN(n814) );
  XNOR2_X1 U867 ( .A(KEYINPUT95), .B(KEYINPUT36), .ZN(n791) );
  NAND2_X1 U868 ( .A1(n894), .A2(G116), .ZN(n780) );
  XNOR2_X1 U869 ( .A(n780), .B(KEYINPUT94), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G128), .A2(n521), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(KEYINPUT35), .ZN(n789) );
  XNOR2_X1 U873 ( .A(KEYINPUT93), .B(KEYINPUT34), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G104), .A2(n897), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G140), .A2(n898), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U877 ( .A(n787), .B(n786), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U879 ( .A(n791), .B(n790), .ZN(n890) );
  NOR2_X1 U880 ( .A1(n814), .A2(n890), .ZN(n925) );
  NOR2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n825) );
  NAND2_X1 U882 ( .A1(n925), .A2(n825), .ZN(n794) );
  XNOR2_X1 U883 ( .A(n794), .B(KEYINPUT96), .ZN(n823) );
  XNOR2_X1 U884 ( .A(KEYINPUT97), .B(G1991), .ZN(n958) );
  NAND2_X1 U885 ( .A1(G107), .A2(n894), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G95), .A2(n897), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G119), .A2(n521), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G131), .A2(n898), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n884) );
  OR2_X1 U892 ( .A1(n958), .A2(n884), .ZN(n811) );
  NAND2_X1 U893 ( .A1(G129), .A2(n521), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G117), .A2(n894), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U896 ( .A(KEYINPUT98), .B(n804), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n897), .A2(G105), .ZN(n805) );
  XNOR2_X1 U898 ( .A(n805), .B(KEYINPUT38), .ZN(n807) );
  NAND2_X1 U899 ( .A1(G141), .A2(n898), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n889) );
  OR2_X1 U902 ( .A1(n815), .A2(n889), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n940) );
  NAND2_X1 U904 ( .A1(n825), .A2(n940), .ZN(n818) );
  XNOR2_X1 U905 ( .A(KEYINPUT99), .B(n818), .ZN(n812) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n986) );
  NAND2_X1 U907 ( .A1(n525), .A2(n813), .ZN(n828) );
  NAND2_X1 U908 ( .A1(n814), .A2(n890), .ZN(n926) );
  NAND2_X1 U909 ( .A1(n889), .A2(n815), .ZN(n920) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n816) );
  XNOR2_X1 U911 ( .A(KEYINPUT107), .B(n816), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n884), .A2(n958), .ZN(n937) );
  NAND2_X1 U913 ( .A1(n817), .A2(n937), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n920), .A2(n820), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT39), .B(n821), .Z(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n926), .A2(n824), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT40), .B(n829), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U924 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U933 ( .A(G2454), .B(G2446), .ZN(n844) );
  XNOR2_X1 U934 ( .A(G2430), .B(G2443), .ZN(n842) );
  XOR2_X1 U935 ( .A(G2435), .B(KEYINPUT108), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2451), .B(G2438), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U938 ( .A(n838), .B(G2427), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1341), .B(G1348), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n845) );
  NAND2_X1 U943 ( .A1(n845), .A2(G14), .ZN(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT109), .B(n846), .ZN(G401) );
  XOR2_X1 U945 ( .A(G2100), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2072), .B(KEYINPUT110), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n849), .B(G2678), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2090), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U951 ( .A(KEYINPUT42), .B(G2096), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1976), .B(G1961), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1966), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U958 ( .A(G1971), .B(G1956), .Z(n859) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U962 ( .A(KEYINPUT111), .B(G2474), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n865) );
  XOR2_X1 U964 ( .A(G1981), .B(KEYINPUT41), .Z(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(G229) );
  XOR2_X1 U966 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n867) );
  NAND2_X1 U967 ( .A1(G124), .A2(n521), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n874) );
  NAND2_X1 U969 ( .A1(G112), .A2(n894), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G100), .A2(n897), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n870), .B(KEYINPUT113), .ZN(n872) );
  NAND2_X1 U973 ( .A1(G136), .A2(n898), .ZN(n871) );
  NAND2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G103), .A2(n897), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G139), .A2(n898), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G127), .A2(n521), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G115), .A2(n894), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT114), .B(n879), .Z(n880) );
  XNOR2_X1 U983 ( .A(KEYINPUT47), .B(n880), .ZN(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n928) );
  XNOR2_X1 U985 ( .A(G164), .B(n928), .ZN(n883) );
  XNOR2_X1 U986 ( .A(n883), .B(G162), .ZN(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n886) );
  XNOR2_X1 U988 ( .A(n884), .B(n936), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n888), .B(n887), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n906) );
  NAND2_X1 U993 ( .A1(G130), .A2(n521), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G118), .A2(n894), .ZN(n895) );
  NAND2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U996 ( .A1(G106), .A2(n897), .ZN(n900) );
  NAND2_X1 U997 ( .A1(G142), .A2(n898), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U999 ( .A(KEYINPUT45), .B(n901), .Z(n902) );
  NOR2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(G160), .B(n904), .Z(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(n908) );
  XOR2_X1 U1004 ( .A(KEYINPUT115), .B(n908), .Z(G395) );
  XOR2_X1 U1005 ( .A(n909), .B(G286), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G171), .B(n989), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(n978), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n913), .ZN(G397) );
  OR2_X1 U1010 ( .A1(n919), .A2(G401), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n919), .ZN(G319) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1019 ( .A(G2090), .B(G162), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n922), .B(KEYINPUT51), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT116), .B(n923), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n934) );
  XOR2_X1 U1025 ( .A(n928), .B(KEYINPUT117), .Z(n929) );
  XOR2_X1 U1026 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1029 ( .A(KEYINPUT50), .B(n932), .Z(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n942) );
  XOR2_X1 U1031 ( .A(G2084), .B(G160), .Z(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(KEYINPUT118), .B(n943), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT52), .B(n944), .Z(n946) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n948) );
  XOR2_X1 U1041 ( .A(KEYINPUT119), .B(n948), .Z(n1030) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(n951), .B(G27), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT121), .B(n956), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(G28), .ZN(n961) );
  XOR2_X1 U1051 ( .A(KEYINPUT120), .B(n958), .Z(n959) );
  XNOR2_X1 U1052 ( .A(G25), .B(n959), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1054 ( .A(KEYINPUT53), .B(n962), .Z(n965) );
  XOR2_X1 U1055 ( .A(KEYINPUT54), .B(G34), .Z(n963) );
  XNOR2_X1 U1056 ( .A(G2084), .B(n963), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(KEYINPUT55), .B(n968), .ZN(n970) );
  INV_X1 U1061 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n971), .A2(G11), .ZN(n1028) );
  INV_X1 U1064 ( .A(G16), .ZN(n1024) );
  XOR2_X1 U1065 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n972) );
  XNOR2_X1 U1066 ( .A(n1024), .B(n972), .ZN(n1000) );
  XOR2_X1 U1067 ( .A(G1966), .B(G168), .Z(n973) );
  XNOR2_X1 U1068 ( .A(KEYINPUT123), .B(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT57), .ZN(n998) );
  XOR2_X1 U1071 ( .A(G1341), .B(KEYINPUT125), .Z(n977) );
  XNOR2_X1 U1072 ( .A(n978), .B(n977), .ZN(n996) );
  XOR2_X1 U1073 ( .A(G1956), .B(G299), .Z(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n988) );
  NAND2_X1 U1076 ( .A1(G1971), .A2(G303), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(n989), .B(G1348), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G171), .B(G1961), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1084 ( .A(KEYINPUT124), .B(n994), .Z(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  XOR2_X1 U1088 ( .A(G1986), .B(G24), .Z(n1003) );
  XNOR2_X1 U1089 ( .A(KEYINPUT127), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(n1001), .B(G1971), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1006), .Z(n1021) );
  XOR2_X1 U1095 ( .A(G1961), .B(G5), .Z(n1016) );
  XNOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(G4), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(G6), .B(G1981), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G20), .B(G1956), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G21), .B(G1966), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(KEYINPUT126), .B(n1019), .Z(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

