//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n206), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n202), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT66), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n208), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n217), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n250), .A2(new_n252), .B1(new_n201), .B2(new_n206), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n206), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n253), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n215), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G50), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n260), .B1(new_n205), .B2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n270), .B2(new_n267), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT9), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n262), .A2(KEYINPUT9), .A3(new_n271), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT10), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  AND2_X1   g0077(.A1(G1), .A2(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G226), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n281), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n291), .A2(G222), .ZN(new_n292));
  AND2_X1   g0092(.A1(G223), .A2(G1698), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n202), .B2(new_n290), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT68), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n285), .B1(new_n295), .B2(new_n296), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n287), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G190), .ZN(new_n300));
  INV_X1    g0100(.A(new_n299), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n275), .A2(new_n276), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n300), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n273), .A2(new_n274), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT10), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n309), .B1(G169), .B2(new_n299), .C1(new_n262), .C2(new_n271), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n220), .B1(new_n270), .B2(KEYINPUT12), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n206), .A2(G68), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(G50), .B2(new_n251), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n202), .B2(new_n256), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n260), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n313), .B1(new_n318), .B2(KEYINPUT11), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT12), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n320), .A2(new_n263), .A3(G1), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n320), .A2(new_n265), .B1(new_n321), .B2(new_n314), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT73), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n324), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n312), .B1(new_n323), .B2(new_n317), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT73), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT72), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n283), .B1(new_n221), .B2(new_n286), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n236), .A2(G1698), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n336), .B1(G226), .B2(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G97), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n285), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n333), .B1(new_n335), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n285), .B1(new_n339), .B2(new_n340), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n345), .A2(new_n334), .A3(KEYINPUT13), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n332), .B(G169), .C1(new_n344), .C2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n335), .A2(new_n343), .A3(new_n333), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT13), .B1(new_n345), .B2(new_n334), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(G179), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G169), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n348), .B2(new_n349), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n332), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n331), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n347), .A2(new_n350), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n357), .A2(new_n354), .A3(KEYINPUT72), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n330), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n326), .A2(new_n327), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n348), .A2(new_n349), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(G200), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n348), .A2(new_n349), .A3(G190), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT74), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n284), .B2(G1698), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n290), .B1(G33), .B2(G87), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n366), .B1(new_n369), .B2(new_n285), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n284), .A2(G1698), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G223), .B2(G1698), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n337), .A2(new_n338), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(KEYINPUT74), .A3(new_n342), .ZN(new_n376));
  INV_X1    g0176(.A(G190), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n285), .A2(G232), .A3(new_n281), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n283), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n370), .A2(new_n376), .A3(new_n377), .A4(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n369), .A2(new_n285), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n288), .A2(new_n206), .A3(new_n289), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT7), .B1(new_n374), .B2(new_n206), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G58), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n220), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n251), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n386), .A2(new_n387), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n374), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n220), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n402), .B2(new_n396), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(new_n403), .A3(new_n260), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n255), .A2(new_n265), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n269), .B2(new_n255), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n385), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT17), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n385), .A2(new_n404), .A3(new_n406), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n404), .A2(new_n406), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n283), .A2(new_n378), .A3(new_n308), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n370), .A2(new_n376), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n370), .A2(new_n376), .A3(KEYINPUT75), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n380), .B1(new_n285), .B2(new_n369), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n352), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n412), .A2(new_n418), .A3(new_n423), .A4(new_n420), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n411), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT70), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n254), .B(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(new_n252), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n260), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT71), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n270), .B2(new_n202), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n269), .A2(KEYINPUT71), .A3(G77), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n266), .A2(new_n202), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G238), .A2(G1698), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n290), .B(new_n439), .C1(new_n236), .C2(G1698), .ZN(new_n440));
  INV_X1    g0240(.A(G107), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n374), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n342), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n285), .A2(G244), .A3(new_n281), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n283), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n352), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n443), .A2(new_n308), .A3(new_n283), .A4(new_n445), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n438), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n431), .A2(new_n260), .B1(new_n202), .B2(new_n266), .ZN(new_n450));
  OAI21_X1  g0250(.A(G200), .B1(new_n444), .B2(new_n446), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n443), .A2(G190), .A3(new_n283), .A4(new_n445), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n450), .A2(new_n436), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NOR4_X1   g0254(.A1(new_n311), .A2(new_n365), .A3(new_n425), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G116), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G20), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT23), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n206), .B2(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n441), .A2(KEYINPUT23), .A3(G20), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n206), .B(G87), .C1(new_n337), .C2(new_n338), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n462), .A2(KEYINPUT22), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(KEYINPUT22), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT24), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n462), .B(KEYINPUT22), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(new_n461), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n260), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n205), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n261), .A2(new_n265), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n441), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT25), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n265), .B2(G107), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n473), .A2(G107), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G250), .B(new_n291), .C1(new_n337), .C2(new_n338), .ZN(new_n478));
  AND2_X1   g0278(.A1(G257), .A2(G1698), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n337), .B2(new_n338), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G294), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n342), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  INV_X1    g0285(.A(G41), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G41), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G264), .A3(new_n285), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n205), .B(G45), .C1(new_n486), .C2(KEYINPUT5), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n488), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n280), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n483), .A2(new_n377), .A3(new_n491), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n483), .A2(new_n491), .A3(new_n495), .ZN(new_n497));
  AOI22_X1  g0297(.A1(KEYINPUT84), .A2(new_n496), .B1(new_n497), .B2(new_n382), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n497), .A2(KEYINPUT84), .A3(new_n382), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n470), .B(new_n477), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n497), .A2(G179), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n352), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n465), .A2(KEYINPUT24), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n468), .A2(new_n467), .A3(new_n461), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n261), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n477), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n501), .B(new_n502), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT85), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n500), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n500), .B2(new_n507), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G303), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n288), .A2(new_n513), .A3(new_n289), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G264), .A2(G1698), .ZN(new_n515));
  INV_X1    g0315(.A(G257), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(G1698), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n514), .B(new_n342), .C1(new_n374), .C2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G270), .B(new_n285), .C1(new_n492), .C2(new_n493), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT80), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n490), .A2(KEYINPUT80), .A3(G270), .A4(new_n285), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n495), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n519), .A2(new_n520), .B1(new_n494), .B2(new_n280), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT81), .B1(new_n526), .B2(new_n522), .ZN(new_n527));
  OAI211_X1 g0327(.A(G190), .B(new_n518), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n266), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT82), .B1(new_n265), .B2(G116), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n473), .A2(G116), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  INV_X1    g0335(.A(G97), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n206), .C1(G33), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(G20), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n260), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT20), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n534), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n260), .A2(new_n538), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(KEYINPUT83), .A3(KEYINPUT20), .A4(new_n537), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n539), .A2(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n533), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n518), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n523), .A2(new_n524), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n526), .A2(KEYINPUT81), .A3(new_n522), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n528), .B(new_n547), .C1(new_n382), .C2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n518), .B1(new_n525), .B2(new_n527), .ZN(new_n553));
  NAND2_X1  g0353(.A1(KEYINPUT21), .A2(G169), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n533), .B2(new_n545), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n518), .A2(G179), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n549), .B2(new_n550), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n553), .A2(new_n555), .B1(new_n557), .B2(new_n546), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n546), .A2(G169), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(new_n551), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n552), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n265), .A2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n472), .B2(new_n536), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n441), .B1(new_n400), .B2(new_n401), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n568));
  OR2_X1    g0368(.A1(KEYINPUT6), .A2(G97), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n441), .A2(KEYINPUT76), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT76), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(G107), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(new_n568), .ZN(new_n574));
  XNOR2_X1  g0374(.A(KEYINPUT76), .B(G107), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n206), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n252), .A2(new_n202), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n567), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n566), .B1(new_n579), .B2(new_n261), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n490), .A2(G257), .A3(new_n285), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n495), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G250), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n288), .B2(new_n289), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT4), .ZN(new_n585));
  OAI21_X1  g0385(.A(G1698), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n374), .B2(new_n222), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n585), .A2(G1698), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(G244), .C1(new_n338), .C2(new_n337), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n586), .A2(new_n535), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n582), .B1(new_n590), .B2(new_n342), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n308), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n222), .B1(new_n288), .B2(new_n289), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n589), .B(new_n535), .C1(new_n593), .C2(KEYINPUT4), .ZN(new_n594));
  OAI21_X1  g0394(.A(G250), .B1(new_n337), .B2(new_n338), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n291), .B1(new_n595), .B2(KEYINPUT4), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n342), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n582), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n352), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n580), .A2(new_n592), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n576), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n574), .A2(new_n575), .ZN(new_n603));
  OAI21_X1  g0403(.A(G20), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(G107), .B1(new_n388), .B2(new_n389), .ZN(new_n605));
  INV_X1    g0405(.A(new_n578), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n565), .B1(new_n607), .B2(new_n260), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n591), .A2(G190), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n599), .A2(G200), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n613));
  AND2_X1   g0413(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n614));
  NOR2_X1   g0414(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n615));
  OAI211_X1 g0415(.A(G33), .B(G97), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n613), .B1(new_n616), .B2(new_n206), .ZN(new_n617));
  OR2_X1    g0417(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n618));
  NAND2_X1  g0418(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n618), .B(new_n619), .C1(new_n256), .C2(new_n536), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n206), .B(G68), .C1(new_n337), .C2(new_n338), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n260), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n473), .A2(new_n427), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n266), .A2(new_n426), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT79), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT79), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n623), .A2(new_n624), .A3(new_n628), .A4(new_n625), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n285), .B(G250), .C1(G1), .C2(new_n484), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n285), .A2(G274), .A3(new_n485), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT77), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n280), .A2(KEYINPUT77), .A3(new_n485), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n221), .A2(new_n291), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n222), .A2(G1698), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n637), .B(new_n638), .C1(new_n337), .C2(new_n338), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n456), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n342), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n636), .A2(new_n308), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n634), .A2(new_n635), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n641), .A3(new_n630), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n352), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n627), .A2(new_n629), .A3(new_n642), .A4(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n644), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G190), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(G200), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n473), .A2(G87), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n623), .A2(new_n650), .A3(new_n625), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n612), .A2(new_n654), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n455), .A2(new_n512), .A3(new_n562), .A4(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n449), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n364), .A2(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n359), .A2(new_n658), .B1(new_n408), .B2(new_n410), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n422), .A2(new_n424), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n307), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(new_n310), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT87), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n648), .A2(new_n652), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n632), .A2(new_n633), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT77), .B1(new_n280), .B2(new_n485), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n630), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT86), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n668), .A2(new_n669), .B1(new_n342), .B2(new_n640), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n636), .A2(KEYINPUT86), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n382), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(G169), .B1(new_n670), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n642), .A2(new_n626), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n665), .A2(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n663), .B(new_n664), .C1(new_n675), .C2(new_n601), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n646), .A2(new_n653), .ZN(new_n677));
  INV_X1    g0477(.A(new_n601), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(KEYINPUT26), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n670), .A2(new_n671), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G200), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n651), .B1(G190), .B2(new_n647), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n674), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n641), .B1(new_n636), .B2(KEYINPUT86), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n668), .A2(new_n669), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n352), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n678), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n663), .B1(new_n690), .B2(new_n664), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n601), .A2(new_n611), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n682), .A2(new_n683), .B1(new_n685), .B2(new_n688), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n500), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n558), .A2(new_n507), .A3(new_n561), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n689), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n455), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n662), .A2(new_n700), .ZN(G369));
  NAND2_X1  g0501(.A1(new_n264), .A2(new_n206), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT88), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n702), .B(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(G213), .B1(new_n704), .B2(KEYINPUT27), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n702), .B(KEYINPUT88), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT27), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n558), .B2(new_n561), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n512), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n507), .ZN(new_n713));
  INV_X1    g0513(.A(new_n710), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n470), .A2(new_n477), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n511), .B1(new_n718), .B2(new_n710), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n713), .B2(new_n710), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n558), .A2(new_n561), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n710), .A2(new_n546), .ZN(new_n722));
  MUX2_X1   g0522(.A(new_n721), .B(new_n562), .S(new_n722), .Z(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n717), .B1(new_n720), .B2(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n209), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n613), .A2(new_n530), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n727), .A2(new_n205), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n214), .B2(new_n727), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n714), .C1(new_n692), .C2(new_n698), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT89), .B1(new_n695), .B2(new_n697), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n500), .A2(new_n601), .A3(new_n611), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT89), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n694), .A4(new_n696), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n690), .A2(KEYINPUT26), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n677), .A2(new_n664), .A3(new_n678), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n739), .A2(new_n689), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n710), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n733), .B1(new_n742), .B2(new_n732), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G330), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n549), .A2(new_n550), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n483), .A2(G179), .A3(new_n491), .A4(new_n518), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n644), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n746), .A2(new_n748), .A3(new_n591), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n497), .A2(new_n308), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n591), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(new_n553), .A3(new_n681), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n746), .A2(new_n748), .A3(KEYINPUT30), .A4(new_n591), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n751), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT31), .B1(new_n756), .B2(new_n710), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n612), .A2(new_n654), .A3(new_n710), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n760), .B(new_n562), .C1(new_n509), .C2(new_n510), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n745), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n744), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n731), .B1(new_n765), .B2(G1), .ZN(G364));
  INV_X1    g0566(.A(new_n727), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n263), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G45), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n767), .A2(G1), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n723), .B2(G330), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n723), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n726), .A2(new_n374), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G355), .B1(new_n530), .B2(new_n726), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n245), .A2(new_n484), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n209), .A2(new_n374), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT90), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n213), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n775), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT91), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n215), .B1(G20), .B2(new_n352), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n782), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G179), .A2(G200), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n206), .B1(new_n790), .B2(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n536), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n206), .A2(G190), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n382), .A2(G179), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G87), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n206), .A2(new_n377), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n794), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n290), .B1(new_n795), .B2(new_n441), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n377), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n792), .B(new_n799), .C1(G50), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n308), .A2(G200), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT92), .ZN(new_n804));
  AND3_X1   g0604(.A1(new_n803), .A2(new_n793), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n803), .B2(new_n793), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n797), .A2(new_n803), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n807), .A2(new_n202), .B1(new_n391), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT93), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n793), .A2(new_n790), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n814));
  XNOR2_X1  g0614(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n800), .A2(G190), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(G68), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n809), .A2(KEYINPUT93), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n802), .A2(new_n810), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n807), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G311), .ZN(new_n821));
  INV_X1    g0621(.A(new_n795), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n290), .B1(new_n822), .B2(G283), .ZN(new_n823));
  INV_X1    g0623(.A(new_n798), .ZN(new_n824));
  INV_X1    g0624(.A(new_n811), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G303), .A2(new_n824), .B1(new_n825), .B2(G329), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n791), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G326), .B2(new_n801), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n821), .A2(new_n823), .A3(new_n826), .A4(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n816), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT33), .B(G317), .Z(new_n832));
  INV_X1    g0632(.A(G322), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n831), .A2(new_n832), .B1(new_n808), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT95), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n819), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n770), .B1(new_n836), .B2(new_n787), .ZN(new_n837));
  INV_X1    g0637(.A(new_n786), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n789), .B(new_n837), .C1(new_n723), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n773), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  NAND2_X1  g0641(.A1(new_n438), .A2(new_n710), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n449), .A2(new_n453), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT98), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n657), .A2(new_n710), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT98), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n449), .A2(new_n842), .A3(new_n846), .A4(new_n453), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT99), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n848), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n699), .B2(new_n714), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n851), .A2(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n844), .A2(new_n847), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n714), .B(new_n853), .C1(new_n692), .C2(new_n698), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n851), .B2(KEYINPUT100), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(new_n763), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(KEYINPUT101), .A3(new_n763), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n857), .A2(new_n770), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n856), .A2(new_n763), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n787), .A2(new_n784), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n770), .B1(new_n202), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n822), .A2(G87), .B1(new_n825), .B2(G311), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(KEYINPUT96), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(G116), .B2(new_n820), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n801), .A2(G303), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n792), .B1(new_n816), .B2(G283), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n374), .B1(new_n798), .B2(new_n441), .C1(new_n827), .C2(new_n808), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(KEYINPUT96), .B2(new_n865), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n808), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(G143), .B1(G150), .B2(new_n816), .ZN(new_n874));
  INV_X1    g0674(.A(G137), .ZN(new_n875));
  INV_X1    g0675(.A(new_n801), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .C1(new_n807), .C2(new_n812), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT34), .Z(new_n878));
  AOI22_X1  g0678(.A1(G50), .A2(new_n824), .B1(new_n825), .B2(G132), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n374), .B1(new_n822), .B2(G68), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n879), .B(new_n880), .C1(new_n391), .C2(new_n791), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n872), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT97), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n787), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n882), .A2(KEYINPUT97), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n864), .B1(new_n785), .B2(new_n848), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n862), .A2(new_n886), .ZN(G384));
  NOR2_X1   g0687(.A1(new_n602), .A2(new_n603), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n889), .A2(KEYINPUT35), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(KEYINPUT35), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(G116), .A3(new_n216), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT36), .Z(new_n893));
  OAI211_X1 g0693(.A(new_n214), .B(G77), .C1(new_n391), .C2(new_n220), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n267), .A2(G68), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n205), .B(G13), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n705), .A2(new_n708), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n412), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n421), .A2(new_n407), .A3(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n421), .A2(new_n900), .A3(new_n407), .A4(new_n902), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT105), .ZN(new_n908));
  INV_X1    g0708(.A(new_n900), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n908), .B1(new_n425), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n425), .A2(new_n909), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n908), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n905), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(KEYINPUT104), .B1(new_n425), .B2(new_n909), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT104), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n921), .A3(new_n905), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(KEYINPUT38), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n898), .B1(new_n917), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n325), .A2(new_n329), .A3(new_n710), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT102), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n359), .A2(new_n927), .A3(new_n364), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n351), .A2(new_n355), .A3(new_n331), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT72), .B1(new_n357), .B2(new_n354), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n364), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n330), .A3(new_n710), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n925), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n759), .A2(new_n761), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT106), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n935), .A2(KEYINPUT106), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n924), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n919), .A2(KEYINPUT104), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(new_n922), .A3(new_n912), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n916), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n923), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n898), .B1(new_n943), .B2(new_n935), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n938), .A2(G330), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n455), .A2(new_n762), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT107), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n938), .A2(new_n944), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n455), .A2(new_n934), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND4_X1   g0752(.A1(KEYINPUT38), .A2(new_n939), .A3(new_n922), .A4(new_n912), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT38), .B1(new_n920), .B2(new_n922), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT39), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT39), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n912), .A2(KEYINPUT105), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n957), .A2(new_n910), .A3(new_n907), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n923), .B(new_n956), .C1(new_n958), .C2(KEYINPUT38), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n359), .A2(new_n710), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n928), .A2(new_n932), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n449), .A2(new_n710), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n963), .B1(new_n854), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n966), .A2(new_n942), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n899), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n660), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n743), .A2(new_n455), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n662), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n971), .B(new_n973), .Z(new_n974));
  OAI22_X1  g0774(.A1(new_n952), .A2(new_n974), .B1(new_n205), .B2(new_n768), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n952), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n897), .B1(new_n975), .B2(new_n976), .ZN(G367));
  XOR2_X1   g0777(.A(new_n727), .B(KEYINPUT41), .Z(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  MUX2_X1   g0779(.A(new_n720), .B(new_n512), .S(new_n711), .Z(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n724), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(new_n764), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n678), .A2(new_n710), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT108), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n693), .B1(new_n608), .B2(new_n714), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n716), .A2(new_n987), .A3(KEYINPUT109), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT109), .B1(new_n716), .B2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n716), .A2(new_n987), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n716), .A2(KEYINPUT44), .A3(new_n987), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n720), .A2(new_n724), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT110), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n995), .A2(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n988), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n992), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n997), .A2(new_n998), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n982), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n979), .B1(new_n1005), .B2(new_n764), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n769), .A2(G1), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n710), .A2(new_n651), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n694), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n689), .B2(new_n1010), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n986), .A2(new_n512), .A3(new_n711), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT42), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n678), .B1(new_n986), .B2(new_n713), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n1016), .B2(new_n710), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1014), .A2(KEYINPUT42), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1019), .B(new_n1020), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n997), .A2(new_n986), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1009), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n791), .A2(new_n220), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n374), .B(new_n1025), .C1(G77), .C2(new_n822), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n820), .A2(G50), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G143), .A2(new_n801), .B1(new_n816), .B2(G159), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n808), .A2(new_n250), .B1(new_n811), .B2(new_n875), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G58), .B2(new_n824), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n290), .B1(new_n825), .B2(G317), .ZN(new_n1032));
  INV_X1    g0832(.A(G283), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n536), .B2(new_n795), .C1(new_n807), .C2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n798), .A2(new_n530), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT46), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n831), .B2(new_n827), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1035), .A2(KEYINPUT46), .B1(new_n441), .B2(new_n791), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n873), .A2(G303), .B1(G311), .B2(new_n801), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT111), .Z(new_n1041));
  OAI21_X1  g0841(.A(new_n1031), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT47), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n787), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n778), .A2(new_n240), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n788), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n726), .B2(new_n427), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n770), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1044), .B(new_n1048), .C1(new_n838), .C2(new_n1012), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1024), .A2(new_n1049), .ZN(G387));
  NAND2_X1  g0850(.A1(new_n981), .A2(new_n764), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n982), .A2(new_n727), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n720), .A2(new_n786), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n824), .A2(G77), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n250), .B2(new_n811), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G50), .B2(new_n873), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n791), .A2(new_n426), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n290), .B1(new_n795), .B2(new_n536), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(G159), .C2(new_n801), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n820), .A2(G68), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n255), .A2(new_n816), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n290), .B1(new_n825), .B2(G326), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n798), .A2(new_n827), .B1(new_n791), .B2(new_n1033), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n873), .A2(G317), .B1(G311), .B2(new_n816), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n833), .B2(new_n876), .C1(new_n513), .C2(new_n807), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT49), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1063), .B1(new_n530), .B2(new_n795), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1062), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n787), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n774), .A2(new_n728), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(G107), .B2(new_n209), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n237), .A2(G45), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n778), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n430), .A2(G50), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  AOI211_X1 g0880(.A(G45), .B(new_n728), .C1(G68), .C2(G77), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1076), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n771), .B1(new_n1083), .B2(new_n1046), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT112), .Z(new_n1085));
  NAND3_X1  g0885(.A1(new_n1053), .A2(new_n1074), .A3(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1052), .B(new_n1086), .C1(new_n1008), .C2(new_n981), .ZN(G393));
  NOR2_X1   g0887(.A1(new_n1005), .A2(new_n767), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n982), .A2(new_n1004), .A3(new_n1003), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n430), .A2(new_n807), .ZN(new_n1091));
  INV_X1    g0891(.A(G143), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n798), .A2(new_n220), .B1(new_n811), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(KEYINPUT113), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n791), .A2(new_n202), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n290), .B1(new_n795), .B2(new_n796), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G50), .C2(new_n816), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1094), .B(new_n1097), .C1(KEYINPUT113), .C2(new_n1093), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n873), .A2(G159), .B1(G150), .B2(new_n801), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n798), .A2(new_n1033), .B1(new_n811), .B2(new_n833), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n290), .B(new_n1101), .C1(G107), .C2(new_n822), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n791), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1103), .A2(G116), .B1(G303), .B2(new_n816), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(new_n827), .C2(new_n807), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n873), .A2(G311), .B1(G317), .B2(new_n801), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1098), .A2(new_n1100), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n787), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n788), .B1(new_n536), .B2(new_n209), .C1(new_n1078), .C2(new_n248), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n771), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n987), .B2(new_n786), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n1007), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1090), .A2(new_n1114), .ZN(G390));
  NAND2_X1  g0915(.A1(new_n933), .A2(new_n762), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT114), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n966), .A2(new_n961), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n960), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n738), .A2(new_n741), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n714), .A3(new_n853), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n963), .B1(new_n1122), .B2(new_n965), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n961), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT38), .B1(new_n911), .B2(new_n914), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n953), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1123), .A2(new_n1126), .B1(KEYINPUT114), .B2(new_n1116), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1118), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1116), .A2(KEYINPUT114), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n961), .B1(new_n917), .B2(new_n923), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n928), .A2(new_n932), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n853), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n710), .B(new_n1132), .C1(new_n738), .C2(new_n741), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1131), .B1(new_n1133), .B2(new_n964), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1129), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n955), .B(new_n959), .C1(new_n966), .C2(new_n961), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1136), .A3(new_n1117), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1128), .A2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n745), .B(new_n925), .C1(new_n759), .C2(new_n761), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT115), .B1(new_n1139), .B2(new_n1131), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n934), .A2(G330), .A3(new_n848), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT115), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n963), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1116), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n854), .A2(new_n965), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1133), .A2(new_n964), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n762), .A2(new_n850), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1148), .A2(new_n963), .B1(new_n762), .B2(new_n933), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n972), .A2(new_n662), .A3(new_n946), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT116), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1144), .A2(new_n1145), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT116), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n1152), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1138), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1141), .A2(new_n963), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1159), .A2(KEYINPUT115), .B1(new_n762), .B2(new_n933), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1160), .A2(new_n1143), .B1(new_n854), .B2(new_n965), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1150), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1153), .B(KEYINPUT116), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1156), .B1(new_n1155), .B2(new_n1152), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1128), .A4(new_n1137), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1158), .A2(new_n727), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n955), .A2(new_n959), .A3(new_n784), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n863), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n771), .B1(new_n255), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n290), .B(new_n1095), .C1(G87), .C2(new_n824), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n820), .A2(G97), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G107), .A2(new_n816), .B1(new_n801), .B2(G283), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n795), .A2(new_n220), .B1(new_n811), .B2(new_n827), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G116), .B2(new_n873), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(G125), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n290), .B1(new_n811), .B2(new_n1176), .C1(new_n267), .C2(new_n795), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT117), .Z(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT54), .B(G143), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n820), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n798), .A2(new_n250), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1183), .A2(KEYINPUT53), .B1(new_n816), .B2(G137), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT53), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1182), .A2(new_n1185), .B1(G128), .B2(new_n801), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n873), .A2(G132), .B1(new_n1103), .B2(G159), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1181), .A2(new_n1184), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1175), .B1(new_n1178), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1169), .B1(new_n1189), .B2(new_n787), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1138), .A2(new_n1007), .B1(new_n1167), .B2(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1166), .A2(KEYINPUT118), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT118), .B1(new_n1166), .B2(new_n1191), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(G378));
  INV_X1    g0994(.A(KEYINPUT123), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n262), .A2(new_n271), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n969), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT121), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n307), .B2(new_n310), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n307), .A2(new_n310), .A3(new_n1200), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1196), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1203), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1196), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1201), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n971), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n945), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n970), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n960), .B2(new_n961), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1208), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n968), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1209), .A2(new_n1210), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1213), .B1(new_n1212), .B2(new_n968), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1124), .B1(new_n955), .B2(new_n959), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1217), .A2(new_n967), .A3(new_n1211), .A4(new_n1208), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n945), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1158), .A2(new_n1153), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1195), .B1(new_n1220), .B2(KEYINPUT57), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n767), .B1(new_n1220), .B2(KEYINPUT57), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1152), .B1(new_n1226), .B2(new_n1138), .ZN(new_n1227));
  OAI211_X1 g1027(.A(KEYINPUT123), .B(new_n1223), .C1(new_n1225), .C2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1221), .A2(new_n1222), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1224), .A2(new_n1007), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n771), .B1(G50), .B2(new_n1168), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n820), .A2(G137), .B1(G132), .B2(new_n816), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT119), .ZN(new_n1233));
  INV_X1    g1033(.A(G128), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1234), .A2(new_n808), .B1(new_n798), .B2(new_n1179), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G150), .B2(new_n1103), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1233), .B(new_n1236), .C1(new_n1176), .C2(new_n876), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT120), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n822), .A2(G159), .ZN(new_n1242));
  AOI211_X1 g1042(.A(G33), .B(G41), .C1(new_n825), .C2(G124), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n795), .A2(new_n391), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G107), .B2(new_n873), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n1033), .B2(new_n811), .C1(new_n807), .C2(new_n426), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n290), .A2(G41), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1054), .A2(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n831), .A2(new_n536), .B1(new_n876), .B2(new_n530), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(new_n1247), .A2(new_n1025), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT58), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1248), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1253), .B(new_n267), .C1(G33), .C2(G41), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1251), .A2(KEYINPUT58), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1244), .A2(new_n1252), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1231), .B1(new_n1256), .B2(new_n787), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1208), .A2(new_n784), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT122), .B1(new_n1230), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT122), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1259), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n1224), .C2(new_n1007), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1229), .A2(new_n1264), .ZN(G375));
  NOR2_X1   g1065(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1155), .A2(new_n1152), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n979), .A3(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT124), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n374), .B(new_n1245), .C1(G132), .C2(new_n801), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n820), .A2(G150), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G50), .A2(new_n1103), .B1(new_n1180), .B2(new_n816), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n808), .A2(new_n875), .B1(new_n811), .B2(new_n1234), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G159), .B2(new_n824), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n290), .B(new_n1057), .C1(G77), .C2(new_n822), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n820), .A2(G107), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(G116), .A2(new_n816), .B1(new_n801), .B2(G294), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n798), .A2(new_n536), .B1(new_n811), .B2(new_n513), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(G283), .B2(new_n873), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .A4(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1275), .A2(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n787), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n770), .B1(new_n220), .B2(new_n863), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1285), .B(new_n1286), .C1(new_n1131), .C2(new_n785), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n1155), .B2(new_n1008), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1269), .A2(new_n1289), .ZN(G381));
  NAND4_X1  g1090(.A1(new_n1024), .A2(new_n1049), .A3(new_n1090), .A4(new_n1114), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n862), .A2(new_n886), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1166), .A2(new_n1191), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  OR4_X1    g1095(.A1(G375), .A2(new_n1291), .A3(G381), .A4(new_n1295), .ZN(G407));
  NAND2_X1  g1096(.A1(new_n709), .A2(G213), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1293), .A2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G407), .B(G213), .C1(G375), .C2(new_n1299), .ZN(G409));
  NAND3_X1  g1100(.A1(new_n1155), .A2(KEYINPUT60), .A3(new_n1152), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n727), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1266), .A2(KEYINPUT60), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n1267), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1292), .B1(new_n1304), .B2(new_n1288), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1304), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(G384), .A3(new_n1289), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1229), .A2(G378), .A3(new_n1264), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1220), .A2(new_n979), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(new_n1230), .A3(new_n1259), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1293), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1310), .A2(new_n1311), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1311), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1297), .B(new_n1309), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1310), .A2(new_n1314), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(new_n1297), .A3(new_n1309), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1321), .A2(new_n1318), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1023), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1049), .ZN(new_n1325));
  OAI21_X1  g1125(.A(G390), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1291), .A2(new_n1326), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(G393), .B(new_n840), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1328), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1291), .A2(new_n1326), .A3(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1329), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1322), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT127), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1335), .B(new_n1297), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1336));
  INV_X1    g1136(.A(G2897), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1308), .B1(new_n1337), .B2(new_n1297), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1305), .A2(new_n1307), .A3(G2897), .A4(new_n1298), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1336), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1320), .A2(KEYINPUT126), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1310), .A2(new_n1314), .A3(new_n1311), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1335), .B1(new_n1344), .B2(new_n1297), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1319), .B(new_n1334), .C1(new_n1341), .C2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1321), .A2(KEYINPUT62), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1320), .A2(new_n1297), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1340), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1349), .A2(new_n1330), .A3(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1347), .B1(new_n1348), .B2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1346), .A2(new_n1353), .ZN(G405));
  NAND2_X1  g1154(.A1(G375), .A2(new_n1293), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1310), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1309), .ZN(new_n1357));
  XNOR2_X1  g1157(.A(new_n1357), .B(new_n1347), .ZN(G402));
endmodule


