//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1258, new_n1259, new_n1260;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT64), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n449), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT65), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G137), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n469), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(new_n465), .A3(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n462), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR3_X1   g061(.A1(new_n486), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n469), .A2(KEYINPUT66), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n465), .C1(new_n460), .C2(new_n461), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n485), .A2(new_n488), .B1(KEYINPUT4), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n465), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n490), .A2(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n511), .A2(KEYINPUT69), .A3(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n504), .A2(new_n506), .B1(new_n503), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT67), .A3(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(new_n521), .B1(KEYINPUT6), .B2(new_n518), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(G88), .A2(new_n523), .B1(new_n524), .B2(G50), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n514), .A2(new_n515), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G51), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT70), .B(KEYINPUT7), .Z(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(new_n522), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n528), .B(new_n529), .C1(new_n535), .C2(KEYINPUT71), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(KEYINPUT71), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(G168));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n522), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n534), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n518), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n509), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT72), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n551), .A3(G651), .ZN(new_n552));
  AOI22_X1  g127(.A1(G81), .A2(new_n523), .B1(new_n524), .B2(G43), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n516), .A2(new_n522), .A3(G91), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT73), .B(G65), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n516), .A2(new_n562), .B1(G78), .B2(G543), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n563), .B2(new_n518), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n519), .A2(new_n521), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n566), .A2(G53), .A3(G543), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n522), .A2(new_n570), .A3(G53), .A4(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n565), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  OAI21_X1  g150(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n516), .A2(new_n522), .A3(G87), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n522), .A2(G49), .A3(G543), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT74), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n509), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n523), .A2(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n524), .A2(G48), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G305));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n534), .A2(new_n588), .B1(new_n540), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n518), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n590), .A2(new_n592), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G301), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n516), .A2(new_n522), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT75), .Z(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n509), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n524), .B2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n598), .A2(KEYINPUT76), .A3(new_n603), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n595), .B1(new_n608), .B2(new_n594), .ZN(G284));
  AOI21_X1  g184(.A(new_n595), .B1(new_n608), .B2(new_n594), .ZN(G321));
  NAND2_X1  g185(.A1(G299), .A2(new_n594), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G168), .B2(new_n594), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(G168), .B2(new_n594), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n608), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND3_X1  g190(.A1(new_n606), .A2(new_n614), .A3(new_n607), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT77), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT77), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n606), .A2(new_n619), .A3(new_n614), .A4(new_n607), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n618), .A2(new_n594), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n594), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n469), .A2(new_n466), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n475), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n463), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n465), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n630), .A3(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT79), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT78), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2430), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n647), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n628), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n636), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n674), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  AOI211_X1 g253(.A(new_n676), .B(new_n678), .C1(new_n671), .C2(new_n675), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT80), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n681), .A2(new_n683), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n681), .A2(new_n683), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G6), .ZN(new_n693));
  INV_X1    g268(.A(G305), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n692), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(KEYINPUT82), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(KEYINPUT82), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT32), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n695), .A2(KEYINPUT82), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT32), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(new_n701), .A3(new_n696), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n699), .A2(new_n702), .A3(G1981), .ZN(new_n703));
  AOI21_X1  g278(.A(G1981), .B1(new_n699), .B2(new_n702), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n692), .A2(G22), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G303), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT83), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G288), .B2(new_n692), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT84), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n713));
  INV_X1    g288(.A(G1976), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n708), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT34), .B1(new_n705), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n721));
  INV_X1    g296(.A(new_n708), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n713), .A2(new_n715), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G1976), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n722), .B1(new_n724), .B2(new_n716), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT34), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n725), .B(new_n726), .C1(new_n703), .C2(new_n704), .ZN(new_n727));
  NOR2_X1   g302(.A1(G25), .A2(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n475), .A2(G119), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n463), .A2(G131), .ZN(new_n730));
  OR2_X1    g305(.A1(G95), .A2(G2105), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n731), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT81), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n735), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G24), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n590), .A2(new_n592), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n738), .B1(G1986), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G1986), .B2(new_n741), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n720), .A2(new_n721), .A3(new_n727), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT85), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n720), .A2(new_n746), .A3(new_n727), .A4(new_n743), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n745), .A2(KEYINPUT36), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n744), .A2(KEYINPUT85), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n751), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT29), .B(G2090), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n756), .B2(KEYINPUT24), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(KEYINPUT24), .B2(new_n756), .ZN(new_n758));
  INV_X1    g333(.A(G160), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n751), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G11), .ZN(new_n763));
  INV_X1    g338(.A(G28), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(KEYINPUT30), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n751), .B1(new_n766), .B2(G28), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n763), .B1(new_n765), .B2(new_n767), .C1(new_n635), .C2(new_n751), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(new_n465), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n771));
  NAND2_X1  g346(.A1(G103), .A2(G2104), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n463), .A2(G139), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n770), .A2(G29), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G29), .B2(G33), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n762), .A2(new_n768), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G32), .ZN(new_n781));
  AOI21_X1  g356(.A(KEYINPUT92), .B1(new_n751), .B2(new_n781), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n463), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n475), .A2(G129), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT91), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G29), .ZN(new_n789));
  MUX2_X1   g364(.A(KEYINPUT92), .B(new_n782), .S(new_n789), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n755), .B(new_n780), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n751), .A2(G26), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT89), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT28), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n463), .A2(G140), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT87), .Z(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT88), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G128), .B2(new_n475), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2067), .ZN(new_n805));
  INV_X1    g380(.A(G1961), .ZN(new_n806));
  NOR2_X1   g381(.A1(G171), .A2(new_n692), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G5), .B2(new_n692), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n751), .A2(G27), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G164), .B2(new_n751), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G2078), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n777), .A2(new_n778), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT90), .Z(new_n814));
  NOR4_X1   g389(.A1(new_n793), .A2(new_n809), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n692), .A2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G168), .B2(new_n692), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1966), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n692), .A2(G19), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n555), .B2(new_n692), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1341), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n790), .A2(new_n792), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n808), .A2(new_n806), .B1(new_n761), .B2(new_n760), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT93), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n815), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n608), .A2(new_n692), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G4), .B2(new_n692), .ZN(new_n829));
  INV_X1    g404(.A(G1348), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n831), .B(new_n832), .C1(KEYINPUT93), .C2(new_n825), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n692), .A2(G20), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT94), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT23), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G299), .B2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT95), .ZN(new_n838));
  INV_X1    g413(.A(G1956), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n827), .A2(new_n833), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n748), .A2(new_n750), .A3(new_n841), .ZN(G311));
  NAND3_X1  g417(.A1(new_n748), .A2(new_n750), .A3(new_n841), .ZN(G150));
  NAND2_X1  g418(.A1(new_n608), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  INV_X1    g420(.A(G93), .ZN(new_n846));
  INV_X1    g421(.A(G55), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n534), .A2(new_n846), .B1(new_n540), .B2(new_n847), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n518), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n554), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n845), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  INV_X1    g432(.A(new_n851), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(G145));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT96), .B1(new_n494), .B2(new_n497), .ZN(new_n863));
  OR2_X1    g438(.A1(G102), .A2(G2105), .ZN(new_n864));
  INV_X1    g439(.A(G114), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G2105), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n866), .A3(G2104), .ZN(new_n867));
  AND2_X1   g442(.A1(G126), .A2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n460), .B2(new_n461), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n862), .B1(new_n490), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n462), .A2(new_n482), .A3(new_n484), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT66), .B1(new_n469), .B2(new_n487), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n877), .A2(KEYINPUT97), .A3(new_n863), .A4(new_n871), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n788), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n733), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n770), .A2(KEYINPUT98), .A3(new_n775), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n803), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n475), .A2(G130), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n465), .A2(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(G142), .B2(new_n463), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n626), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n883), .B(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n881), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(G160), .B(new_n635), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n480), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n897), .A3(new_n892), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n604), .A2(G299), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n598), .A2(new_n565), .A3(new_n572), .A4(new_n603), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n907), .A2(KEYINPUT41), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n913), .B2(new_n904), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n852), .B1(new_n617), .B2(new_n620), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n617), .A2(new_n620), .A3(new_n852), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n907), .B(KEYINPUT100), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n617), .A2(new_n620), .A3(new_n852), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n920), .B2(new_n915), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(KEYINPUT101), .A3(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(KEYINPUT101), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n925));
  NAND2_X1  g500(.A1(G290), .A2(G288), .ZN(new_n926));
  INV_X1    g501(.A(G288), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n740), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT103), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G166), .A2(G305), .ZN(new_n930));
  NAND2_X1  g505(.A1(G303), .A2(new_n694), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n926), .A2(new_n928), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n930), .B(new_n931), .C1(new_n936), .C2(new_n929), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n925), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n931), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n935), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n926), .A2(KEYINPUT103), .A3(new_n928), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n942), .A2(KEYINPUT42), .A3(new_n932), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n924), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n922), .A2(new_n923), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n922), .B2(new_n923), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n938), .A2(new_n943), .A3(new_n924), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT105), .B1(new_n948), .B2(new_n594), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n950));
  INV_X1    g525(.A(new_n947), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n922), .A2(new_n923), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n944), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n950), .B(G868), .C1(new_n953), .C2(new_n945), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n858), .A2(new_n594), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(G295));
  NAND3_X1  g531(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(G331));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NOR2_X1   g533(.A1(G171), .A2(KEYINPUT106), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n852), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n555), .A2(new_n851), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n554), .A2(new_n858), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G286), .B1(KEYINPUT106), .B2(G171), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n961), .A3(new_n964), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n914), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n942), .A2(new_n932), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n908), .A3(new_n969), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n971), .B2(new_n974), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n958), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n970), .A2(new_n913), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(new_n972), .C1(new_n919), .C2(new_n970), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n981), .A2(KEYINPUT43), .A3(new_n976), .A4(new_n975), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT43), .B1(new_n977), .B2(new_n978), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n981), .A2(new_n958), .A3(new_n976), .A4(new_n975), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(G397));
  OAI21_X1  g565(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n991));
  INV_X1    g566(.A(G40), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n468), .A2(new_n472), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n995));
  OAI211_X1 g570(.A(new_n994), .B(new_n995), .C1(new_n490), .C2(new_n872), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n991), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(KEYINPUT120), .A2(G2084), .ZN(new_n998));
  AND2_X1   g573(.A1(KEYINPUT120), .A2(G2084), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(KEYINPUT45), .B(new_n994), .C1(new_n490), .C2(new_n499), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n470), .A2(new_n471), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1004), .B(G40), .C1(new_n465), .C2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n994), .B1(new_n490), .B2(new_n872), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1003), .B1(new_n1009), .B2(KEYINPUT118), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n870), .B1(new_n867), .B2(new_n869), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n1014), .B2(new_n877), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(KEYINPUT45), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1011), .B1(new_n1016), .B2(new_n1006), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1966), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT119), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT118), .B(new_n993), .C1(new_n1015), .C2(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1002), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT118), .B1(new_n1023), .B2(new_n993), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT119), .B(new_n1019), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(G168), .B(new_n1001), .C1(new_n1020), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(KEYINPUT123), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(KEYINPUT123), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1027), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1001), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(G8), .A3(G286), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1032), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT62), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1019), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g616(.A(G286), .B(new_n1000), .C1(new_n1041), .C2(new_n1025), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1030), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1031), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1035), .A4(new_n1033), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G303), .A2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n873), .A2(new_n878), .A3(KEYINPUT45), .A4(new_n994), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1008), .B1(G164), .B2(G1384), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n993), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1971), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(KEYINPUT110), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT112), .B1(new_n997), .B2(G2090), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1006), .B1(new_n1015), .B2(new_n995), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n1057));
  INV_X1    g632(.A(G2090), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n991), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1054), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT110), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1061));
  OAI211_X1 g636(.A(G8), .B(new_n1049), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT113), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT110), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1066), .A2(new_n1054), .A3(new_n1055), .A4(new_n1059), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(G8), .A4(new_n1049), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1015), .A2(new_n993), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n1028), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n583), .A2(G651), .B1(new_n524), .B2(G48), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n585), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT114), .B(G86), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n523), .A2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT49), .B(new_n1077), .C1(new_n1080), .C2(new_n1076), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT49), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G305), .A2(G1981), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1076), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1074), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n927), .A2(G1976), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1072), .A2(G8), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(G288), .B2(new_n714), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1072), .A2(new_n1090), .A3(G8), .A4(new_n1087), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1071), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1092), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1074), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(KEYINPUT117), .A3(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1097));
  INV_X1    g672(.A(new_n995), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1006), .B1(new_n1007), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n993), .B1(new_n1015), .B2(new_n995), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT116), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1058), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1028), .B1(new_n1104), .B2(new_n1064), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1049), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1093), .A2(new_n1096), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1052), .B2(G2078), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n997), .A2(new_n806), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(G2078), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1110), .B(new_n1111), .C1(new_n1018), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G171), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1070), .A2(new_n1108), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1038), .A2(new_n1046), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1000), .B1(new_n1041), .B2(new_n1025), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1119), .A2(new_n1028), .A3(G286), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1070), .A2(new_n1108), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1067), .A2(G8), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1107), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1086), .A2(new_n1122), .A3(new_n1092), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1070), .A2(new_n1120), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n873), .A2(new_n878), .A3(new_n994), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1113), .B1(new_n1129), .B2(new_n1008), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n993), .A3(new_n1050), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1110), .A2(new_n1111), .A3(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1132), .A2(G171), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT54), .B1(new_n1133), .B2(new_n1115), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  AOI21_X1  g710(.A(G1956), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n569), .A2(new_n571), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n1137), .B2(new_n564), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n572), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n516), .A2(new_n562), .ZN(new_n1141));
  NAND2_X1  g716(.A1(G78), .A2(G543), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G651), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n572), .A3(new_n1145), .A4(new_n561), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1138), .A2(new_n1140), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1140), .B1(new_n1138), .B2(new_n1146), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT56), .B(G2072), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1050), .A2(new_n993), .A3(new_n1051), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1136), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1140), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1138), .A2(new_n1140), .A3(new_n1146), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1100), .B(new_n993), .C1(new_n1015), .C2(new_n995), .ZN(new_n1159));
  OR3_X1    g734(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n839), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1158), .B1(new_n1163), .B2(new_n1151), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1135), .B1(new_n1153), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1149), .B1(new_n1136), .B2(new_n1152), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1163), .A2(new_n1158), .A3(new_n1151), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT61), .ZN(new_n1168));
  INV_X1    g743(.A(G2067), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n997), .A2(new_n830), .B1(new_n1073), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n604), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n598), .A2(KEYINPUT60), .A3(new_n603), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT58), .B(G1341), .Z(new_n1177));
  NAND2_X1  g752(.A1(new_n1072), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1052), .B2(G1996), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n555), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1182), .A3(new_n555), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1165), .A2(new_n1168), .A3(new_n1176), .A4(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1170), .A2(new_n604), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1164), .B1(new_n1167), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1134), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1044), .A2(new_n1035), .A3(new_n1033), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1192), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1132), .A2(G171), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1194), .B(KEYINPUT54), .C1(G171), .C2(new_n1114), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1114), .A2(G171), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1198), .A2(new_n1194), .A3(KEYINPUT124), .A4(KEYINPUT54), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1188), .A2(new_n1189), .A3(new_n1193), .A4(new_n1200), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1070), .A2(new_n1086), .A3(new_n1092), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1203));
  NOR2_X1   g778(.A1(G288), .A2(G1976), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT115), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1077), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1206), .A2(new_n1074), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1118), .A2(new_n1128), .A3(new_n1201), .A4(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1129), .A2(new_n1008), .A3(new_n993), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT107), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1129), .A2(KEYINPUT107), .A3(new_n1008), .A4(new_n993), .ZN(new_n1213));
  INV_X1    g788(.A(G1996), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n788), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT108), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1212), .A2(new_n1215), .A3(KEYINPUT108), .A4(new_n1213), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n803), .B(new_n1169), .ZN(new_n1221));
  INV_X1    g796(.A(new_n788), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1221), .B1(G1996), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1224));
  INV_X1    g799(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  AND3_X1   g801(.A1(new_n1220), .A2(KEYINPUT109), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g802(.A(KEYINPUT109), .B1(new_n1220), .B2(new_n1226), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n733), .B(new_n736), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1229), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g806(.A(G290), .B(G1986), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1231), .B1(new_n1225), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1209), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT46), .ZN(new_n1235));
  OAI211_X1 g810(.A(new_n1221), .B(new_n788), .C1(new_n1235), .C2(G1996), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1225), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1235), .B1(new_n1224), .B2(G1996), .ZN(new_n1238));
  AND2_X1   g813(.A1(new_n1238), .A2(KEYINPUT127), .ZN(new_n1239));
  NOR2_X1   g814(.A1(new_n1238), .A2(KEYINPUT127), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1237), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g816(.A(new_n1241), .B(KEYINPUT47), .ZN(new_n1242));
  NOR3_X1   g817(.A1(new_n1224), .A2(G1986), .A3(G290), .ZN(new_n1243));
  XNOR2_X1  g818(.A(new_n1243), .B(KEYINPUT48), .ZN(new_n1244));
  OAI21_X1  g819(.A(new_n1242), .B1(new_n1231), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n734), .A2(new_n736), .ZN(new_n1246));
  XNOR2_X1  g821(.A(new_n1246), .B(KEYINPUT125), .ZN(new_n1247));
  INV_X1    g822(.A(new_n1247), .ZN(new_n1248));
  NOR3_X1   g823(.A1(new_n1227), .A2(new_n1228), .A3(new_n1248), .ZN(new_n1249));
  NOR2_X1   g824(.A1(new_n803), .A2(G2067), .ZN(new_n1250));
  OAI21_X1  g825(.A(new_n1225), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1251), .A2(KEYINPUT126), .ZN(new_n1252));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1253));
  OAI211_X1 g828(.A(new_n1253), .B(new_n1225), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1254));
  AOI21_X1  g829(.A(new_n1245), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g830(.A1(new_n1234), .A2(new_n1255), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g831(.A(G319), .ZN(new_n1258));
  OR2_X1    g832(.A1(new_n1258), .A2(G227), .ZN(new_n1259));
  NOR3_X1   g833(.A1(G229), .A2(G401), .A3(new_n1259), .ZN(new_n1260));
  AND3_X1   g834(.A1(new_n1260), .A2(new_n987), .A3(new_n902), .ZN(G308));
  NAND3_X1  g835(.A1(new_n1260), .A2(new_n987), .A3(new_n902), .ZN(G225));
endmodule


