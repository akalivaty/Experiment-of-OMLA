//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  INV_X1    g000(.A(G131), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n190), .B2(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n188), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(new_n187), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT65), .A2(G131), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n200), .A2(new_n191), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n194), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(new_n197), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n191), .A3(new_n201), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT66), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n193), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT70), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n212), .A3(G128), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT70), .A4(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n211), .A2(G146), .ZN(new_n221));
  OAI21_X1  g035(.A(G128), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n219), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n215), .A2(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n198), .A2(new_n202), .A3(new_n194), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT66), .B1(new_n204), .B2(new_n205), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n196), .A2(new_n197), .A3(new_n191), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n225), .A2(new_n226), .B1(G131), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n209), .A2(G143), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n229), .B(new_n230), .C1(new_n221), .C2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT0), .A4(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI22_X1  g048(.A1(new_n207), .A2(new_n224), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT72), .A3(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n238), .A2(KEYINPUT71), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n245), .A3(G116), .ZN(new_n246));
  INV_X1    g060(.A(G113), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT2), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G113), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n242), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n242), .B2(new_n246), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n236), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n242), .A2(new_n246), .ZN(new_n255));
  INV_X1    g069(.A(new_n251), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n242), .A2(new_n246), .A3(new_n251), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(KEYINPUT73), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n235), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n232), .A2(new_n263), .A3(new_n233), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n232), .B2(new_n233), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT67), .B1(new_n266), .B2(new_n228), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n232), .A2(new_n263), .A3(new_n233), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n227), .A2(G131), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n203), .B2(new_n206), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n224), .B1(new_n207), .B2(KEYINPUT68), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n192), .B1(new_n225), .B2(new_n226), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT30), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n260), .B1(new_n235), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n262), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(G237), .A2(G953), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G210), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT27), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT26), .B(G101), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n284), .A2(KEYINPUT76), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT76), .B1(new_n284), .B2(new_n290), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n266), .A2(new_n228), .A3(KEYINPUT67), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n273), .B1(new_n270), .B2(new_n272), .ZN(new_n295));
  INV_X1    g109(.A(new_n279), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n215), .A2(new_n220), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n222), .A2(new_n223), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n277), .B2(new_n278), .ZN(new_n300));
  OAI22_X1  g114(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n260), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT28), .B1(new_n235), .B2(new_n260), .ZN(new_n303));
  INV_X1    g117(.A(new_n234), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n304), .A2(new_n272), .B1(new_n299), .B2(new_n277), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n306));
  INV_X1    g120(.A(new_n260), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n293), .B1(new_n310), .B2(new_n290), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n291), .A2(new_n292), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n305), .A2(new_n307), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n303), .B2(new_n308), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n290), .A2(new_n293), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(KEYINPUT77), .A3(new_n315), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G472), .B1(new_n312), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n261), .A2(new_n290), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n324), .B(new_n325), .C1(new_n281), .C2(new_n283), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT75), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n307), .B1(new_n305), .B2(KEYINPUT30), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n267), .A2(new_n274), .B1(new_n276), .B2(new_n279), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(KEYINPUT30), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n325), .A4(new_n324), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n283), .B1(new_n301), .B2(new_n282), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n262), .A2(new_n289), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT31), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT74), .B(KEYINPUT31), .C1(new_n334), .C2(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n310), .A2(new_n290), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n333), .A2(new_n338), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(G472), .A2(G902), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT32), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n339), .A2(new_n340), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n330), .A2(new_n324), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT74), .B1(new_n348), .B2(KEYINPUT31), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n343), .B1(new_n350), .B2(new_n333), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n323), .B(new_n346), .C1(new_n351), .C2(KEYINPUT32), .ZN(new_n352));
  INV_X1    g166(.A(G128), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n238), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT71), .B(G119), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(new_n353), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT24), .B(G110), .Z(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G125), .ZN(new_n360));
  INV_X1    g174(.A(G125), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G140), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n363));
  OR3_X1    g177(.A1(new_n361), .A2(KEYINPUT16), .A3(G140), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G146), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(G146), .B1(new_n363), .B2(new_n364), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n358), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G110), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT23), .B(new_n354), .C1(new_n355), .C2(new_n353), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(new_n355), .B2(G128), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n369), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n356), .A2(new_n357), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n369), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n360), .A2(new_n362), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n378), .A2(KEYINPUT78), .A3(G146), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n380));
  XNOR2_X1  g194(.A(G125), .B(G140), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(new_n209), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n365), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n377), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT22), .B(G137), .ZN(new_n386));
  INV_X1    g200(.A(G953), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(G221), .A3(G234), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n386), .B(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n374), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n368), .A2(new_n373), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n383), .B1(new_n375), .B2(new_n376), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n394), .A3(new_n321), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT25), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n390), .A2(new_n394), .A3(KEYINPUT25), .A4(new_n321), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G217), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(G234), .B2(new_n321), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(KEYINPUT79), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT79), .B1(new_n399), .B2(new_n401), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n390), .A2(new_n394), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n401), .A2(G902), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n407), .B(KEYINPUT80), .Z(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT81), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT9), .B(G234), .ZN(new_n413));
  OAI21_X1  g227(.A(G221), .B1(new_n413), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G469), .ZN(new_n416));
  XNOR2_X1  g230(.A(G104), .B(G107), .ZN(new_n417));
  INV_X1    g231(.A(G101), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT83), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT82), .B(G101), .ZN(new_n420));
  INV_X1    g234(.A(G104), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT3), .B1(new_n421), .B2(G107), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(G107), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n424));
  INV_X1    g238(.A(G107), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(G104), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n420), .A2(new_n422), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n421), .A2(G107), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n425), .A2(G104), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n428), .B(G101), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n419), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(new_n297), .A3(new_n298), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n219), .B2(G128), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n215), .B2(new_n220), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(new_n432), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n272), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT12), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n439), .A2(KEYINPUT84), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(KEYINPUT84), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G110), .B(G140), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n387), .A2(G227), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n432), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n299), .A2(new_n447), .A3(KEYINPUT10), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT10), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n436), .B2(new_n432), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n427), .A2(KEYINPUT4), .B1(G101), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(KEYINPUT4), .A3(G101), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n304), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n448), .A2(new_n450), .A3(new_n228), .A4(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n432), .A2(new_n297), .A3(new_n298), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n432), .B2(new_n436), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n458), .A2(KEYINPUT84), .A3(new_n439), .A4(new_n272), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n442), .A2(new_n446), .A3(new_n456), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n448), .A2(new_n455), .A3(new_n450), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n272), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n446), .B1(new_n462), .B2(new_n456), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n460), .B1(new_n463), .B2(KEYINPUT85), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n465), .B(new_n446), .C1(new_n462), .C2(new_n456), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n416), .B(new_n321), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n416), .A2(new_n321), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n442), .A2(new_n456), .A3(new_n459), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n456), .A2(new_n446), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n469), .A2(new_n445), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n468), .B1(new_n471), .B2(G469), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n415), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT86), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n352), .A2(new_n412), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n432), .A2(new_n252), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n255), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n477), .ZN(new_n479));
  OAI21_X1  g293(.A(G113), .B1(new_n479), .B2(new_n246), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT89), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT89), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n476), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT82), .B(G101), .Z(new_n486));
  OAI21_X1  g300(.A(KEYINPUT4), .B1(new_n451), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n451), .A2(G101), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI221_X4 g303(.A(new_n485), .B1(new_n489), .B2(new_n453), .C1(new_n254), .C2(new_n259), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n453), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT87), .B1(new_n260), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n484), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G110), .B(G122), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n494), .B(new_n484), .C1(new_n490), .C2(new_n492), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(KEYINPUT6), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n499), .A3(new_n495), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n224), .A2(new_n361), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n234), .A2(G125), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G224), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(G953), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n503), .B(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n498), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n508), .A2(KEYINPUT91), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n501), .A2(new_n502), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n508), .B2(new_n505), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n505), .A2(new_n508), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n501), .A2(new_n502), .A3(new_n512), .A4(new_n509), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n242), .A2(new_n246), .A3(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n476), .B1(new_n480), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n483), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n252), .B1(new_n517), .B2(new_n481), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n518), .B2(new_n447), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n494), .B(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n514), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(G902), .B1(new_n522), .B2(new_n497), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n507), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT92), .ZN(new_n525));
  OAI21_X1  g339(.A(G210), .B1(G237), .B2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n507), .A2(new_n528), .A3(new_n523), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n507), .A2(new_n523), .A3(new_n526), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G214), .B1(G237), .B2(G902), .ZN(new_n533));
  AND2_X1   g347(.A1(KEYINPUT65), .A2(G131), .ZN(new_n534));
  NOR2_X1   g348(.A1(KEYINPUT65), .A2(G131), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n285), .A2(G143), .A3(G214), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G143), .B1(new_n285), .B2(G214), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G237), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n387), .A3(G214), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n211), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n538), .A3(new_n536), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(KEYINPUT94), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n544), .A2(new_n547), .A3(new_n536), .A4(new_n538), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n537), .B(KEYINPUT17), .C1(new_n539), .C2(new_n540), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n553), .A2(new_n367), .A3(new_n366), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G113), .B(G122), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(new_n421), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT18), .B(G131), .C1(new_n539), .C2(new_n540), .ZN(new_n558));
  NAND2_X1  g372(.A1(KEYINPUT18), .A2(G131), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n544), .A2(new_n538), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT78), .B1(new_n378), .B2(G146), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n381), .A2(new_n380), .A3(new_n209), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n562), .A2(new_n563), .B1(G146), .B2(new_n378), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT93), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n379), .A2(new_n382), .B1(new_n209), .B2(new_n381), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n560), .A4(new_n558), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n555), .A2(new_n557), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n557), .B1(new_n555), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n321), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G475), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT20), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n378), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n381), .A2(KEYINPUT19), .ZN(new_n577));
  AOI21_X1  g391(.A(G146), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n366), .B1(new_n578), .B2(KEYINPUT95), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n548), .A4(new_n546), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n569), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n557), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n555), .A2(new_n557), .A3(new_n569), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(G475), .A2(G902), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n574), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n587), .ZN(new_n589));
  AOI211_X1 g403(.A(KEYINPUT20), .B(new_n589), .C1(new_n584), .C2(new_n585), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n573), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n387), .A2(G952), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(G234), .B2(G237), .ZN(new_n594));
  NAND2_X1  g408(.A1(G234), .A2(G237), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(G902), .A3(G953), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT21), .B(G898), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G478), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n211), .A2(G128), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n353), .A2(G143), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(G128), .B(G143), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n190), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n606), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n612), .A3(G134), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G122), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G116), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n240), .A2(G122), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(G107), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT97), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n617), .A2(new_n621), .A3(KEYINPUT14), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n617), .B2(KEYINPUT14), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n616), .B1(new_n617), .B2(KEYINPUT14), .ZN(new_n626));
  OAI21_X1  g440(.A(G107), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n614), .A2(new_n620), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n608), .A2(KEYINPUT13), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n629), .B(G134), .C1(KEYINPUT13), .C2(new_n603), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n425), .B1(new_n616), .B2(new_n617), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n610), .B(new_n630), .C1(new_n631), .C2(new_n619), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n413), .A2(new_n400), .A3(G953), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n628), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n628), .B2(new_n632), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n321), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n602), .B1(new_n636), .B2(KEYINPUT99), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(KEYINPUT99), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n639), .B(new_n321), .C1(new_n634), .C2(new_n635), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n637), .B1(new_n641), .B2(new_n602), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n592), .A2(new_n600), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n532), .A2(new_n533), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n475), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n420), .ZN(G3));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n327), .A2(new_n332), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n321), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(G472), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n467), .A2(new_n472), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n414), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT86), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n341), .A2(new_n342), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT86), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n473), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n652), .A2(new_n655), .A3(new_n656), .A4(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n648), .B1(new_n659), .B2(new_n411), .ZN(new_n660));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n341), .B2(new_n321), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n351), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n474), .A2(new_n663), .A3(KEYINPUT100), .A4(new_n412), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n507), .A2(new_n523), .A3(new_n526), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n526), .B1(new_n507), .B2(new_n523), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n533), .B(new_n600), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n601), .A2(G902), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT33), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT33), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n628), .A2(new_n632), .ZN(new_n672));
  INV_X1    g486(.A(new_n633), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n628), .A2(new_n632), .A3(new_n633), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n669), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n636), .A2(new_n678), .A3(new_n601), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n636), .B2(new_n601), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n591), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n668), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n665), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT34), .B(G104), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G6));
  NOR2_X1   g500(.A1(new_n642), .A2(new_n591), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n668), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n665), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  NAND2_X1  g506(.A1(new_n399), .A2(new_n401), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT79), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n374), .A2(new_n385), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n391), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n408), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n695), .A2(new_n402), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n532), .A2(new_n533), .A3(new_n644), .A4(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n659), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT37), .B(G110), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G12));
  OAI21_X1  g518(.A(new_n533), .B1(new_n666), .B2(new_n667), .ZN(new_n705));
  INV_X1    g519(.A(new_n594), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n596), .A2(G900), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n687), .A2(new_n700), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n352), .A2(new_n710), .A3(new_n474), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G128), .ZN(G30));
  INV_X1    g526(.A(new_n474), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n708), .B(KEYINPUT39), .Z(new_n714));
  OR3_X1    g528(.A1(new_n713), .A2(KEYINPUT40), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT40), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n532), .B(KEYINPUT38), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n284), .A2(new_n289), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n313), .A2(new_n261), .A3(new_n289), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(G902), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n661), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n346), .B(new_n722), .C1(new_n351), .C2(KEYINPUT32), .ZN(new_n723));
  INV_X1    g537(.A(new_n700), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n588), .A2(new_n590), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n642), .B1(new_n725), .B2(new_n573), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n533), .A2(new_n723), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  AND3_X1   g543(.A1(new_n591), .A2(new_n681), .A3(new_n708), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT102), .B1(new_n705), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n533), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n524), .A2(new_n527), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n734), .B2(new_n531), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT102), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n730), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n352), .A3(new_n474), .A4(new_n700), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  OAI21_X1  g554(.A(new_n321), .B1(new_n464), .B2(new_n466), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n414), .A3(new_n467), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n683), .A2(new_n352), .A3(new_n412), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  NAND4_X1  g561(.A1(new_n689), .A2(new_n352), .A3(new_n412), .A4(new_n744), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT103), .B(G116), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G18));
  NOR2_X1   g564(.A1(new_n705), .A2(new_n743), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n352), .A2(new_n751), .A3(new_n644), .A4(new_n700), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  XNOR2_X1  g567(.A(new_n342), .B(KEYINPUT104), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n314), .A2(new_n289), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(KEYINPUT31), .B2(new_n348), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n755), .B1(new_n333), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n662), .A2(new_n411), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n668), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n743), .A2(new_n592), .A3(new_n642), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NOR3_X1   g577(.A1(new_n705), .A2(new_n731), .A3(new_n743), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n662), .A2(new_n724), .A3(new_n758), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  NOR2_X1   g581(.A1(new_n666), .A2(new_n733), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n530), .A2(new_n473), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n352), .A3(new_n412), .A4(new_n730), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n530), .A2(new_n768), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n654), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT105), .B1(new_n351), .B2(KEYINPUT32), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT105), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n656), .A2(new_n777), .A3(new_n344), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n776), .A2(new_n346), .A3(new_n778), .A4(new_n323), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(new_n779), .A3(new_n412), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  INV_X1    g596(.A(new_n708), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n688), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n769), .A2(new_n352), .A3(new_n412), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  NAND3_X1  g600(.A1(new_n592), .A2(KEYINPUT43), .A3(new_n681), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT106), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n591), .B1(new_n788), .B2(new_n681), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n788), .B2(new_n681), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT43), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n790), .A2(KEYINPUT107), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT107), .B1(new_n790), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n663), .A2(new_n724), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n773), .B1(new_n797), .B2(KEYINPUT44), .ZN(new_n798));
  INV_X1    g612(.A(new_n467), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n471), .A2(KEYINPUT45), .ZN(new_n800));
  OAI21_X1  g614(.A(G469), .B1(new_n471), .B2(KEYINPUT45), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n800), .A2(new_n801), .B1(new_n416), .B2(new_n321), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT46), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n803), .B2(new_n802), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n414), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n714), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n796), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n798), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  XOR2_X1   g624(.A(KEYINPUT108), .B(G137), .Z(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(G39));
  AND3_X1   g626(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n414), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT47), .B1(new_n805), .B2(new_n414), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n352), .ZN(new_n816));
  INV_X1    g630(.A(new_n773), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n411), .A3(new_n730), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(new_n359), .ZN(G42));
  AND3_X1   g634(.A1(new_n794), .A2(new_n594), .A3(new_n759), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n751), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT116), .ZN(new_n823));
  INV_X1    g637(.A(new_n723), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n773), .A2(new_n743), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n594), .A4(new_n412), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n826), .A2(KEYINPUT114), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(KEYINPUT114), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n682), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n593), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n794), .A2(new_n594), .A3(new_n825), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT48), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n777), .B1(new_n656), .B2(new_n344), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n323), .A2(new_n346), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n411), .B1(new_n837), .B2(new_n778), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n833), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n834), .B1(new_n833), .B2(new_n838), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n823), .B(new_n831), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n717), .A2(new_n533), .A3(new_n743), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n821), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT50), .ZN(new_n844));
  INV_X1    g658(.A(new_n681), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n827), .A2(new_n592), .A3(new_n845), .A4(new_n828), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n833), .A2(new_n765), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n821), .A2(new_n842), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n844), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n815), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n742), .A2(new_n467), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n414), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n821), .A2(new_n817), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT51), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n841), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n851), .A2(KEYINPUT113), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n853), .B1(new_n851), .B2(KEYINPUT113), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n855), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n859), .B1(new_n850), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(KEYINPUT115), .B(new_n859), .C1(new_n850), .C2(new_n862), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n726), .B(new_n533), .C1(new_n666), .C2(new_n667), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n654), .A2(new_n700), .A3(new_n783), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n723), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n352), .A2(new_n474), .A3(new_n700), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n876), .B2(new_n738), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n352), .A2(new_n474), .A3(new_n710), .ZN(new_n878));
  INV_X1    g692(.A(new_n758), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n652), .A2(new_n700), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n735), .A2(new_n744), .A3(new_n730), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT109), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT109), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n766), .A2(new_n711), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n877), .A2(new_n883), .A3(KEYINPUT52), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n723), .A2(new_n872), .A3(new_n873), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n732), .A2(new_n737), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n875), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n766), .A2(new_n711), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n870), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n870), .A3(new_n892), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n745), .A2(new_n748), .A3(new_n752), .A4(new_n762), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n772), .B2(new_n780), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n475), .A2(new_n645), .B1(new_n701), .B2(new_n659), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n688), .A2(new_n682), .ZN(new_n900));
  AND4_X1   g714(.A1(new_n533), .A2(new_n532), .A3(new_n600), .A4(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n665), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n592), .A2(new_n642), .A3(new_n708), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n530), .A2(new_n768), .A3(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(new_n352), .A3(new_n474), .A4(new_n700), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n769), .A2(new_n765), .A3(new_n730), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n785), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n898), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n908), .A2(KEYINPUT53), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT111), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n766), .A2(new_n711), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(KEYINPUT52), .A3(new_n739), .A4(new_n888), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n892), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n745), .A2(new_n748), .A3(new_n752), .A4(new_n762), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(new_n781), .A3(new_n907), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n352), .A2(new_n412), .A3(new_n474), .ZN(new_n917));
  INV_X1    g731(.A(new_n645), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n526), .B1(new_n524), .B2(KEYINPUT92), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n666), .B1(new_n919), .B2(new_n529), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n920), .A2(new_n733), .A3(new_n643), .A4(new_n724), .ZN(new_n921));
  INV_X1    g735(.A(new_n659), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n917), .A2(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n660), .A2(new_n901), .A3(new_n664), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n892), .A2(new_n912), .A3(new_n910), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n914), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n896), .A2(new_n909), .B1(new_n928), .B2(KEYINPUT53), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n907), .A2(new_n923), .A3(KEYINPUT53), .A4(new_n924), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT112), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n838), .A2(new_n775), .B1(new_n770), .B2(new_n771), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n897), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n915), .A2(new_n781), .A3(KEYINPUT112), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n886), .A2(new_n870), .A3(new_n892), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n893), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT53), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n928), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g756(.A1(KEYINPUT54), .A2(new_n929), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n869), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n867), .A2(new_n868), .ZN(new_n945));
  OAI22_X1  g759(.A1(new_n944), .A2(new_n945), .B1(G952), .B2(G953), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n845), .A2(new_n733), .A3(new_n415), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n412), .A2(new_n947), .A3(new_n592), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n852), .A2(KEYINPUT49), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(KEYINPUT49), .B2(new_n852), .ZN(new_n951));
  OR3_X1    g765(.A1(new_n951), .A2(new_n717), .A3(new_n723), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n946), .A2(new_n952), .ZN(G75));
  NOR2_X1   g767(.A1(new_n908), .A2(new_n913), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT53), .B1(new_n954), .B2(new_n927), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n785), .A2(new_n905), .A3(new_n906), .A4(KEYINPUT53), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n925), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n932), .A2(new_n931), .A3(new_n897), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT112), .B1(new_n915), .B2(new_n781), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n895), .B2(new_n894), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n321), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT56), .B1(new_n963), .B2(G210), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n498), .A2(new_n500), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT118), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n506), .B(KEYINPUT55), .Z(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n387), .A2(G952), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n964), .B2(new_n968), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n969), .A2(new_n972), .ZN(G51));
  OAI21_X1  g787(.A(KEYINPUT119), .B1(new_n939), .B2(new_n955), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT54), .B1(new_n955), .B2(new_n961), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT119), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n942), .A2(new_n976), .A3(new_n938), .A4(new_n937), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n468), .B(KEYINPUT57), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n466), .B2(new_n464), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n800), .A2(new_n801), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n963), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n970), .B1(new_n981), .B2(new_n983), .ZN(G54));
  AND2_X1   g798(.A1(KEYINPUT58), .A2(G475), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n963), .A2(new_n586), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n586), .B1(new_n963), .B2(new_n985), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n986), .A2(new_n987), .A3(new_n970), .ZN(G60));
  OR2_X1    g802(.A1(new_n670), .A2(new_n676), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n991));
  NAND2_X1  g805(.A1(G478), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n990), .B1(new_n943), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n990), .A2(new_n993), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n970), .B1(new_n978), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT121), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI211_X1 g812(.A(KEYINPUT121), .B(new_n970), .C1(new_n978), .C2(new_n995), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(G63));
  XNOR2_X1  g814(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G217), .A2(G902), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n962), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n698), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1005), .B(new_n971), .C1(new_n406), .C2(new_n1004), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1004), .A2(new_n406), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1009), .A2(KEYINPUT61), .A3(new_n971), .A4(new_n1005), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(G66));
  OAI21_X1  g825(.A(G953), .B1(new_n598), .B2(new_n504), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT123), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n925), .A2(new_n897), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1013), .B1(new_n1014), .B2(G953), .ZN(new_n1015));
  INV_X1    g829(.A(new_n966), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1016), .B1(G898), .B2(new_n387), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1015), .B(new_n1017), .ZN(G69));
  AOI21_X1  g832(.A(new_n387), .B1(G227), .B2(G900), .ZN(new_n1019));
  INV_X1    g833(.A(new_n819), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n810), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n883), .A2(new_n739), .A3(new_n885), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n807), .A2(new_n838), .A3(new_n872), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n781), .A2(new_n1023), .A3(new_n785), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n387), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n281), .B1(KEYINPUT30), .B2(new_n305), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n576), .A2(new_n577), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(G900), .A2(G953), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1019), .B1(new_n1031), .B2(KEYINPUT125), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n816), .A2(new_n411), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n900), .B(KEYINPUT124), .Z(new_n1034));
  NOR2_X1   g848(.A1(new_n713), .A2(new_n714), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n817), .ZN(new_n1036));
  AND3_X1   g850(.A1(new_n810), .A2(new_n1020), .A3(new_n1036), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n728), .A2(new_n883), .A3(new_n739), .A4(new_n885), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AND2_X1   g855(.A1(new_n1041), .A2(new_n387), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1031), .B1(new_n1042), .B2(new_n1029), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1032), .B(new_n1043), .Z(G72));
  NAND4_X1  g858(.A1(new_n1037), .A2(new_n1039), .A3(new_n1014), .A4(new_n1040), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  NAND3_X1  g861(.A1(new_n1045), .A2(KEYINPUT126), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n718), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT127), .ZN(new_n1051));
  AOI21_X1  g865(.A(KEYINPUT126), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1052));
  OR3_X1    g866(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1051), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1054));
  INV_X1    g868(.A(new_n1047), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1055), .B1(new_n1025), .B2(new_n1014), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n330), .A2(new_n262), .A3(new_n290), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n971), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n291), .A2(new_n292), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1055), .B1(new_n1059), .B2(new_n348), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n1058), .B1(new_n929), .B2(new_n1060), .ZN(new_n1061));
  AND3_X1   g875(.A1(new_n1053), .A2(new_n1054), .A3(new_n1061), .ZN(G57));
endmodule


