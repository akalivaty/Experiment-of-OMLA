//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n597,
    new_n598, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n458), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n458), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(new_n468), .ZN(G160));
  NOR2_X1   g044(.A1(new_n463), .A2(new_n464), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G136), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n458), .A2(G112), .ZN(new_n473));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n476), .B1(new_n470), .B2(new_n458), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n459), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n475), .B1(G124), .B2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT68), .Z(G162));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n483));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n484), .A2(new_n486), .A3(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n463), .B2(new_n464), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n490), .B(new_n493), .C1(new_n464), .C2(new_n463), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n488), .B1(new_n492), .B2(new_n494), .ZN(G164));
  OR2_X1    g070(.A1(KEYINPUT5), .A2(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT69), .B(G88), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n501), .A2(new_n507), .ZN(G303));
  INV_X1    g083(.A(G303), .ZN(G166));
  INV_X1    g084(.A(new_n498), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n502), .A2(G89), .ZN(new_n511));
  NAND2_X1  g086(.A1(G63), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT70), .B(G51), .Z(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n505), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n513), .A2(new_n517), .ZN(G168));
  AOI22_X1  g093(.A1(new_n498), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n500), .ZN(new_n520));
  INV_X1    g095(.A(G90), .ZN(new_n521));
  INV_X1    g096(.A(G52), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n503), .A2(new_n521), .B1(new_n505), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n520), .A2(new_n523), .ZN(G301));
  INV_X1    g099(.A(G301), .ZN(G171));
  AOI22_X1  g100(.A1(new_n498), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n500), .ZN(new_n527));
  INV_X1    g102(.A(G81), .ZN(new_n528));
  INV_X1    g103(.A(G43), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n503), .A2(new_n528), .B1(new_n505), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n532), .B1(new_n505), .B2(new_n529), .C1(new_n528), .C2(new_n503), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n527), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND4_X1  g114(.A1(G319), .A2(G483), .A3(G661), .A4(new_n539), .ZN(G188));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  INV_X1    g116(.A(G53), .ZN(new_n542));
  NOR3_X1   g117(.A1(new_n505), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT9), .ZN(new_n544));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(KEYINPUT6), .A2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(KEYINPUT6), .A2(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT73), .B1(new_n548), .B2(G53), .ZN(new_n549));
  NOR3_X1   g124(.A1(new_n543), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n503), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G91), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n541), .B(new_n544), .C1(new_n505), .C2(new_n542), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n496), .B2(new_n497), .ZN(new_n555));
  AND2_X1   g130(.A1(G78), .A2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n552), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  OR2_X1    g136(.A1(new_n498), .A2(G74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(G49), .B2(new_n548), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n551), .B2(G87), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n503), .A2(KEYINPUT74), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(G288));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n496), .B2(new_n497), .ZN(new_n570));
  AND2_X1   g145(.A1(G73), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n498), .A2(new_n502), .A3(G86), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n548), .A2(G48), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT75), .ZN(G305));
  AOI22_X1  g151(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n500), .ZN(new_n578));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n503), .A2(new_n579), .B1(new_n505), .B2(new_n580), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n578), .A2(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n498), .A2(new_n502), .A3(G92), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n548), .A2(G54), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n498), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n500), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n583), .B1(new_n591), .B2(G868), .ZN(G284));
  OAI21_X1  g167(.A(new_n583), .B1(new_n591), .B2(G868), .ZN(G321));
  NAND2_X1  g168(.A1(G286), .A2(G868), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n559), .B2(G868), .ZN(G297));
  OAI21_X1  g170(.A(new_n594), .B1(new_n559), .B2(G868), .ZN(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n591), .B1(new_n597), .B2(G860), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT76), .ZN(G148));
  NAND2_X1  g174(.A1(new_n591), .A2(new_n597), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G868), .B2(new_n534), .ZN(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g178(.A1(new_n459), .A2(new_n466), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT78), .ZN(new_n605));
  XNOR2_X1  g180(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(G2100), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n471), .A2(G135), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n458), .A2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  INV_X1    g189(.A(G123), .ZN(new_n615));
  OAI221_X1 g190(.A(new_n612), .B1(new_n613), .B2(new_n614), .C1(new_n479), .C2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT80), .B(G2096), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n610), .A2(new_n611), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT81), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT82), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n627), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(new_n635), .A3(G14), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  INV_X1    g212(.A(KEYINPUT18), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2096), .B(G2100), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n641), .B2(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT83), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(G227));
  XNOR2_X1  g225(.A(G1961), .B(G1966), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n652), .A2(new_n654), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n661), .A2(new_n657), .A3(new_n655), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n659), .B(new_n662), .C1(new_n657), .C2(new_n661), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT85), .Z(new_n664));
  XOR2_X1   g239(.A(G1981), .B(G1986), .Z(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n664), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G229));
  MUX2_X1   g246(.A(G6), .B(G305), .S(G16), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT32), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G288), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n676), .B2(G23), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT33), .B(G1976), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n676), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(G1971), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(G1971), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n674), .A2(new_n681), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT34), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n480), .A2(G119), .ZN(new_n694));
  OAI21_X1  g269(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n695));
  INV_X1    g270(.A(G107), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G2105), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n471), .B2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n693), .B1(new_n700), .B2(new_n692), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(KEYINPUT86), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(KEYINPUT86), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n676), .A2(G24), .ZN(new_n707));
  INV_X1    g282(.A(G290), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n676), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n690), .A2(new_n691), .A3(new_n705), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT36), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n692), .A2(G35), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G162), .B2(new_n692), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2090), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n692), .A2(G26), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT28), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n471), .A2(G140), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n458), .A2(G116), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n723));
  INV_X1    g298(.A(G128), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n721), .B1(new_n722), .B2(new_n723), .C1(new_n479), .C2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G2067), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n692), .A2(G33), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n471), .A2(G139), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n459), .A2(G127), .ZN(new_n736));
  NAND2_X1  g311(.A1(G115), .A2(G2104), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n458), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT87), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n729), .B1(new_n740), .B2(new_n692), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2072), .ZN(new_n742));
  INV_X1    g317(.A(G1341), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n534), .A2(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G16), .B2(G19), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n742), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n728), .B(new_n746), .C1(new_n743), .C2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n480), .A2(G129), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n466), .A2(G105), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT26), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n749), .B(new_n751), .C1(G141), .C2(new_n471), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(new_n692), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n692), .B2(G32), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n676), .A2(G4), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n591), .B2(new_n676), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n756), .A2(new_n757), .B1(G1348), .B2(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(G1348), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n760), .B(new_n761), .C1(new_n756), .C2(new_n757), .ZN(new_n762));
  NOR2_X1   g337(.A1(G168), .A2(new_n676), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n676), .B2(G21), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G160), .A2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G34), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(KEYINPUT24), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n767), .B2(KEYINPUT24), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(KEYINPUT88), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(KEYINPUT88), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n765), .A2(G1966), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n616), .A2(new_n692), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT89), .Z(new_n776));
  NOR2_X1   g351(.A1(G5), .A2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT90), .Z(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G301), .B2(new_n676), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1961), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n781), .A2(G28), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n692), .B1(new_n781), .B2(G28), .ZN(new_n783));
  AND2_X1   g358(.A1(KEYINPUT31), .A2(G11), .ZN(new_n784));
  NOR2_X1   g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  OAI22_X1  g360(.A1(new_n782), .A2(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G1966), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n764), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n774), .A2(new_n776), .A3(new_n780), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G27), .A2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G164), .B2(G29), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT91), .B(G2078), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n793), .B1(new_n773), .B2(new_n772), .C1(new_n741), .C2(G2072), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n676), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT93), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT23), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G299), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1956), .Z(new_n799));
  NOR4_X1   g374(.A1(new_n762), .A2(new_n789), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n718), .A2(new_n747), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n713), .A2(new_n801), .ZN(G150));
  INV_X1    g377(.A(G150), .ZN(G311));
  NAND2_X1  g378(.A1(new_n548), .A2(G55), .ZN(new_n804));
  INV_X1    g379(.A(G93), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n498), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n804), .B1(new_n503), .B2(new_n805), .C1(new_n806), .C2(new_n500), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT94), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G860), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT97), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n534), .A2(new_n807), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n808), .B2(new_n534), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT95), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(new_n813), .C1(new_n808), .C2(new_n534), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n597), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n818), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n823), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n812), .B1(new_n824), .B2(new_n826), .ZN(G145));
  XNOR2_X1  g402(.A(new_n616), .B(G160), .ZN(new_n828));
  XNOR2_X1  g403(.A(G162), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n699), .B(KEYINPUT100), .ZN(new_n831));
  INV_X1    g406(.A(new_n607), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n480), .A2(G130), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT99), .Z(new_n836));
  OR2_X1    g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n471), .A2(G142), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n831), .A2(new_n832), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n834), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n842), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n831), .A2(new_n832), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n833), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n830), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n842), .B1(new_n834), .B2(new_n843), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n845), .A3(new_n833), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n849), .A2(KEYINPUT101), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n753), .B(new_n725), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n492), .A2(new_n494), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n483), .A2(new_n487), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n856), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n857), .B(new_n858), .C1(new_n738), .C2(new_n735), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n853), .A2(new_n856), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n740), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n829), .B1(new_n852), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(KEYINPUT102), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n849), .A2(new_n850), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n859), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n852), .A2(new_n864), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n863), .B1(new_n851), .B2(new_n848), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n829), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g451(.A(new_n818), .B(new_n600), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n591), .A2(G299), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n819), .A2(new_n559), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT103), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n819), .A2(new_n559), .A3(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT104), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n877), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n878), .A2(new_n879), .A3(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n877), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G305), .B(G288), .ZN(new_n893));
  XNOR2_X1  g468(.A(G303), .B(G290), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n888), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n888), .B2(new_n892), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n901));
  INV_X1    g476(.A(G868), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n808), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(G295));
  NAND2_X1  g481(.A1(new_n900), .A2(new_n903), .ZN(G331));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n891), .B1(new_n883), .B2(KEYINPUT41), .ZN(new_n909));
  XNOR2_X1  g484(.A(G301), .B(G168), .ZN(new_n910));
  INV_X1    g485(.A(new_n817), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n531), .A2(new_n533), .ZN(new_n912));
  INV_X1    g487(.A(new_n527), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n807), .A2(KEYINPUT94), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n807), .A2(KEYINPUT94), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n816), .B1(new_n917), .B2(new_n813), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n910), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  INV_X1    g495(.A(new_n910), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n815), .A2(new_n817), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n815), .A2(KEYINPUT106), .A3(new_n817), .A4(new_n921), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n909), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(KEYINPUT107), .A3(new_n922), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n815), .A2(new_n927), .A3(new_n817), .A4(new_n921), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n882), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G37), .B1(new_n930), .B2(new_n895), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(new_n895), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n889), .B1(new_n878), .B2(new_n879), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n882), .B2(new_n889), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n926), .A2(new_n936), .A3(new_n928), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n923), .A2(new_n924), .B1(new_n884), .B2(new_n886), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n934), .B1(new_n925), .B2(new_n929), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n933), .B1(new_n931), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n909), .A2(new_n923), .A3(new_n924), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n926), .A2(new_n928), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n895), .B(new_n943), .C1(new_n944), .C2(new_n882), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n939), .A2(new_n945), .A3(new_n933), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT108), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n908), .B(new_n940), .C1(new_n942), .C2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT43), .B1(new_n931), .B2(new_n941), .ZN(new_n950));
  AND4_X1   g525(.A1(KEYINPUT43), .A2(new_n939), .A3(new_n945), .A4(new_n946), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G164), .B2(G1384), .ZN(new_n955));
  INV_X1    g530(.A(G125), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n470), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n461), .ZN(new_n958));
  OAI21_X1  g533(.A(G2105), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n468), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(G40), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n725), .B(new_n727), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n754), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n963), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT46), .B1(new_n963), .B2(G1996), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n753), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n700), .A2(new_n702), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n699), .A2(new_n703), .ZN(new_n973));
  AND4_X1   g548(.A1(new_n964), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(new_n963), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT126), .ZN(new_n976));
  INV_X1    g551(.A(G1986), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n962), .A2(new_n977), .A3(new_n708), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT48), .Z(new_n979));
  NOR2_X1   g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n971), .A2(new_n964), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n981), .A2(new_n972), .B1(G2067), .B2(new_n725), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n969), .B(new_n980), .C1(new_n962), .C2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n462), .A2(new_n984), .A3(new_n468), .ZN(new_n985));
  AOI21_X1  g560(.A(G1384), .B1(new_n854), .B2(new_n855), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(KEYINPUT45), .ZN(new_n987));
  NOR3_X1   g562(.A1(G164), .A2(new_n954), .A3(G1384), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n787), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n856), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n990), .A2(new_n993), .A3(new_n773), .A4(new_n985), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(G8), .A3(G286), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n989), .B2(new_n994), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(KEYINPUT120), .A3(G286), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n1003));
  AOI22_X1  g578(.A1(G286), .A2(G8), .B1(new_n1003), .B2(KEYINPUT51), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(KEYINPUT51), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n990), .A2(new_n993), .A3(new_n985), .ZN(new_n1006));
  INV_X1    g581(.A(new_n494), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n493), .B1(new_n459), .B2(new_n490), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT45), .B(new_n992), .C1(new_n1009), .C2(new_n488), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n955), .A2(new_n985), .A3(new_n1010), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1006), .A2(new_n773), .B1(new_n1011), .B2(new_n787), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1004), .B(new_n1005), .C1(new_n1012), .C2(new_n999), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1005), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1004), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1000), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT122), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1002), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1002), .B2(new_n1017), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT62), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1002), .A2(new_n1017), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT122), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT62), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1002), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n999), .B1(new_n985), .B2(new_n986), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1028), .B(new_n1029), .C1(new_n1027), .C2(G288), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1029), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G288), .A2(new_n1027), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n574), .A2(new_n573), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n572), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n572), .A2(new_n1036), .A3(new_n573), .A4(new_n574), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT112), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n572), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1037), .A2(new_n1039), .B1(new_n1040), .B2(G1981), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1029), .B1(new_n1041), .B2(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(G1981), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1030), .B(new_n1033), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1971), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT109), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n856), .A2(new_n1048), .A3(KEYINPUT45), .A4(new_n992), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(new_n955), .A3(new_n985), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n986), .B2(KEYINPUT45), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT111), .B(G2090), .Z(new_n1053));
  NAND2_X1  g628(.A1(new_n1006), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT55), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1046), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(KEYINPUT110), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(new_n1047), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(new_n1062), .A3(new_n1054), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1058), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(G8), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1059), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1011), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(G2078), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n990), .A2(new_n993), .A3(new_n985), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1070), .A2(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n992), .B1(new_n1009), .B2(new_n488), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n961), .B1(new_n1076), .B2(new_n954), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1010), .A2(KEYINPUT109), .ZN(new_n1078));
  INV_X1    g653(.A(G2078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1049), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1071), .ZN(new_n1081));
  AOI21_X1  g656(.A(G301), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1021), .A2(new_n1026), .A3(new_n1069), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1065), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT63), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1012), .A2(new_n999), .A3(G286), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1063), .A2(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1058), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1046), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT113), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n1093), .B(new_n1046), .C1(new_n1089), .C2(new_n1058), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1088), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1085), .B1(new_n1096), .B2(new_n1087), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1027), .B(new_n675), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1031), .B1(new_n1099), .B2(new_n1043), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1083), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1080), .A2(new_n1071), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1072), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1105), .B(G301), .C1(new_n1011), .C2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1077), .A2(new_n1078), .A3(new_n1049), .A4(new_n1072), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1109), .A2(new_n1105), .ZN(new_n1110));
  AOI21_X1  g685(.A(G301), .B1(new_n1110), .B2(new_n1081), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1103), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1105), .ZN(new_n1113));
  OAI21_X1  g688(.A(G171), .B1(new_n1104), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1075), .A2(new_n1081), .A3(G301), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(KEYINPUT124), .A3(KEYINPUT54), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1082), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(G301), .A3(new_n1081), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1117), .B(new_n1122), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1096), .A2(KEYINPUT123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1059), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT125), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1112), .A2(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1069), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1077), .A2(new_n1078), .A3(new_n1049), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT116), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1049), .A2(new_n955), .A3(new_n985), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1078), .A4(new_n1133), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT115), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n559), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT115), .B(KEYINPUT57), .C1(new_n550), .C2(new_n558), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT114), .B(G1956), .Z(new_n1145));
  NOR2_X1   g720(.A1(new_n1006), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1139), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT61), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1144), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT118), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G1348), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1073), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n985), .A2(new_n986), .A3(new_n727), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1155), .A2(new_n819), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n819), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT60), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n819), .A2(KEYINPUT60), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1155), .A2(new_n1160), .A3(new_n1156), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n534), .A2(KEYINPUT117), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1077), .A2(new_n1078), .A3(new_n970), .A4(new_n1049), .ZN(new_n1164));
  XOR2_X1   g739(.A(KEYINPUT58), .B(G1341), .Z(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1076), .B2(new_n961), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT59), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1162), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1148), .B1(new_n1151), .B2(new_n1150), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1139), .B2(new_n1147), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT118), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1173), .B(new_n1174), .C1(new_n1151), .C2(new_n1150), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1153), .A2(new_n1169), .A3(new_n1172), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1148), .B1(new_n1152), .B2(new_n1158), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1102), .B1(new_n1132), .B2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G290), .B(new_n977), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n963), .B1(new_n974), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n983), .B1(new_n1182), .B2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g760(.A(G319), .ZN(new_n1187));
  NOR2_X1   g761(.A1(G227), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n670), .A2(new_n636), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1189), .B1(new_n871), .B2(new_n874), .ZN(new_n1190));
  OAI211_X1 g764(.A(new_n1190), .B(new_n940), .C1(new_n942), .C2(new_n948), .ZN(G225));
  INV_X1    g765(.A(G225), .ZN(G308));
endmodule


