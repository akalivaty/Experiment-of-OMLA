//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT0), .A3(G128), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n200), .A2(new_n202), .A3(new_n206), .A4(new_n203), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n205), .A2(KEYINPUT67), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT67), .B1(new_n205), .B2(new_n207), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n197), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n214), .A2(new_n215), .B1(KEYINPUT2), .B2(G113), .ZN(new_n216));
  INV_X1    g030(.A(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G116), .ZN(new_n218));
  INV_X1    g032(.A(G116), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G119), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT66), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n216), .B2(new_n222), .ZN(new_n224));
  INV_X1    g038(.A(new_n216), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT66), .A3(new_n221), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n195), .A2(new_n228), .A3(G128), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT64), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n230), .B1(new_n235), .B2(new_n188), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n229), .B1(new_n236), .B2(new_n195), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n199), .A2(G137), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n201), .A2(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n207), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT68), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n207), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n237), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n210), .A2(new_n227), .A3(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n210), .A2(KEYINPUT30), .A3(new_n245), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n216), .A2(new_n222), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n223), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n241), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n205), .A2(new_n207), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n237), .A2(new_n250), .B1(new_n197), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n249), .B1(new_n252), .B2(KEYINPUT30), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n246), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G237), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT27), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n197), .A2(new_n251), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n189), .A2(G146), .ZN(new_n265));
  OAI21_X1  g079(.A(G128), .B1(new_n228), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n188), .A2(new_n190), .A3(G128), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n266), .A2(new_n191), .B1(new_n228), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n268), .B2(new_n241), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n249), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n246), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n260), .B(KEYINPUT69), .Z(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n210), .A2(new_n245), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n249), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n210), .A2(KEYINPUT71), .A3(new_n245), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT28), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n262), .B(new_n263), .C1(new_n276), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n194), .A2(new_n196), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n251), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n205), .A2(KEYINPUT67), .A3(new_n207), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n237), .A2(new_n242), .A3(new_n244), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT72), .B(new_n249), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n246), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT72), .B1(new_n277), .B2(new_n249), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT28), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n227), .A3(new_n280), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n292), .A2(KEYINPUT29), .A3(new_n296), .A4(new_n260), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n282), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G472), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n274), .ZN(new_n302));
  INV_X1    g116(.A(new_n275), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n246), .B(new_n260), .C1(new_n247), .C2(new_n253), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT30), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n269), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n308), .B(new_n249), .C1(new_n277), .C2(new_n307), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n309), .A2(KEYINPUT31), .A3(new_n246), .A4(new_n260), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n302), .A2(new_n303), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G472), .A2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n301), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n313), .A2(new_n301), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n311), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n310), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n272), .B1(new_n246), .B2(new_n270), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n303), .B1(new_n281), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n300), .A2(new_n314), .A3(new_n318), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(G234), .B2(new_n298), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n217), .B2(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n217), .A2(G128), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n230), .A2(KEYINPUT23), .A3(G119), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G110), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n230), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT24), .B(G110), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT74), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n334), .A2(new_n341), .A3(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n344), .A2(KEYINPUT16), .A3(G140), .ZN(new_n345));
  XNOR2_X1  g159(.A(G125), .B(G140), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(KEYINPUT16), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G146), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n187), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n347), .B(G146), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n332), .A2(new_n333), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n336), .A2(new_n337), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G137), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n256), .A2(G221), .A3(G234), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n358), .B(new_n359), .Z(new_n360));
  NAND3_X1  g174(.A1(new_n352), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n360), .ZN(new_n362));
  INV_X1    g176(.A(new_n357), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n350), .B1(new_n340), .B2(new_n342), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n365), .A3(new_n298), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n361), .A2(new_n365), .A3(KEYINPUT25), .A4(new_n298), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n327), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n361), .A2(new_n365), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n326), .A2(G902), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n324), .A2(KEYINPUT75), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT75), .B1(new_n324), .B2(new_n374), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G221), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT9), .B(G234), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n380), .B2(new_n298), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT76), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(new_n298), .ZN(new_n384));
  XNOR2_X1  g198(.A(G110), .B(G140), .ZN(new_n385));
  INV_X1    g199(.A(G227), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G953), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n385), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(new_n389), .B2(G107), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT77), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G104), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT77), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n392), .A3(G104), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n397), .A2(new_n392), .A3(KEYINPUT78), .A4(G104), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n392), .A2(G104), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(G101), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n197), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n395), .A2(new_n391), .B1(new_n400), .B2(new_n401), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n403), .A2(G101), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(G101), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n404), .A2(new_n393), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n410), .A2(new_n411), .B1(G101), .B2(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n195), .A2(new_n228), .A3(G128), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT79), .B1(new_n265), .B2(new_n231), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n188), .A2(new_n419), .A3(KEYINPUT1), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(G128), .A3(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n421), .A2(new_n191), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n416), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n409), .A2(new_n414), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n208), .A2(new_n209), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n396), .A2(new_n402), .A3(new_n411), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n415), .A2(G101), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n427), .A2(KEYINPUT81), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT81), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT10), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n268), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT82), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n428), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n427), .A2(KEYINPUT81), .A3(new_n428), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n437), .A2(KEYINPUT82), .A3(new_n438), .A4(new_n433), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n425), .B(new_n426), .C1(new_n434), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n268), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n423), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n251), .A2(KEYINPUT12), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n426), .B1(new_n423), .B2(new_n442), .ZN(new_n445));
  OAI22_X1  g259(.A1(new_n443), .A2(new_n444), .B1(new_n445), .B2(KEYINPUT12), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n417), .B1(new_n191), .B2(new_n421), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n424), .B1(new_n435), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G101), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n410), .B2(new_n404), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n449), .B1(new_n453), .B2(new_n408), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n437), .A2(new_n438), .A3(new_n433), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n457), .B2(new_n439), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n388), .B1(new_n458), .B2(new_n426), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n425), .B1(new_n434), .B2(new_n440), .ZN(new_n460));
  INV_X1    g274(.A(new_n426), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n388), .A2(new_n447), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n384), .B1(new_n463), .B2(G469), .ZN(new_n464));
  INV_X1    g278(.A(new_n388), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n462), .B2(new_n441), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n441), .A2(new_n465), .A3(new_n446), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n383), .B(new_n298), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n382), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G214), .B1(G237), .B2(G902), .ZN(new_n470));
  OAI21_X1  g284(.A(G210), .B1(G237), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n249), .A2(new_n407), .A3(new_n414), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n474));
  OAI21_X1  g288(.A(G113), .B1(new_n474), .B2(new_n218), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n222), .A2(new_n474), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n476), .A2(new_n477), .B1(new_n216), .B2(new_n222), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n437), .A2(new_n478), .A3(new_n438), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G122), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(KEYINPUT6), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n472), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT84), .B(new_n484), .C1(new_n473), .C2(new_n479), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT6), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n481), .B1(new_n473), .B2(new_n479), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n483), .A2(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n283), .A2(G125), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n344), .B(new_n229), .C1(new_n236), .C2(new_n195), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n256), .A2(G224), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT85), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n484), .B1(new_n473), .B2(new_n479), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n472), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n499));
  INV_X1    g313(.A(new_n495), .ZN(new_n500));
  INV_X1    g314(.A(new_n488), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n486), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT7), .B1(new_n256), .B2(G224), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n490), .B2(new_n491), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n481), .B(KEYINPUT8), .Z(new_n509));
  AND3_X1   g323(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT5), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n225), .A2(new_n221), .B1(new_n475), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n416), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n478), .A2(new_n435), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n507), .B1(new_n493), .B2(new_n494), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n298), .B1(new_n505), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT86), .B(new_n298), .C1(new_n505), .C2(new_n516), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n471), .B1(new_n504), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n471), .ZN(new_n524));
  AOI211_X1 g338(.A(new_n524), .B(new_n521), .C1(new_n496), .C2(new_n503), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n469), .B(new_n470), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n347), .B(new_n187), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n255), .A2(new_n256), .A3(G214), .ZN(new_n528));
  NOR2_X1   g342(.A1(KEYINPUT87), .A2(G143), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(KEYINPUT87), .A2(G143), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n528), .B1(new_n531), .B2(new_n529), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n206), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n530), .A2(new_n532), .A3(new_n206), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n530), .A2(new_n532), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT17), .A3(G131), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(KEYINPUT89), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n533), .B2(KEYINPUT17), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n527), .B(new_n537), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n533), .A2(KEYINPUT18), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n346), .B(new_n187), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT18), .A2(G131), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n530), .A2(new_n532), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(G104), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT90), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n543), .A2(KEYINPUT90), .A3(new_n554), .A4(new_n551), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n298), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G475), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT20), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n534), .A2(new_n536), .ZN(new_n561));
  INV_X1    g375(.A(new_n346), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT19), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n562), .A2(KEYINPUT88), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT88), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT19), .B1(new_n346), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n187), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n561), .A2(new_n348), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n554), .B1(new_n545), .B2(new_n549), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n554), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n552), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(G475), .A2(G902), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n560), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n554), .B1(new_n543), .B2(new_n551), .ZN(new_n575));
  INV_X1    g389(.A(new_n573), .ZN(new_n576));
  NOR4_X1   g390(.A1(new_n575), .A2(new_n570), .A3(KEYINPUT20), .A4(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n559), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G122), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G116), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n580), .B(KEYINPUT14), .Z(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(KEYINPUT91), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G122), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n219), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G107), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n580), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n582), .A2(new_n584), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n392), .B(new_n587), .C1(new_n588), .C2(new_n219), .ZN(new_n589));
  XNOR2_X1  g403(.A(G128), .B(G143), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n199), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n586), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G107), .B1(new_n585), .B2(new_n580), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT13), .B1(new_n230), .B2(G143), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n199), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(new_n590), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n594), .A2(new_n597), .A3(KEYINPUT92), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT92), .B1(new_n594), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n592), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n379), .A2(new_n325), .A3(G953), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n592), .B(new_n601), .C1(new_n598), .C2(new_n599), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(KEYINPUT93), .A3(new_n298), .ZN(new_n606));
  INV_X1    g420(.A(G478), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(KEYINPUT15), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n603), .B2(new_n604), .ZN(new_n610));
  INV_X1    g424(.A(new_n608), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(KEYINPUT93), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G952), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(G953), .ZN(new_n615));
  NAND2_X1  g429(.A1(G234), .A2(G237), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(G902), .A3(G953), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT21), .B(G898), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n578), .A2(new_n613), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n526), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n377), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  NAND2_X1  g441(.A1(new_n464), .A2(new_n468), .ZN(new_n628));
  INV_X1    g442(.A(new_n382), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n322), .A2(new_n298), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G472), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n632), .B(new_n374), .C1(new_n311), .C2(new_n313), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n470), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n504), .A2(new_n522), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n524), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n504), .A2(new_n471), .A3(new_n522), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n622), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n607), .A2(G902), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n603), .A2(new_n643), .A3(new_n604), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n603), .B2(new_n604), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n641), .B(new_n642), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n642), .ZN(new_n648));
  INV_X1    g462(.A(new_n646), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n644), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT94), .B1(new_n610), .B2(G478), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n568), .A2(new_n569), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n540), .A2(new_n542), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n537), .A2(new_n527), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n550), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n653), .B(new_n573), .C1(new_n656), .C2(new_n554), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT20), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n572), .A2(new_n560), .A3(new_n573), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n658), .A2(new_n659), .B1(G475), .B2(new_n558), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n634), .A2(new_n639), .A3(new_n640), .A4(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT95), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n660), .A2(new_n613), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n634), .A2(new_n639), .A3(new_n640), .A4(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  INV_X1    g484(.A(KEYINPUT97), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n368), .A2(new_n369), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n326), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT96), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n352), .B2(new_n357), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n362), .A2(KEYINPUT36), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n352), .A2(new_n674), .A3(new_n357), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT96), .ZN(new_n680));
  OAI22_X1  g494(.A1(new_n680), .A2(new_n675), .B1(KEYINPUT36), .B2(new_n362), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n373), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n671), .B1(new_n673), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n373), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n679), .B2(new_n681), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n370), .A2(new_n686), .A3(KEYINPUT97), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n311), .A2(new_n313), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(G472), .B2(new_n631), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n639), .A2(new_n691), .A3(new_n469), .A4(new_n623), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT98), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n692), .B(new_n694), .ZN(G12));
  NAND2_X1  g509(.A1(new_n324), .A2(new_n688), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n620), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n617), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n660), .A2(new_n613), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n639), .A3(new_n469), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT99), .B(G128), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G30));
  NOR2_X1   g518(.A1(new_n370), .A2(new_n686), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n470), .A3(new_n578), .A4(new_n613), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n318), .A2(new_n323), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n303), .B1(new_n290), .B2(new_n291), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n304), .B1(new_n708), .B2(KEYINPUT100), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n298), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G472), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n314), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n699), .B(KEYINPUT39), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n469), .A2(new_n715), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n706), .B(new_n714), .C1(KEYINPUT40), .C2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n525), .A2(new_n523), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT38), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n717), .B(new_n720), .C1(KEYINPUT40), .C2(new_n716), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT101), .B(G143), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G45));
  INV_X1    g537(.A(new_n699), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n652), .A2(new_n660), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n324), .A2(new_n688), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n639), .A3(new_n727), .A4(new_n469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n324), .A2(new_n688), .A3(new_n725), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT102), .B1(new_n526), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  NAND3_X1  g546(.A1(new_n639), .A2(new_n640), .A3(new_n661), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n324), .A2(new_n374), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n298), .B1(new_n466), .B2(new_n467), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n737));
  INV_X1    g551(.A(new_n381), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n468), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n738), .A3(new_n468), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n734), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n733), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT41), .B(G113), .Z(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G15));
  NAND3_X1  g559(.A1(new_n639), .A2(new_n640), .A3(new_n667), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n742), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n219), .ZN(G18));
  NAND2_X1  g562(.A1(new_n741), .A2(new_n739), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n470), .B1(new_n525), .B2(new_n523), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n624), .A4(new_n696), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n217), .ZN(G21));
  INV_X1    g566(.A(new_n749), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n609), .A2(new_n612), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(new_n660), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n578), .A2(new_n613), .A3(KEYINPUT105), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n640), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT104), .B(G472), .Z(new_n760));
  NAND2_X1  g574(.A1(new_n631), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n319), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n275), .B1(new_n292), .B2(new_n296), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n312), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n374), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n753), .A2(new_n754), .A3(new_n639), .A4(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n639), .A2(new_n766), .A3(new_n739), .A4(new_n741), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT106), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT107), .B(G122), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G24));
  INV_X1    g586(.A(new_n725), .ZN(new_n773));
  INV_X1    g587(.A(new_n705), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n761), .A2(new_n774), .A3(new_n764), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(new_n639), .A3(new_n739), .A4(new_n741), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  NOR3_X1   g592(.A1(new_n525), .A2(new_n523), .A3(new_n635), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n773), .A2(KEYINPUT42), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n381), .B1(new_n464), .B2(new_n468), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n734), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n637), .A2(new_n781), .A3(new_n470), .A4(new_n638), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n300), .A2(new_n314), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n311), .A2(new_n317), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n725), .B(new_n374), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT42), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  XNOR2_X1  g603(.A(new_n700), .B(KEYINPUT108), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n779), .A2(new_n734), .A3(new_n781), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  OR2_X1    g606(.A1(new_n652), .A2(new_n578), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT43), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n690), .A2(new_n705), .ZN(new_n796));
  OR3_X1    g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n779), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n468), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n463), .A2(KEYINPUT45), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n383), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n463), .A2(KEYINPUT45), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n384), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n802), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(KEYINPUT46), .A3(new_n807), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n381), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(new_n715), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n797), .A2(KEYINPUT109), .A3(new_n779), .A4(new_n798), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n801), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  OR2_X1    g630(.A1(new_n812), .A2(KEYINPUT47), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n812), .A2(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n773), .A2(new_n324), .A3(new_n374), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n637), .A2(new_n470), .A3(new_n638), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n819), .A2(KEYINPUT110), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT110), .B1(new_n819), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(G140), .Z(G42));
  NAND2_X1  g640(.A1(new_n736), .A2(new_n468), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n374), .A2(new_n470), .A3(new_n629), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n793), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n714), .A2(new_n828), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n720), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n817), .B(new_n818), .C1(new_n629), .C2(new_n827), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n794), .A2(new_n617), .A3(new_n765), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n836), .A2(new_n779), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n749), .A2(new_n821), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(new_n618), .A3(new_n374), .A4(new_n714), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n660), .A3(new_n652), .A4(new_n843), .ZN(new_n844));
  OR2_X1    g658(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n837), .A2(new_n635), .A3(new_n719), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n846), .A2(new_n749), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n846), .B2(new_n749), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n794), .A2(new_n617), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n839), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n851), .A2(new_n775), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n844), .A2(new_n848), .A3(new_n849), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n835), .B1(new_n838), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n848), .A2(new_n849), .A3(new_n852), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n836), .A2(new_n779), .A3(new_n837), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT51), .A4(new_n844), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n374), .B1(new_n784), .B2(new_n785), .ZN(new_n859));
  OR3_X1    g673(.A1(new_n851), .A2(KEYINPUT48), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT48), .B1(new_n851), .B2(new_n859), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n842), .A2(new_n661), .A3(new_n843), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n837), .A2(new_n639), .A3(new_n753), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n615), .A4(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT116), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  INV_X1    g682(.A(new_n751), .ZN(new_n869));
  INV_X1    g683(.A(new_n661), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n750), .A2(new_n622), .A3(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n750), .A2(new_n622), .A3(new_n666), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n734), .B(new_n753), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n770), .A2(new_n869), .A3(new_n873), .A4(new_n788), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n781), .A2(new_n705), .A3(new_n699), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n757), .A2(new_n758), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n639), .A3(new_n713), .A4(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n731), .A2(new_n702), .A3(new_n777), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT52), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n702), .A2(new_n777), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n731), .A4(new_n878), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n626), .A2(new_n662), .A3(new_n668), .A4(new_n692), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n779), .A2(new_n776), .A3(new_n781), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n791), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n756), .A2(new_n660), .A3(new_n887), .A4(new_n699), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n609), .A2(new_n612), .A3(new_n699), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT111), .B1(new_n889), .B2(new_n578), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n469), .A2(new_n324), .A3(new_n891), .A4(new_n688), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n779), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n469), .A2(new_n891), .A3(new_n324), .A4(new_n688), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT112), .B1(new_n895), .B2(new_n821), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n884), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n875), .A2(new_n880), .A3(new_n883), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n884), .A2(new_n898), .A3(new_n901), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n875), .A3(new_n880), .A4(new_n883), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n868), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT113), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n791), .A2(new_n885), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n894), .B2(new_n896), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n375), .A2(new_n376), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n639), .A2(new_n469), .A3(new_n623), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n662), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n668), .A2(new_n692), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n909), .A2(new_n914), .A3(KEYINPUT53), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n874), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n880), .A2(new_n883), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT113), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n907), .A2(new_n918), .B1(new_n901), .B2(new_n900), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n905), .B1(new_n919), .B2(new_n868), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n867), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(G952), .A2(G953), .ZN(new_n922));
  OAI211_X1 g736(.A(KEYINPUT117), .B(new_n834), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n867), .B2(new_n920), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n833), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n926), .ZN(G75));
  XNOR2_X1  g741(.A(new_n489), .B(new_n500), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT55), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT113), .B1(new_n916), .B2(new_n917), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n880), .A2(new_n883), .ZN(new_n932));
  NOR4_X1   g746(.A1(new_n932), .A2(new_n915), .A3(new_n906), .A4(new_n874), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n902), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(G210), .A2(G902), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT118), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n907), .A2(new_n918), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n935), .B1(new_n940), .B2(new_n902), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT118), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n930), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n614), .A2(G953), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT119), .Z(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n929), .A2(KEYINPUT56), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT120), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT56), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n941), .B2(KEYINPUT118), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n937), .A2(new_n938), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n929), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT120), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n955), .A3(new_n948), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n950), .A2(new_n956), .ZN(G51));
  NAND2_X1  g771(.A1(new_n919), .A2(new_n868), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n934), .A2(KEYINPUT54), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT121), .ZN(new_n960));
  OR3_X1    g774(.A1(new_n919), .A2(KEYINPUT121), .A3(new_n868), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n384), .B(KEYINPUT57), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n466), .A2(new_n467), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n919), .A2(new_n298), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(new_n805), .A3(new_n804), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n946), .B1(new_n965), .B2(new_n967), .ZN(G54));
  NAND3_X1  g782(.A1(new_n966), .A2(KEYINPUT58), .A3(G475), .ZN(new_n969));
  INV_X1    g783(.A(new_n572), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n972), .A3(new_n946), .ZN(G60));
  NOR2_X1   g787(.A1(new_n645), .A2(new_n646), .ZN(new_n974));
  NAND2_X1  g788(.A1(G478), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT59), .Z(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n920), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n945), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n960), .A2(new_n961), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n974), .A2(new_n976), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G63));
  XNOR2_X1  g795(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n325), .A2(new_n298), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n934), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n946), .B1(new_n985), .B2(new_n371), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n987));
  INV_X1    g801(.A(new_n984), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n919), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n987), .B1(new_n989), .B2(new_n682), .ZN(new_n990));
  INV_X1    g804(.A(new_n682), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n985), .A2(KEYINPUT123), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n986), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(KEYINPUT61), .B(new_n986), .C1(new_n990), .C2(new_n992), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(G66));
  INV_X1    g811(.A(G224), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n621), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n742), .B1(new_n733), .B2(new_n746), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(new_n751), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n914), .A2(new_n1001), .A3(new_n770), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n489), .B1(G898), .B2(new_n256), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G69));
  OAI21_X1  g820(.A(G953), .B1(new_n386), .B2(new_n697), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n308), .B1(new_n277), .B2(new_n307), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT124), .Z(new_n1009));
  NOR2_X1   g823(.A1(new_n564), .A2(new_n566), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1009), .B(new_n1010), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n881), .A2(new_n731), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n639), .A2(new_n877), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1014), .A2(new_n859), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n813), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n788), .A2(new_n791), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n815), .A2(new_n1013), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n256), .B1(new_n825), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n256), .A2(G900), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(KEYINPUT126), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1019), .A2(KEYINPUT126), .A3(new_n1021), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1012), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1013), .A2(new_n721), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n716), .B1(new_n870), .B2(new_n666), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n377), .A2(new_n779), .A3(new_n1028), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n1027), .A2(new_n815), .A3(new_n1029), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(KEYINPUT125), .B1(new_n1032), .B2(new_n825), .ZN(new_n1033));
  INV_X1    g847(.A(new_n825), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT125), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1034), .A2(new_n1035), .A3(new_n1031), .A4(new_n1030), .ZN(new_n1036));
  AOI211_X1 g850(.A(G953), .B(new_n1011), .C1(new_n1033), .C2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1007), .B1(new_n1025), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1024), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1011), .B1(new_n1039), .B2(new_n1022), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1041), .A2(new_n256), .A3(new_n1012), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1007), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1038), .A2(new_n1044), .ZN(G72));
  XNOR2_X1  g859(.A(new_n254), .B(KEYINPUT127), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n260), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1033), .A2(new_n1003), .A3(new_n1036), .ZN(new_n1048));
  NAND2_X1  g862(.A1(G472), .A2(G902), .ZN(new_n1049));
  XOR2_X1   g863(.A(new_n1049), .B(KEYINPUT63), .Z(new_n1050));
  AOI21_X1  g864(.A(new_n1047), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OR3_X1    g865(.A1(new_n825), .A2(new_n1002), .A3(new_n1018), .ZN(new_n1052));
  AOI211_X1 g866(.A(new_n260), .B(new_n1046), .C1(new_n1052), .C2(new_n1050), .ZN(new_n1053));
  AND2_X1   g867(.A1(new_n902), .A2(new_n904), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n262), .A2(new_n304), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1055), .A2(new_n1050), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n945), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g871(.A1(new_n1051), .A2(new_n1053), .A3(new_n1057), .ZN(G57));
endmodule


