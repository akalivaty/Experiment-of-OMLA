//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(KEYINPUT65), .B1(G567), .B2(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(G137), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G125), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(new_n482), .B1(G113), .B2(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(KEYINPUT67), .A3(G125), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n475), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(G160));
  XNOR2_X1  g062(.A(new_n469), .B(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n472), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  INV_X1    g066(.A(new_n475), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  NOR2_X1   g069(.A1(G100), .A2(G2105), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT71), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT72), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  XOR2_X1   g074(.A(new_n499), .B(KEYINPUT73), .Z(G162));
  NAND3_X1  g075(.A1(new_n470), .A2(G126), .A3(G2105), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n473), .A2(G138), .A3(new_n474), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n469), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n475), .A2(new_n507), .A3(G138), .A4(new_n480), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(G164));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  INV_X1    g088(.A(G75), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT75), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR3_X1    g091(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT75), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT74), .B1(new_n519), .B2(G651), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT6), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(new_n523), .B1(new_n519), .B2(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(G50), .A2(G543), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n518), .A2(G651), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n512), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n528), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n534), .A2(new_n535), .B1(new_n512), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n519), .A2(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n521), .B1(KEYINPUT6), .B2(new_n522), .ZN(new_n540));
  NOR3_X1   g115(.A1(new_n519), .A2(KEYINPUT74), .A3(G651), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n524), .A2(KEYINPUT76), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n544), .A2(G543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G51), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n538), .A2(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  AOI22_X1  g124(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n522), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT77), .Z(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n527), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n546), .A2(G52), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n512), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n528), .A2(G81), .B1(new_n560), .B2(G651), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n544), .A2(new_n545), .A3(G43), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT78), .ZN(G188));
  NAND4_X1  g145(.A1(new_n544), .A2(new_n545), .A3(G53), .A4(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n558), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n528), .A2(G91), .B1(new_n575), .B2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  OAI21_X1  g153(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n527), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n546), .B2(G49), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n524), .A2(G48), .A3(G543), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n585), .B2(new_n522), .C1(new_n527), .C2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n546), .A2(G47), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n558), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n528), .A2(G85), .B1(new_n591), .B2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G290));
  XOR2_X1   g168(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT80), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n524), .A2(G92), .A3(new_n512), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND4_X1  g172(.A1(new_n544), .A2(new_n545), .A3(G54), .A4(G543), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n522), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(KEYINPUT81), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT81), .B1(new_n598), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G321));
  XNOR2_X1  g182(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(new_n576), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n609), .B1(new_n613), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n609), .B1(new_n613), .B2(G868), .ZN(G280));
  XNOR2_X1  g190(.A(new_n595), .B(new_n596), .ZN(new_n616));
  INV_X1    g191(.A(new_n603), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n601), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  NOR2_X1   g195(.A1(new_n564), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n618), .A2(new_n619), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI221_X1 g200(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n475), .C2(G111), .ZN(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  INV_X1    g202(.A(G123), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n488), .A2(new_n492), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n626), .B1(new_n489), .B2(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(G2096), .ZN(new_n632));
  INV_X1    g207(.A(new_n478), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n480), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n631), .A2(new_n632), .A3(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT84), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n645), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(G14), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT85), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  AOI211_X1 g252(.A(new_n674), .B(new_n677), .C1(new_n669), .C2(new_n673), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1981), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT87), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n680), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G25), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT88), .ZN(new_n689));
  OAI21_X1  g264(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n690));
  INV_X1    g265(.A(G107), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n492), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n490), .B2(G131), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n493), .B2(G119), .ZN(new_n695));
  INV_X1    g270(.A(G119), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n629), .A2(KEYINPUT89), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n693), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n689), .B1(new_n698), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT35), .B(G1991), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G6), .B(G305), .S(G16), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n703), .A2(G23), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n582), .B2(new_n703), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT33), .B(G1976), .Z(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n707), .A2(new_n710), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT34), .Z(new_n717));
  NOR2_X1   g292(.A1(G16), .A2(G24), .ZN(new_n718));
  XNOR2_X1  g293(.A(G290), .B(KEYINPUT91), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G1986), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n702), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT36), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n687), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  OAI221_X1 g301(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n475), .C2(G116), .ZN(new_n727));
  INV_X1    g302(.A(G140), .ZN(new_n728));
  INV_X1    g303(.A(G128), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n727), .B1(new_n489), .B2(new_n728), .C1(new_n729), .C2(new_n629), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n726), .B1(new_n731), .B2(new_n687), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT93), .B(G2067), .Z(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(G160), .A2(G29), .ZN(new_n735));
  INV_X1    g310(.A(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n736), .B2(KEYINPUT24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(KEYINPUT24), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n490), .A2(G141), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n493), .A2(G129), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT26), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n746), .A2(new_n747), .B1(G105), .B2(new_n633), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n742), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n687), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n687), .B2(G32), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n734), .B(new_n741), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n703), .A2(G19), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n564), .B2(new_n703), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NOR2_X1   g332(.A1(G171), .A2(new_n703), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G5), .B2(new_n703), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(new_n760), .B2(G1961), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n703), .A2(G20), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n613), .B2(new_n703), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G164), .A2(new_n687), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G27), .B2(new_n687), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G28), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT30), .ZN(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n772), .B2(KEYINPUT30), .ZN(new_n774));
  OR2_X1    g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n769), .A2(new_n770), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n630), .A2(new_n687), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n771), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n733), .B2(new_n732), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n754), .A2(new_n761), .A3(new_n767), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n703), .A2(G4), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n618), .B2(new_n703), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT92), .B(G1348), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n784), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(G168), .A2(G16), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G21), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(KEYINPUT95), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(KEYINPUT95), .B2(new_n788), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n687), .A2(G33), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT25), .Z(new_n796));
  AOI22_X1  g371(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n797));
  INV_X1    g372(.A(G139), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n796), .B1(new_n475), .B2(new_n797), .C1(new_n798), .C2(new_n489), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT94), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n794), .B1(new_n800), .B2(new_n687), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2072), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n782), .A2(new_n787), .A3(new_n793), .A4(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n759), .A2(new_n804), .B1(new_n740), .B2(new_n739), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n752), .B2(new_n753), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT96), .ZN(new_n807));
  NOR2_X1   g382(.A1(G29), .A2(G35), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G162), .B2(G29), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G2090), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n724), .A2(new_n803), .A3(new_n807), .A4(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NOR2_X1   g390(.A1(new_n604), .A2(new_n619), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(G80), .A2(G543), .ZN(new_n819));
  INV_X1    g394(.A(G67), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n558), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n528), .A2(G93), .B1(new_n821), .B2(G651), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT100), .B(G55), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n544), .A2(new_n545), .A3(G543), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n563), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n563), .A2(new_n825), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n818), .B(new_n828), .Z(new_n829));
  AND2_X1   g404(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n830), .A2(new_n831), .A3(G860), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n825), .A2(G860), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n832), .A2(new_n834), .ZN(G145));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n698), .B(KEYINPUT103), .ZN(new_n837));
  OAI221_X1 g412(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n475), .C2(G118), .ZN(new_n838));
  INV_X1    g413(.A(G130), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n629), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G142), .B2(new_n490), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n837), .B(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n635), .B(KEYINPUT102), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n501), .A2(new_n503), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT101), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT101), .B1(new_n506), .B2(new_n508), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n730), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n749), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n799), .ZN(new_n851));
  INV_X1    g426(.A(new_n800), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n844), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(G160), .B(new_n630), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G162), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n851), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n842), .A2(new_n843), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n842), .A2(new_n843), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n856), .B1(new_n854), .B2(new_n860), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n836), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n866), .A2(KEYINPUT40), .A3(new_n862), .A4(new_n861), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(G395));
  NAND2_X1  g443(.A1(new_n825), .A2(new_n605), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT104), .B1(new_n618), .B2(G299), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n604), .A2(new_n613), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n604), .A2(new_n613), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n622), .B(new_n828), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n874), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n870), .A2(new_n872), .A3(KEYINPUT41), .A4(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n870), .A2(KEYINPUT105), .A3(new_n872), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n874), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n879), .B1(new_n883), .B2(KEYINPUT41), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n877), .B1(new_n884), .B2(new_n876), .ZN(new_n885));
  XNOR2_X1  g460(.A(G288), .B(G290), .ZN(new_n886));
  XOR2_X1   g461(.A(G303), .B(G305), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT42), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n885), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n869), .B1(new_n890), .B2(new_n605), .ZN(G295));
  OAI21_X1  g466(.A(new_n869), .B1(new_n890), .B2(new_n605), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n893));
  NOR3_X1   g468(.A1(G168), .A2(new_n826), .A3(new_n827), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n563), .A2(new_n825), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n563), .A2(new_n825), .ZN(new_n896));
  AOI21_X1  g471(.A(G286), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(G301), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n828), .A2(G286), .ZN(new_n899));
  OAI21_X1  g474(.A(G168), .B1(new_n826), .B2(new_n827), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(G171), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n879), .B(new_n902), .C1(new_n883), .C2(KEYINPUT41), .ZN(new_n903));
  INV_X1    g478(.A(new_n875), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n888), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n862), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n888), .B1(new_n903), .B2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n905), .ZN(new_n912));
  INV_X1    g487(.A(new_n888), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n862), .A3(new_n906), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n898), .A2(new_n901), .A3(KEYINPUT41), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n875), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n888), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n883), .A2(new_n918), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n862), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n908), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT107), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n926));
  NOR4_X1   g501(.A1(new_n908), .A2(new_n922), .A3(new_n926), .A4(KEYINPUT43), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n893), .B1(new_n917), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n908), .B2(new_n922), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n930), .A2(KEYINPUT109), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n893), .B1(new_n930), .B2(KEYINPUT109), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n907), .A2(new_n908), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n924), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n915), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n931), .B(new_n932), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n929), .A2(new_n937), .ZN(G397));
  XNOR2_X1  g513(.A(KEYINPUT110), .B(G1384), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT45), .B1(new_n848), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n486), .A2(G40), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1996), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n749), .B(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G2067), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n730), .B(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n698), .A2(new_n701), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n698), .A2(new_n701), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(G290), .A2(G1986), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n588), .A2(new_n721), .A3(new_n592), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n943), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n486), .A2(G40), .ZN(new_n956));
  NOR2_X1   g531(.A1(G164), .A2(G1384), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n506), .A2(new_n508), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT101), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n504), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n960), .B1(new_n965), .B2(G1384), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n848), .A2(KEYINPUT112), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n959), .B1(new_n969), .B2(new_n958), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n766), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n848), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT111), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n848), .A2(new_n974), .A3(KEYINPUT45), .A4(new_n939), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n956), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n845), .A2(new_n961), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT45), .B1(new_n977), .B2(new_n967), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT56), .B(G2072), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n613), .B(KEYINPUT57), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n971), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n956), .B1(new_n966), .B2(new_n968), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n946), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n965), .A2(new_n960), .A3(G1384), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT112), .B1(new_n848), .B2(new_n967), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n958), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n977), .A2(new_n967), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n956), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n786), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n618), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT119), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT120), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n956), .B(new_n978), .C1(new_n973), .C2(new_n975), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n996), .A2(new_n980), .B1(new_n970), .B2(new_n766), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n997), .B2(new_n982), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n982), .B1(new_n971), .B2(new_n981), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT120), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n983), .B1(new_n994), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n971), .A2(new_n981), .ZN(new_n1004));
  INV_X1    g579(.A(new_n982), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n983), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT61), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n971), .A2(new_n981), .A3(new_n982), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1003), .B(new_n1008), .C1(new_n1010), .C2(new_n999), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n986), .A2(new_n992), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT50), .B1(new_n966), .B2(new_n968), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n941), .B1(new_n957), .B2(new_n958), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n604), .B(new_n985), .C1(new_n1018), .C2(new_n786), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n993), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1020), .B2(KEYINPUT60), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n969), .A2(new_n941), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT58), .B(G1341), .Z(new_n1023));
  AOI22_X1  g598(.A1(new_n996), .A2(new_n944), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT59), .B1(new_n1024), .B2(new_n563), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n976), .A2(new_n979), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1027), .B2(G1996), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n564), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT122), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n983), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n971), .A2(new_n981), .A3(KEYINPUT122), .A4(new_n982), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(KEYINPUT61), .A3(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1021), .B(new_n1031), .C1(new_n1001), .C2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1002), .B1(new_n1013), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1038), .B(new_n1039), .Z(new_n1040));
  AOI21_X1  g615(.A(G1971), .B1(new_n976), .B2(new_n979), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1016), .A2(new_n1017), .A3(G2090), .ZN(new_n1042));
  OAI211_X1 g617(.A(G8), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n984), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n582), .B2(G1976), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1045), .B(new_n1048), .C1(new_n1049), .C2(G288), .ZN(new_n1050));
  AND2_X1   g625(.A1(G305), .A2(G1981), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G305), .A2(G1981), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT116), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT115), .B1(new_n1056), .B2(KEYINPUT49), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1055), .A2(KEYINPUT49), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1045), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1022), .B(G8), .C1(new_n1049), .C2(G288), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1043), .A2(new_n1050), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1027), .A2(new_n706), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n812), .B(new_n959), .C1(new_n969), .C2(new_n958), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1040), .B1(new_n1065), .B2(G8), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n989), .A2(new_n991), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n940), .A2(new_n1069), .A3(G2078), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1068), .A2(new_n804), .B1(new_n976), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n973), .A2(new_n975), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1072), .A2(new_n770), .A3(new_n941), .A4(new_n979), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1069), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1071), .A2(new_n1074), .A3(G301), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n804), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n966), .A2(new_n1077), .A3(new_n968), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n956), .B1(new_n957), .B2(KEYINPUT45), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(KEYINPUT53), .A3(new_n770), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1076), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1074), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1075), .B1(new_n1084), .B2(G171), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1067), .B1(new_n1085), .B2(KEYINPUT54), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n792), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1018), .A2(new_n740), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(KEYINPUT117), .A3(new_n792), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1090), .A2(G168), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1093), .A2(new_n1094), .A3(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n1087), .B2(new_n792), .ZN(new_n1097));
  OAI21_X1  g672(.A(G286), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(G8), .A3(new_n1093), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(KEYINPUT51), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1086), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(G171), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT53), .B1(new_n996), .B2(new_n770), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT123), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1076), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1105), .B1(new_n1110), .B2(G301), .ZN(new_n1111));
  OAI211_X1 g686(.A(G301), .B(new_n1074), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(KEYINPUT124), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT125), .B(new_n1104), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1104), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AND4_X1   g692(.A1(new_n1037), .A2(new_n1101), .A3(new_n1114), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1100), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1093), .A2(G8), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1094), .B1(new_n1121), .B2(new_n1098), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT62), .B1(new_n1122), .B2(new_n1095), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1061), .A2(new_n1050), .A3(new_n1059), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1044), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1124), .B(new_n1043), .C1(new_n1125), .C2(new_n1040), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1126), .A2(G301), .A3(new_n1110), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1120), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1058), .A2(G1976), .A3(G288), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1045), .B1(new_n1129), .B2(new_n1052), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1124), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n1043), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G286), .A2(new_n1044), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1135), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1133), .B1(new_n1139), .B2(new_n1126), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1062), .ZN(new_n1141));
  OAI21_X1  g716(.A(G8), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1040), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1133), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1141), .B(new_n1144), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1132), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1128), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n955), .B1(new_n1118), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n943), .A2(new_n944), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT46), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n947), .A2(new_n750), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n942), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT126), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1153), .A2(KEYINPUT47), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(KEYINPUT47), .ZN(new_n1155));
  INV_X1    g730(.A(new_n949), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n948), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n731), .A2(new_n946), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n942), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n942), .A2(new_n953), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n951), .A2(new_n943), .B1(KEYINPUT48), .B2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1160), .A2(KEYINPUT48), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1154), .A2(new_n1155), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1148), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g740(.A1(new_n917), .A2(new_n928), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n461), .A2(G227), .ZN(new_n1168));
  NOR2_X1   g742(.A1(new_n1168), .A2(KEYINPUT127), .ZN(new_n1169));
  AND2_X1   g743(.A1(new_n1168), .A2(KEYINPUT127), .ZN(new_n1170));
  NOR4_X1   g744(.A1(G229), .A2(G401), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g745(.A(new_n1171), .B1(new_n863), .B2(new_n864), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1167), .A2(new_n1172), .ZN(G308));
  OAI221_X1 g747(.A(new_n1171), .B1(new_n863), .B2(new_n864), .C1(new_n917), .C2(new_n928), .ZN(G225));
endmodule


