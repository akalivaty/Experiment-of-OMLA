//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067;
  INV_X1    g000(.A(KEYINPUT0), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n187), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT64), .B1(new_n190), .B2(G146), .ZN(new_n196));
  OAI211_X1 g010(.A(G128), .B(new_n189), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(new_n187), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT65), .A2(G131), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT65), .A2(G131), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n212), .A2(new_n204), .A3(new_n206), .A4(new_n207), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n209), .A2(new_n213), .A3(KEYINPUT70), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT70), .B1(new_n209), .B2(new_n213), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n201), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G116), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G119), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT69), .B(G116), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G119), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n218), .B1(new_n222), .B2(KEYINPUT68), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n219), .A2(KEYINPUT69), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G116), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n226), .A3(G119), .ZN(new_n227));
  INV_X1    g041(.A(new_n220), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n217), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n190), .A2(G146), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n188), .B2(G143), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(G128), .ZN(new_n240));
  OAI21_X1  g054(.A(G128), .B1(new_n234), .B2(new_n239), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n192), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n205), .A2(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n207), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G131), .ZN(new_n247));
  XNOR2_X1  g061(.A(G134), .B(G137), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT66), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n243), .A2(new_n213), .A3(new_n247), .A4(new_n250), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n216), .A2(new_n233), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n233), .B1(new_n216), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT28), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n216), .A2(new_n233), .A3(new_n251), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT73), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n259), .A3(new_n256), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n254), .A2(new_n258), .A3(new_n260), .A4(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(G902), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n213), .A2(new_n250), .A3(new_n247), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n213), .A2(new_n250), .A3(new_n247), .A4(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n243), .A3(new_n275), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n198), .A2(new_n200), .B1(new_n213), .B2(new_n209), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n256), .A2(new_n255), .B1(new_n279), .B2(new_n232), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n216), .A2(new_n233), .A3(new_n251), .A4(KEYINPUT28), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n265), .A4(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n216), .A2(KEYINPUT30), .A3(new_n251), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT71), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n216), .A2(new_n286), .A3(new_n251), .A4(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n233), .B1(new_n279), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n252), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n283), .B1(new_n291), .B2(new_n265), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n279), .A2(new_n232), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n257), .A2(new_n293), .A3(new_n265), .A4(new_n282), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n267), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n271), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G472), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT32), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n265), .B1(new_n280), .B2(new_n282), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n272), .A2(KEYINPUT67), .B1(new_n242), .B2(new_n240), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n277), .B1(new_n302), .B2(new_n275), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n232), .B1(new_n303), .B2(KEYINPUT30), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n287), .B2(new_n285), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n255), .A2(new_n265), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n288), .A2(new_n290), .ZN(new_n308));
  INV_X1    g122(.A(new_n306), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT31), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n300), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G472), .A2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n299), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n300), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT31), .B1(new_n308), .B2(new_n309), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n301), .B(new_n306), .C1(new_n288), .C2(new_n290), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT32), .A3(new_n312), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n298), .A2(new_n314), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G217), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n270), .B2(G234), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT25), .ZN(new_n324));
  INV_X1    g138(.A(G953), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(G221), .A3(G234), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT76), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT22), .B(G137), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G128), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(G128), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n331), .B(new_n332), .C1(new_n333), .C2(KEYINPUT23), .ZN(new_n334));
  XOR2_X1   g148(.A(KEYINPUT24), .B(G110), .Z(new_n335));
  XNOR2_X1  g149(.A(G119), .B(G128), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n334), .A2(G110), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G125), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G140), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT16), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n340), .A2(G140), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT16), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n345), .A3(G146), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(G146), .B1(new_n342), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n337), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XOR2_X1   g163(.A(KEYINPUT75), .B(G110), .Z(new_n350));
  OAI22_X1  g164(.A1(new_n334), .A2(new_n350), .B1(new_n335), .B2(new_n336), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n338), .A2(G125), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n188), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n346), .A3(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n329), .A2(new_n349), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n329), .B1(new_n349), .B2(new_n355), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n270), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n324), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT25), .B(new_n270), .C1(new_n356), .C2(new_n357), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n323), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n358), .A2(G902), .A3(new_n322), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT9), .B(G234), .ZN(new_n365));
  OAI21_X1  g179(.A(G221), .B1(new_n365), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n214), .A2(new_n215), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(G104), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(KEYINPUT78), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n377), .A3(G104), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G101), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n374), .B(new_n382), .C1(new_n378), .C2(new_n379), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n380), .A2(new_n385), .A3(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n201), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT78), .B(G107), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n373), .B1(new_n388), .B2(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G101), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n243), .A2(KEYINPUT10), .A3(new_n390), .A4(new_n383), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n394), .B(KEYINPUT1), .C1(new_n190), .C2(G146), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G128), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n393), .B1(new_n398), .B2(new_n238), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n189), .B1(new_n195), .B2(new_n196), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(KEYINPUT80), .C1(new_n397), .C2(new_n396), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n240), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n390), .A2(new_n383), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT10), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n369), .B1(new_n392), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT81), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(new_n369), .C1(new_n392), .C2(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G140), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n325), .A2(G227), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n400), .B1(new_n397), .B2(new_n396), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n393), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n403), .B1(new_n417), .B2(new_n401), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n387), .B(new_n391), .C1(new_n418), .C2(KEYINPUT10), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n414), .B1(new_n419), .B2(new_n369), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT12), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n209), .B2(new_n213), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n403), .A2(new_n242), .A3(new_n240), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n402), .A2(new_n404), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n368), .B1(new_n427), .B2(new_n424), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n428), .B2(KEYINPUT12), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n392), .A2(new_n405), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n368), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n410), .A2(new_n421), .B1(new_n432), .B2(new_n413), .ZN(new_n433));
  OAI21_X1  g247(.A(G469), .B1(new_n433), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(G469), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n414), .B1(new_n410), .B2(new_n431), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n369), .B1(new_n418), .B2(new_n425), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n427), .A2(new_n424), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n437), .A2(new_n422), .B1(new_n438), .B2(new_n423), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n420), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n435), .B(new_n270), .C1(new_n436), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n367), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n224), .A2(new_n226), .A3(G122), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT14), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n219), .A2(G122), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n221), .A2(KEYINPUT14), .A3(G122), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(G107), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT95), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n444), .A2(new_n446), .ZN(new_n451));
  XNOR2_X1  g265(.A(G128), .B(G143), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n452), .A2(new_n203), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n203), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n451), .A2(new_n388), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n447), .A2(new_n456), .A3(G107), .A4(new_n448), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n450), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n193), .A2(G143), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n203), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n452), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n451), .A2(new_n388), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n444), .A2(new_n388), .A3(new_n446), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n365), .A2(new_n321), .A3(G953), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n458), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n458), .B2(new_n465), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n443), .B(new_n270), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G478), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n270), .B1(new_n467), .B2(new_n468), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT96), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  INV_X1    g289(.A(new_n471), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G952), .ZN(new_n478));
  AOI211_X1 g292(.A(G953), .B(new_n478), .C1(G234), .C2(G237), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n325), .B(new_n270), .C1(G234), .C2(G237), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(G898), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G902), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n343), .B2(new_n352), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT89), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(G146), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n353), .B2(new_n188), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n486), .A2(new_n489), .A3(G146), .A4(new_n487), .ZN(new_n492));
  AND2_X1   g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n261), .A2(G214), .B1(new_n494), .B2(G143), .ZN(new_n495));
  INV_X1    g309(.A(G214), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n496), .A2(G237), .A3(G953), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(G143), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n190), .A2(KEYINPUT88), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n495), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n493), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n190), .A2(KEYINPUT88), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n494), .A2(G143), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n497), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G237), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n325), .A3(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n498), .ZN(new_n509));
  AND4_X1   g323(.A1(new_n502), .A2(new_n506), .A3(new_n493), .A4(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n491), .B(new_n492), .C1(new_n503), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n212), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n508), .B1(new_n498), .B2(new_n499), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n495), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n506), .A2(new_n212), .A3(new_n509), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n347), .A2(new_n348), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT17), .B(new_n512), .C1(new_n513), .C2(new_n495), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G113), .B(G122), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n521), .B(G104), .Z(new_n522));
  AND3_X1   g336(.A1(new_n511), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n511), .B2(new_n520), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n484), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G475), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n527));
  NOR2_X1   g341(.A1(G475), .A2(G902), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT93), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n347), .B1(new_n514), .B2(new_n516), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n486), .A2(KEYINPUT19), .A3(new_n487), .ZN(new_n532));
  OR2_X1    g346(.A1(KEYINPUT92), .A2(KEYINPUT19), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT92), .A2(KEYINPUT19), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n353), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n188), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n522), .B1(new_n511), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n530), .B1(new_n523), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n527), .B1(new_n539), .B2(KEYINPUT20), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n511), .A2(new_n520), .A3(new_n522), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n491), .A2(new_n492), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT88), .B(G143), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n509), .B(new_n502), .C1(new_n508), .C2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n493), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n542), .A2(new_n546), .B1(new_n536), .B2(new_n531), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n541), .B1(new_n547), .B2(new_n522), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT20), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n548), .A2(KEYINPUT94), .A3(new_n549), .A4(new_n530), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n539), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n540), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n477), .A2(new_n483), .A3(new_n526), .A4(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G214), .B1(G237), .B2(G902), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n384), .A2(new_n232), .A3(new_n386), .ZN(new_n557));
  INV_X1    g371(.A(G113), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT5), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n220), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n229), .B2(new_n559), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n222), .A2(new_n218), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n390), .A3(new_n383), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G122), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT82), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n557), .A2(new_n566), .A3(new_n563), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(KEYINPUT6), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n201), .A2(G125), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n243), .A2(new_n340), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n325), .A2(G224), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT84), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT83), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n573), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT6), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n564), .A2(new_n578), .A3(new_n567), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n570), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n566), .B(KEYINPUT8), .ZN(new_n581));
  INV_X1    g395(.A(new_n563), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n561), .A2(new_n562), .B1(new_n390), .B2(new_n383), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n569), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT85), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n574), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n571), .A2(new_n572), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n574), .A2(KEYINPUT7), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n589), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n571), .A2(new_n572), .A3(new_n591), .A4(new_n587), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n585), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G210), .B1(G237), .B2(G902), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT86), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n580), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n580), .B2(new_n594), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n556), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n555), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n320), .A2(new_n364), .A3(new_n442), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  INV_X1    g417(.A(G472), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n318), .B2(new_n270), .ZN(new_n605));
  INV_X1    g419(.A(new_n364), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n307), .A2(new_n310), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n313), .B1(new_n607), .B2(new_n315), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n442), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT33), .B1(new_n467), .B2(new_n468), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n458), .A2(new_n465), .ZN(new_n613));
  INV_X1    g427(.A(new_n466), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n458), .A2(new_n465), .A3(new_n466), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n359), .A2(new_n470), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n619), .A2(new_n620), .B1(new_n470), .B2(new_n473), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n554), .B2(new_n526), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n580), .A2(new_n594), .A3(new_n595), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n595), .B1(new_n580), .B2(new_n594), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n556), .B(new_n483), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n611), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NAND2_X1  g445(.A1(new_n475), .A2(new_n476), .ZN(new_n632));
  INV_X1    g446(.A(new_n472), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n511), .A2(new_n537), .ZN(new_n635));
  INV_X1    g449(.A(new_n522), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n529), .B1(new_n637), .B2(new_n541), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n551), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n551), .B1(new_n548), .B2(new_n530), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n639), .B1(new_n640), .B2(KEYINPUT97), .ZN(new_n641));
  OR3_X1    g455(.A1(new_n539), .A2(KEYINPUT97), .A3(new_n552), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n634), .A2(new_n643), .A3(new_n526), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n627), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n611), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NOR2_X1   g462(.A1(new_n605), .A2(new_n608), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n329), .A2(KEYINPUT36), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n349), .A2(new_n355), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n652), .A2(new_n484), .A3(new_n323), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n362), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n362), .A2(KEYINPUT98), .A3(new_n653), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n649), .A2(new_n442), .A3(new_n601), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  AND3_X1   g475(.A1(new_n634), .A2(new_n526), .A3(new_n643), .ZN(new_n662));
  INV_X1    g476(.A(new_n556), .ZN(new_n663));
  INV_X1    g477(.A(new_n626), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n624), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n479), .B1(new_n480), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n662), .A2(KEYINPUT99), .A3(new_n665), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n634), .A2(new_n643), .A3(new_n526), .A4(new_n668), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n556), .B1(new_n625), .B2(new_n626), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n320), .A2(new_n442), .A3(new_n658), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n193), .ZN(G30));
  NAND2_X1  g491(.A1(new_n553), .A2(new_n550), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT94), .B1(new_n638), .B2(new_n549), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n526), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n634), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n658), .A2(new_n663), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n305), .A2(new_n306), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n252), .A2(new_n253), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n265), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n484), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G472), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n314), .A2(new_n319), .A3(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n598), .A2(new_n599), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT38), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n682), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n667), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n442), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n190), .ZN(G45));
  NAND2_X1  g511(.A1(new_n619), .A2(new_n620), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n473), .A2(new_n470), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n680), .A2(new_n700), .A3(new_n668), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT100), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n680), .A2(new_n703), .A3(new_n700), .A4(new_n668), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n665), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n656), .A2(new_n657), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n608), .A2(KEYINPUT32), .B1(new_n297), .B2(G472), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n708), .B1(new_n709), .B2(new_n314), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n702), .A2(KEYINPUT101), .A3(new_n665), .A4(new_n704), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n707), .A2(new_n710), .A3(new_n442), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n675), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(KEYINPUT102), .A3(new_n711), .A4(new_n707), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  AOI21_X1  g532(.A(new_n408), .B1(new_n419), .B2(new_n369), .ZN(new_n719));
  INV_X1    g533(.A(new_n409), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n431), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n440), .B1(new_n721), .B2(new_n413), .ZN(new_n722));
  OAI21_X1  g536(.A(G469), .B1(new_n722), .B2(new_n359), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(KEYINPUT103), .A3(new_n441), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n725), .B(G469), .C1(new_n722), .C2(new_n359), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n367), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n606), .B1(new_n709), .B2(new_n314), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n628), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND2_X1  g545(.A1(new_n441), .A2(KEYINPUT103), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n407), .A2(new_n409), .B1(new_n368), .B2(new_n430), .ZN(new_n733));
  OAI22_X1  g547(.A1(new_n733), .A2(new_n414), .B1(new_n420), .B2(new_n439), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n435), .B1(new_n734), .B2(new_n270), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n726), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n366), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n320), .A2(new_n645), .A3(new_n364), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT104), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n727), .A2(new_n728), .A3(new_n741), .A4(new_n645), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  INV_X1    g558(.A(new_n555), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n727), .A2(new_n710), .A3(new_n745), .A4(new_n665), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  NAND3_X1  g561(.A1(new_n254), .A2(new_n258), .A3(new_n260), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n266), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n313), .B1(new_n607), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n605), .A2(new_n606), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n681), .A2(new_n672), .A3(new_n482), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n727), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  OAI211_X1 g568(.A(new_n366), .B(new_n665), .C1(new_n736), .C2(new_n737), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n605), .A2(new_n750), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n658), .A3(new_n704), .A4(new_n702), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n340), .ZN(G27));
  AOI21_X1  g573(.A(new_n703), .B1(new_n622), .B2(new_n668), .ZN(new_n760));
  INV_X1    g574(.A(new_n704), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n434), .A2(new_n441), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n434), .A2(KEYINPUT105), .A3(new_n441), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n598), .A2(new_n599), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n366), .A3(new_n556), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n762), .A2(new_n765), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT32), .B1(new_n318), .B2(new_n312), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n298), .B(new_n319), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n314), .A2(KEYINPUT106), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n364), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT42), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n434), .A2(KEYINPUT105), .A3(new_n441), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT105), .B1(new_n434), .B2(new_n441), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n778), .A3(new_n768), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n702), .A2(new_n704), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT42), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n728), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT107), .B(G131), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G33));
  XNOR2_X1  g599(.A(new_n671), .B(KEYINPUT108), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n779), .A2(new_n728), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n765), .A2(new_n766), .A3(new_n769), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n320), .A2(new_n364), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(KEYINPUT109), .A3(new_n786), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  NOR2_X1   g609(.A1(new_n680), .A2(new_n621), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(KEYINPUT110), .B2(KEYINPUT43), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n680), .B2(new_n621), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n708), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n649), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT44), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(KEYINPUT44), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n767), .A2(new_n556), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n433), .A2(KEYINPUT45), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n420), .B1(new_n409), .B2(new_n407), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n414), .B1(new_n429), .B2(new_n431), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(G469), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(G469), .A2(G902), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT46), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n441), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n813), .A2(KEYINPUT46), .A3(new_n814), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n367), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n692), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n807), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(new_n205), .ZN(G39));
  OR2_X1    g636(.A1(new_n819), .A2(KEYINPUT47), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n819), .A2(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n780), .A2(new_n320), .A3(new_n364), .A4(new_n805), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(KEYINPUT111), .B(G140), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(G42));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n830));
  NOR2_X1   g644(.A1(G952), .A2(G953), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n320), .A2(new_n628), .A3(new_n364), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n751), .A2(new_n752), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n738), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n320), .A2(new_n745), .A3(new_n658), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n755), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n837), .A2(new_n838), .A3(new_n743), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n771), .A2(new_n772), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n314), .A2(KEYINPUT106), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n709), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n779), .A2(new_n364), .A3(new_n762), .A4(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n843), .A2(KEYINPUT42), .B1(new_n792), .B2(new_n781), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n556), .B(new_n483), .C1(new_n598), .C2(new_n599), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(KEYINPUT115), .A3(new_n622), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n623), .B2(new_n845), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n609), .A2(new_n847), .A3(new_n442), .A4(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n471), .B1(new_n474), .B2(new_n469), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n554), .B(new_n526), .C1(new_n851), .C2(new_n472), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n649), .A2(new_n442), .A3(new_n364), .A4(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n850), .A2(new_n602), .A3(new_n659), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n643), .A2(new_n477), .A3(new_n526), .A4(new_n668), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n805), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n320), .A2(new_n857), .A3(new_n442), .A4(new_n658), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n790), .B2(new_n757), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n794), .A2(new_n844), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n838), .B1(new_n837), .B2(new_n743), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n839), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n777), .A2(new_n778), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n362), .A2(new_n653), .A3(new_n367), .A4(new_n667), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n681), .A2(new_n672), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n869), .A3(new_n865), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n867), .A2(new_n688), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n755), .A2(new_n757), .B1(new_n674), .B2(new_n675), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n717), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n872), .B1(new_n714), .B2(new_n716), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n871), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n863), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n602), .A2(new_n659), .A3(new_n854), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n708), .A2(new_n605), .A3(new_n750), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n779), .A2(new_n762), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n881), .A2(new_n850), .A3(new_n883), .A4(new_n858), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n783), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n746), .A2(new_n729), .A3(new_n753), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n742), .B2(new_n740), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n887), .A3(KEYINPUT53), .A4(new_n794), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n876), .B2(new_n878), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n880), .A2(KEYINPUT54), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n892));
  AND4_X1   g706(.A1(KEYINPUT52), .A2(new_n717), .A3(new_n871), .A4(new_n873), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(new_n877), .B2(new_n871), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n834), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n743), .A3(new_n746), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT114), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n837), .A2(new_n838), .A3(new_n743), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n794), .A3(new_n899), .A4(new_n885), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n892), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n863), .A2(new_n879), .A3(KEYINPUT53), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n890), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n724), .A2(new_n726), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n367), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n823), .A2(new_n824), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n479), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n797), .B2(new_n799), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(new_n751), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n806), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n907), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT51), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n690), .A2(new_n556), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n727), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT50), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n910), .A2(KEYINPUT50), .A3(new_n727), .A4(new_n916), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n727), .A2(new_n806), .ZN(new_n922));
  INV_X1    g736(.A(new_n909), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n882), .ZN(new_n925));
  INV_X1    g739(.A(new_n922), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n688), .A2(new_n606), .A3(new_n908), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n680), .A2(new_n700), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT120), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n914), .A2(new_n921), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n922), .A2(new_n775), .A3(new_n923), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT48), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n935), .A2(KEYINPUT48), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n926), .A2(new_n622), .A3(new_n927), .ZN(new_n938));
  INV_X1    g752(.A(new_n755), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n478), .B(G953), .C1(new_n939), .C2(new_n910), .ZN(new_n940));
  AND4_X1   g754(.A1(new_n936), .A2(new_n937), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n930), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n919), .A2(new_n920), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT119), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n943), .A2(KEYINPUT119), .A3(new_n944), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n907), .A2(new_n913), .A3(KEYINPUT118), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT118), .B1(new_n907), .B2(new_n913), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n942), .B1(new_n951), .B2(new_n915), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n831), .B1(new_n904), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n796), .A2(new_n364), .A3(new_n366), .A4(new_n556), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT112), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n955), .A2(new_n688), .A3(new_n690), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT49), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n905), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n724), .A2(KEYINPUT49), .A3(new_n726), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT113), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n830), .B1(new_n953), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n888), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n879), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n901), .A2(new_n891), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n901), .A2(new_n902), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n952), .B(new_n965), .C1(new_n966), .C2(new_n891), .ZN(new_n967));
  INV_X1    g781(.A(new_n831), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n961), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(KEYINPUT121), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n962), .A2(new_n971), .ZN(G75));
  AOI21_X1  g786(.A(new_n270), .B1(new_n901), .B2(new_n964), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n596), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT56), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n570), .A2(new_n579), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(new_n577), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT55), .Z(new_n978));
  AND3_X1   g792(.A1(new_n974), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n974), .B2(new_n975), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n325), .A2(G952), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(G51));
  OAI21_X1  g796(.A(KEYINPUT54), .B1(new_n880), .B2(new_n889), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(KEYINPUT122), .A3(new_n965), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n901), .A2(new_n964), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT122), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT54), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n814), .B(KEYINPUT57), .Z(new_n988));
  NAND3_X1  g802(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n734), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n973), .A2(G469), .A3(new_n808), .A4(new_n812), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(G54));
  NAND3_X1  g806(.A1(new_n973), .A2(KEYINPUT58), .A3(G475), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n993), .A2(new_n541), .A3(new_n637), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n541), .B2(new_n637), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n994), .A2(new_n995), .A3(new_n981), .ZN(G60));
  INV_X1    g810(.A(new_n981), .ZN(new_n997));
  NAND2_X1  g811(.A1(G478), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT59), .Z(new_n999));
  NOR2_X1   g813(.A1(new_n904), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n997), .B1(new_n1000), .B2(new_n619), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n999), .B1(new_n612), .B2(new_n618), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n984), .A2(new_n987), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1001), .A2(new_n1003), .ZN(G63));
  NAND2_X1  g818(.A1(G217), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT60), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n985), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n358), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n985), .A2(new_n652), .A3(new_n1006), .ZN(new_n1009));
  NOR2_X1   g823(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n981), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(G66));
  INV_X1    g828(.A(new_n481), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n325), .B1(new_n1015), .B2(G224), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n839), .A2(new_n862), .ZN(new_n1017));
  INV_X1    g831(.A(new_n855), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1016), .B1(new_n1019), .B2(new_n325), .ZN(new_n1020));
  INV_X1    g834(.A(G898), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n976), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1020), .B(new_n1022), .ZN(G69));
  AOI21_X1  g837(.A(new_n325), .B1(G227), .B2(G900), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n827), .A2(new_n794), .A3(new_n877), .ZN(new_n1025));
  NOR4_X1   g839(.A1(new_n820), .A2(new_n672), .A3(new_n681), .A4(new_n775), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n821), .A2(new_n1026), .A3(new_n783), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1025), .A2(new_n1027), .A3(new_n325), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n288), .B1(KEYINPUT30), .B2(new_n303), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n532), .A2(new_n535), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1028), .B(new_n1031), .C1(new_n666), .C2(new_n325), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n805), .B1(new_n623), .B2(new_n852), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n728), .A2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g849(.A(new_n827), .B1(new_n693), .B2(new_n1035), .C1(new_n820), .C2(new_n807), .ZN(new_n1036));
  INV_X1    g850(.A(new_n696), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(new_n877), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1041), .A2(G953), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1033), .B1(new_n1042), .B2(new_n1031), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1024), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(KEYINPUT124), .B1(new_n1042), .B2(new_n1031), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1024), .ZN(new_n1047));
  INV_X1    g861(.A(KEYINPUT124), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1031), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1048), .B(new_n1049), .C1(new_n1041), .C2(G953), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n1046), .A2(new_n1047), .A3(new_n1032), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1045), .A2(new_n1051), .ZN(G72));
  XOR2_X1   g866(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1053));
  NOR2_X1   g867(.A1(new_n604), .A2(new_n484), .ZN(new_n1054));
  XNOR2_X1  g868(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  INV_X1    g869(.A(new_n1019), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1055), .B1(new_n1041), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n291), .B(KEYINPUT127), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1058), .ZN(new_n1059));
  NOR3_X1   g873(.A1(new_n1057), .A2(new_n266), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g874(.A(new_n291), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n683), .B1(new_n266), .B2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g876(.A1(new_n966), .A2(new_n1055), .A3(new_n1062), .ZN(new_n1063));
  AND2_X1   g877(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1064));
  AOI21_X1  g878(.A(new_n1055), .B1(new_n1064), .B2(new_n1056), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1059), .A2(new_n266), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n997), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g881(.A1(new_n1060), .A2(new_n1063), .A3(new_n1067), .ZN(G57));
endmodule


