

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585;

  NOR2_X2 U320 ( .A1(n496), .A2(n447), .ZN(n448) );
  XNOR2_X2 U321 ( .A(KEYINPUT118), .B(n448), .ZN(n560) );
  XNOR2_X1 U322 ( .A(n353), .B(n352), .ZN(n354) );
  AND2_X1 U323 ( .A1(n563), .A2(n445), .ZN(n446) );
  XOR2_X1 U324 ( .A(n300), .B(n299), .Z(n288) );
  XOR2_X1 U325 ( .A(G29GAT), .B(KEYINPUT7), .Z(n289) );
  XNOR2_X1 U326 ( .A(KEYINPUT105), .B(KEYINPUT47), .ZN(n396) );
  XNOR2_X1 U327 ( .A(n301), .B(n288), .ZN(n302) );
  XNOR2_X1 U328 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U329 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(G85GAT), .B(G92GAT), .Z(n291) );
  XNOR2_X1 U332 ( .A(G99GAT), .B(G106GAT), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n305) );
  XOR2_X1 U334 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n293) );
  NAND2_X1 U335 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U337 ( .A(n294), .B(KEYINPUT11), .Z(n298) );
  XNOR2_X1 U338 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n289), .B(n295), .ZN(n360) );
  XNOR2_X1 U340 ( .A(G36GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n296), .B(KEYINPUT76), .ZN(n332) );
  XNOR2_X1 U342 ( .A(n360), .B(n332), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n303) );
  XOR2_X1 U344 ( .A(G43GAT), .B(G134GAT), .Z(n312) );
  XOR2_X1 U345 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XNOR2_X1 U346 ( .A(n312), .B(n422), .ZN(n301) );
  XOR2_X1 U347 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n300) );
  XNOR2_X1 U348 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n299) );
  XOR2_X1 U349 ( .A(n305), .B(n304), .Z(n555) );
  XOR2_X1 U350 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n307) );
  XNOR2_X1 U351 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U353 ( .A(G169GAT), .B(n308), .Z(n328) );
  XOR2_X1 U354 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n310) );
  XNOR2_X1 U355 ( .A(G190GAT), .B(KEYINPUT82), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U357 ( .A(n312), .B(n311), .Z(n314) );
  NAND2_X1 U358 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U360 ( .A(G176GAT), .B(KEYINPUT84), .Z(n316) );
  XNOR2_X1 U361 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U363 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U364 ( .A(G127GAT), .B(KEYINPUT80), .Z(n320) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n432) );
  XNOR2_X1 U367 ( .A(G99GAT), .B(G71GAT), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n321), .B(G120GAT), .ZN(n348) );
  XNOR2_X1 U369 ( .A(n432), .B(n348), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U371 ( .A(n328), .B(n324), .ZN(n496) );
  XOR2_X1 U372 ( .A(KEYINPUT21), .B(G218GAT), .Z(n326) );
  XNOR2_X1 U373 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U375 ( .A(G197GAT), .B(n327), .Z(n427) );
  XNOR2_X1 U376 ( .A(n328), .B(n427), .ZN(n339) );
  XOR2_X1 U377 ( .A(KEYINPUT73), .B(G64GAT), .Z(n330) );
  XNOR2_X1 U378 ( .A(G176GAT), .B(G92GAT), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U380 ( .A(G204GAT), .B(n331), .Z(n353) );
  XOR2_X1 U381 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n334) );
  XNOR2_X1 U382 ( .A(G8GAT), .B(n332), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U384 ( .A(n353), .B(n335), .Z(n337) );
  NAND2_X1 U385 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U387 ( .A(n339), .B(n338), .ZN(n518) );
  XNOR2_X1 U388 ( .A(KEYINPUT116), .B(n518), .ZN(n408) );
  XOR2_X1 U389 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n378) );
  AND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n378), .B(n340), .ZN(n342) );
  XNOR2_X1 U392 ( .A(G106GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n341), .B(G148GAT), .ZN(n415) );
  XNOR2_X1 U394 ( .A(n342), .B(n415), .ZN(n345) );
  INV_X1 U395 ( .A(n345), .ZN(n343) );
  NAND2_X1 U396 ( .A1(n343), .A2(KEYINPUT31), .ZN(n347) );
  INV_X1 U397 ( .A(KEYINPUT31), .ZN(n344) );
  NAND2_X1 U398 ( .A1(n345), .A2(n344), .ZN(n346) );
  NAND2_X1 U399 ( .A1(n347), .A2(n346), .ZN(n350) );
  XNOR2_X1 U400 ( .A(n348), .B(KEYINPUT72), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U402 ( .A(G85GAT), .B(G57GAT), .Z(n428) );
  XOR2_X1 U403 ( .A(n351), .B(n428), .Z(n355) );
  XNOR2_X1 U404 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n355), .B(n354), .ZN(n400) );
  XNOR2_X1 U406 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n400), .B(n356), .ZN(n548) );
  XNOR2_X1 U408 ( .A(G15GAT), .B(G8GAT), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n357), .B(G1GAT), .ZN(n382) );
  XOR2_X1 U410 ( .A(G141GAT), .B(G22GAT), .Z(n423) );
  XOR2_X1 U411 ( .A(n382), .B(n423), .Z(n359) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(G50GAT), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n364) );
  XOR2_X1 U414 ( .A(n360), .B(KEYINPUT29), .Z(n362) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U417 ( .A(n364), .B(n363), .Z(n372) );
  XOR2_X1 U418 ( .A(G197GAT), .B(G113GAT), .Z(n366) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(G36GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U421 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n368) );
  XNOR2_X1 U422 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n567) );
  NAND2_X1 U426 ( .A1(n548), .A2(n567), .ZN(n374) );
  INV_X1 U427 ( .A(KEYINPUT46), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n393) );
  XOR2_X1 U429 ( .A(G71GAT), .B(G127GAT), .Z(n376) );
  XNOR2_X1 U430 ( .A(G22GAT), .B(G183GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U432 ( .A(n378), .B(n377), .Z(n380) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U435 ( .A(n381), .B(KEYINPUT15), .Z(n384) );
  XNOR2_X1 U436 ( .A(n382), .B(KEYINPUT77), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n392) );
  XOR2_X1 U438 ( .A(G64GAT), .B(G78GAT), .Z(n386) );
  XNOR2_X1 U439 ( .A(G211GAT), .B(G155GAT), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U441 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n388) );
  XNOR2_X1 U442 ( .A(G57GAT), .B(KEYINPUT14), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U444 ( .A(n390), .B(n389), .Z(n391) );
  XNOR2_X1 U445 ( .A(n392), .B(n391), .ZN(n578) );
  NOR2_X1 U446 ( .A1(n393), .A2(n578), .ZN(n394) );
  XOR2_X1 U447 ( .A(n394), .B(KEYINPUT104), .Z(n395) );
  NOR2_X1 U448 ( .A1(n555), .A2(n395), .ZN(n397) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n405) );
  XNOR2_X1 U450 ( .A(n555), .B(KEYINPUT36), .ZN(n581) );
  NAND2_X1 U451 ( .A1(n581), .A2(n578), .ZN(n399) );
  XOR2_X1 U452 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n401) );
  BUF_X1 U454 ( .A(n400), .Z(n573) );
  NAND2_X1 U455 ( .A1(n401), .A2(n573), .ZN(n402) );
  XNOR2_X1 U456 ( .A(KEYINPUT106), .B(n402), .ZN(n403) );
  NOR2_X1 U457 ( .A1(n567), .A2(n403), .ZN(n404) );
  NOR2_X1 U458 ( .A1(n405), .A2(n404), .ZN(n407) );
  INV_X1 U459 ( .A(KEYINPUT48), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n543) );
  NAND2_X1 U461 ( .A1(n408), .A2(n543), .ZN(n409) );
  XNOR2_X1 U462 ( .A(n409), .B(KEYINPUT54), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n410), .B(KEYINPUT117), .ZN(n563) );
  XOR2_X1 U464 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n412) );
  NAND2_X1 U465 ( .A1(G228GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U467 ( .A(n413), .B(KEYINPUT88), .Z(n417) );
  XNOR2_X1 U468 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n414), .B(KEYINPUT2), .ZN(n429) );
  XNOR2_X1 U470 ( .A(n429), .B(n415), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U472 ( .A(G204GAT), .B(KEYINPUT22), .Z(n419) );
  XNOR2_X1 U473 ( .A(KEYINPUT23), .B(KEYINPUT89), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U475 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n464) );
  XOR2_X1 U479 ( .A(n428), .B(G162GAT), .Z(n431) );
  XNOR2_X1 U480 ( .A(G134GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U481 ( .A(n431), .B(n430), .ZN(n436) );
  XOR2_X1 U482 ( .A(n432), .B(KEYINPUT1), .Z(n434) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U485 ( .A(n436), .B(n435), .Z(n444) );
  XOR2_X1 U486 ( .A(G148GAT), .B(G120GAT), .Z(n438) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(G141GAT), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U489 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n440) );
  XNOR2_X1 U490 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U493 ( .A(n444), .B(n443), .ZN(n564) );
  INV_X1 U494 ( .A(n564), .ZN(n516) );
  NOR2_X1 U495 ( .A1(n464), .A2(n516), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n446), .B(KEYINPUT55), .ZN(n447) );
  NAND2_X1 U497 ( .A1(n555), .A2(n560), .ZN(n452) );
  XOR2_X1 U498 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n450) );
  INV_X1 U499 ( .A(G190GAT), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U501 ( .A(KEYINPUT101), .B(n548), .Z(n530) );
  NAND2_X1 U502 ( .A1(n530), .A2(n560), .ZN(n456) );
  XOR2_X1 U503 ( .A(G176GAT), .B(KEYINPUT56), .Z(n454) );
  XNOR2_X1 U504 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n476) );
  NAND2_X1 U507 ( .A1(n567), .A2(n573), .ZN(n487) );
  INV_X1 U508 ( .A(n578), .ZN(n457) );
  NOR2_X1 U509 ( .A1(n555), .A2(n457), .ZN(n458) );
  XOR2_X1 U510 ( .A(KEYINPUT16), .B(n458), .Z(n459) );
  XNOR2_X1 U511 ( .A(KEYINPUT79), .B(n459), .ZN(n474) );
  XOR2_X1 U512 ( .A(n518), .B(KEYINPUT27), .Z(n466) );
  NOR2_X1 U513 ( .A1(n466), .A2(n564), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT92), .ZN(n542) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(n464), .Z(n500) );
  NAND2_X1 U516 ( .A1(n542), .A2(n500), .ZN(n527) );
  XNOR2_X1 U517 ( .A(KEYINPUT85), .B(n496), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n527), .A2(n461), .ZN(n472) );
  INV_X1 U519 ( .A(n518), .ZN(n493) );
  NOR2_X1 U520 ( .A1(n496), .A2(n493), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n464), .A2(n462), .ZN(n463) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n463), .Z(n468) );
  NAND2_X1 U523 ( .A1(n464), .A2(n496), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT26), .ZN(n566) );
  NOR2_X1 U525 ( .A1(n566), .A2(n466), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n469), .A2(n516), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT93), .B(n470), .Z(n471) );
  NOR2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT94), .B(n473), .Z(n484) );
  NAND2_X1 U531 ( .A1(n474), .A2(n484), .ZN(n504) );
  NOR2_X1 U532 ( .A1(n487), .A2(n504), .ZN(n482) );
  NAND2_X1 U533 ( .A1(n482), .A2(n516), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U535 ( .A1(n482), .A2(n518), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n479) );
  INV_X1 U538 ( .A(n496), .ZN(n525) );
  NAND2_X1 U539 ( .A1(n482), .A2(n525), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT95), .Z(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  INV_X1 U543 ( .A(n500), .ZN(n521) );
  NAND2_X1 U544 ( .A1(n482), .A2(n521), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U546 ( .A1(n484), .A2(n581), .ZN(n485) );
  NOR2_X1 U547 ( .A1(n578), .A2(n485), .ZN(n486) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n486), .ZN(n515) );
  NOR2_X1 U549 ( .A1(n515), .A2(n487), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(KEYINPUT97), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(n501) );
  NOR2_X1 U552 ( .A1(n564), .A2(n501), .ZN(n492) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT98), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n490), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n501), .A2(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT99), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  NOR2_X1 U559 ( .A1(n501), .A2(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U562 ( .A(G43GAT), .B(n499), .Z(G1330GAT) );
  NOR2_X1 U563 ( .A1(n501), .A2(n500), .ZN(n502) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n506) );
  INV_X1 U566 ( .A(n567), .ZN(n503) );
  NAND2_X1 U567 ( .A1(n503), .A2(n530), .ZN(n514) );
  NOR2_X1 U568 ( .A1(n514), .A2(n504), .ZN(n510) );
  NAND2_X1 U569 ( .A1(n510), .A2(n516), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n510), .A2(n518), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n525), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(KEYINPUT102), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT103), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U577 ( .A1(n510), .A2(n521), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n513), .Z(G1335GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n522), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n522), .A2(n518), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n525), .A2(n522), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G99GAT), .B(n520), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT107), .Z(n529) );
  NAND2_X1 U591 ( .A1(n525), .A2(n543), .ZN(n526) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n537), .A2(n567), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT108), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U596 ( .A1(n537), .A2(n530), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT109), .Z(n535) );
  NAND2_X1 U600 ( .A1(n537), .A2(n578), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT111), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U604 ( .A1(n537), .A2(n555), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT110), .Z(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  XOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT113), .Z(n547) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n544), .A2(n566), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n545), .B(KEYINPUT112), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n567), .A2(n556), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U615 ( .A1(n556), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n553) );
  NAND2_X1 U619 ( .A1(n556), .A2(n578), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n567), .A2(n560), .ZN(n559) );
  XOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT119), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n578), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  NAND2_X1 U631 ( .A1(n563), .A2(n564), .ZN(n565) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n582) );
  NAND2_X1 U633 ( .A1(n582), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n577) );
  INV_X1 U639 ( .A(n573), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n582), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n582), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

