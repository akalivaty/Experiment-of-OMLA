//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n558, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT69), .B(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(new_n468), .A3(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n465), .A2(KEYINPUT70), .A3(new_n466), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n468), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n472), .B1(new_n481), .B2(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n467), .B(KEYINPUT71), .ZN(new_n487));
  INV_X1    g062(.A(G2105), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n486), .B1(new_n489), .B2(G136), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n487), .A2(new_n482), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n491), .A2(new_n492), .A3(G124), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n491), .B2(G124), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT73), .Z(G162));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n468), .A2(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n479), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n488), .A2(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT4), .A4(G138), .ZN(new_n503));
  NAND2_X1  g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n467), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n488), .A2(G102), .ZN(new_n507));
  NAND2_X1  g082(.A1(G114), .A2(G2105), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n464), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n499), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n515), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  OR3_X1    g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(G166));
  INV_X1    g106(.A(new_n521), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n535), .B(new_n536), .C1(new_n523), .C2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n533), .A2(new_n538), .ZN(G168));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n521), .A2(new_n540), .B1(new_n523), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n528), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  NOR2_X1   g120(.A1(new_n513), .A2(new_n514), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n532), .A2(G81), .B1(G43), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n528), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n548), .B(new_n552), .C1(new_n528), .C2(new_n549), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  XOR2_X1   g132(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n558));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n520), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT80), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n532), .A2(KEYINPUT79), .A3(G91), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n532), .A2(G91), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT78), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n523), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n547), .B(G53), .C1(KEYINPUT78), .C2(new_n572), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n570), .A2(new_n571), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n568), .A2(new_n569), .A3(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(new_n525), .ZN(new_n581));
  INV_X1    g156(.A(new_n530), .ZN(new_n582));
  NOR3_X1   g157(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(G303));
  AOI22_X1  g159(.A1(new_n532), .A2(G87), .B1(G49), .B2(new_n547), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n520), .A2(G74), .ZN(new_n586));
  NOR3_X1   g161(.A1(new_n586), .A2(KEYINPUT82), .A3(new_n528), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n588), .A2(KEYINPUT82), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(new_n547), .A2(G48), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n521), .B2(new_n592), .C1(new_n593), .C2(new_n528), .ZN(G305));
  AOI22_X1  g169(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n528), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT83), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n532), .A2(G85), .B1(G47), .B2(new_n547), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n547), .B(KEYINPUT84), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n532), .A2(G92), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n601), .A2(G54), .B1(new_n602), .B2(KEYINPUT10), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n520), .B(KEYINPUT81), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT85), .B(G66), .Z(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n528), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT86), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n606), .A2(new_n607), .ZN(new_n612));
  INV_X1    g187(.A(new_n609), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n614), .A2(new_n603), .A3(new_n615), .A4(new_n604), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n600), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n600), .B1(new_n617), .B2(G868), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NOR2_X1   g195(.A1(G286), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n570), .A2(new_n571), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n575), .A2(new_n576), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(new_n569), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n528), .B1(new_n564), .B2(new_n566), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n621), .B1(new_n626), .B2(new_n620), .ZN(G297));
  AOI21_X1  g202(.A(new_n621), .B1(new_n626), .B2(new_n620), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n617), .B1(new_n629), .B2(G860), .ZN(G148));
  INV_X1    g205(.A(new_n554), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n617), .A2(new_n629), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n632), .B1(new_n634), .B2(G868), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g211(.A(new_n479), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(new_n470), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT87), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n640), .A2(KEYINPUT13), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(KEYINPUT13), .B2(new_n640), .ZN(new_n644));
  OR3_X1    g219(.A1(new_n644), .A2(new_n641), .A3(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n641), .B2(new_n642), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n489), .A2(G135), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n491), .A2(G123), .ZN(new_n648));
  OAI221_X1 g223(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT88), .Z(G156));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT15), .B(G2435), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2427), .ZN(new_n658));
  INV_X1    g233(.A(G2430), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  XNOR2_X1  g248(.A(G2084), .B(G2090), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT17), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(new_n674), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(new_n671), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n674), .B2(new_n678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n672), .A2(new_n674), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n677), .B1(new_n682), .B2(KEYINPUT17), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n676), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n651), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(new_n642), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n700), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  MUX2_X1   g280(.A(G24), .B(G290), .S(G16), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n489), .A2(G131), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n491), .A2(G119), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g288(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n714));
  OAI221_X1 g289(.A(G2104), .B1(new_n713), .B2(new_n714), .C1(new_n468), .C2(G107), .ZN(new_n715));
  AND3_X1   g290(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT90), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT90), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G25), .A2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n709), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n716), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G29), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(new_n708), .C1(G25), .C2(G29), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n707), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n729));
  NOR2_X1   g304(.A1(G16), .A2(G23), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(G288), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT33), .B(G1976), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(G305), .A2(new_n732), .ZN(new_n736));
  OR2_X1    g311(.A1(G6), .A2(G16), .ZN(new_n737));
  AND3_X1   g312(.A1(new_n736), .A2(KEYINPUT92), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(KEYINPUT92), .B1(new_n736), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT32), .B(G1981), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT91), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n738), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n738), .B2(new_n739), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n735), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G16), .A2(G22), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G166), .B2(G16), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT94), .B(G1971), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n729), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n745), .A2(new_n729), .A3(new_n749), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n728), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT36), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT28), .B1(new_n720), .B2(G26), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n720), .A2(KEYINPUT28), .A3(G26), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n491), .A2(G128), .ZN(new_n757));
  OAI21_X1  g332(.A(KEYINPUT95), .B1(G104), .B2(G2105), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(KEYINPUT95), .A2(G104), .A3(G2105), .ZN(new_n760));
  OAI221_X1 g335(.A(G2104), .B1(new_n759), .B2(new_n760), .C1(new_n468), .C2(G116), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n489), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n755), .B(new_n756), .C1(new_n764), .C2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n732), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n732), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1966), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n765), .A2(new_n766), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n732), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G171), .B2(new_n732), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G1961), .Z(new_n774));
  NAND4_X1  g349(.A1(new_n767), .A2(new_n770), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n720), .A2(G32), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n489), .A2(G141), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n491), .A2(G129), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT26), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n782), .A2(new_n783), .B1(G105), .B2(new_n470), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n778), .A2(new_n779), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n776), .B(new_n777), .C1(new_n786), .C2(new_n720), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT101), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n732), .A2(G19), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n554), .B2(new_n732), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1341), .ZN(new_n791));
  NOR2_X1   g366(.A1(G27), .A2(G29), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G164), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(KEYINPUT24), .A2(G34), .ZN(new_n796));
  NAND2_X1  g371(.A1(KEYINPUT24), .A2(G34), .ZN(new_n797));
  AOI21_X1  g372(.A(G29), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G160), .B2(G29), .ZN(new_n799));
  INV_X1    g374(.A(G2084), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n775), .A2(new_n788), .A3(new_n791), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(G162), .A2(G29), .ZN(new_n804));
  OR2_X1    g379(.A1(G29), .A2(G35), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n804), .A2(KEYINPUT29), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(KEYINPUT29), .B1(new_n804), .B2(new_n805), .ZN(new_n808));
  OAI21_X1  g383(.A(G2090), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n617), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G4), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G1348), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n732), .A2(G20), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT23), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n626), .B2(new_n732), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(G1956), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT31), .B(G11), .Z(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT30), .B(G28), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n720), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n650), .B2(new_n720), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n776), .B1(new_n786), .B2(new_n720), .ZN(new_n823));
  INV_X1    g398(.A(new_n777), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n817), .A2(G1956), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n813), .A2(new_n814), .A3(new_n818), .A4(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n808), .ZN(new_n829));
  INV_X1    g404(.A(G2090), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n829), .A2(new_n830), .A3(new_n806), .ZN(new_n831));
  AND4_X1   g406(.A1(new_n803), .A2(new_n809), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT25), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n487), .A2(new_n488), .ZN(new_n835));
  INV_X1    g410(.A(G139), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT96), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n637), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n468), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(KEYINPUT97), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT97), .B1(new_n838), .B2(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT98), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n838), .A2(new_n840), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n848), .A3(new_n841), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n720), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n720), .A2(G33), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G2072), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n851), .B1(new_n850), .B2(new_n853), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n754), .A2(new_n832), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n854), .A2(new_n856), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n861), .B2(new_n855), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(KEYINPUT100), .A3(G2072), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(G311));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n832), .A2(new_n857), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n754), .A3(new_n866), .ZN(G150));
  NAND2_X1  g442(.A1(new_n617), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  INV_X1    g444(.A(G93), .ZN(new_n870));
  INV_X1    g445(.A(G55), .ZN(new_n871));
  OAI22_X1  g446(.A1(new_n521), .A2(new_n870), .B1(new_n523), .B2(new_n871), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(new_n528), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n554), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n550), .A2(new_n875), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n869), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n881));
  AOI21_X1  g456(.A(G860), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(G860), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT37), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G145));
  NAND2_X1  g461(.A1(new_n764), .A2(new_n511), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n764), .A2(new_n511), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n786), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n762), .A2(new_n763), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G164), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n785), .A3(new_n887), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n844), .A3(new_n849), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n890), .B(new_n893), .C1(new_n843), .C2(new_n842), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n491), .A2(G130), .ZN(new_n898));
  OAI221_X1 g473(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n489), .B2(G142), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n489), .A2(new_n901), .A3(G142), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n717), .A2(new_n639), .A3(new_n718), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n639), .B1(new_n717), .B2(new_n718), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n719), .A2(new_n640), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n725), .A2(new_n639), .ZN(new_n910));
  INV_X1    g485(.A(new_n905), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n897), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(G162), .A2(G160), .ZN(new_n914));
  NAND2_X1  g489(.A1(G162), .A2(G160), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n650), .B(KEYINPUT102), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n908), .A2(new_n912), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n895), .A2(new_n920), .A3(new_n896), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n913), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n895), .A2(new_n920), .A3(new_n896), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n896), .B2(new_n895), .ZN(new_n924));
  OAI22_X1  g499(.A1(new_n923), .A2(new_n924), .B1(new_n918), .B2(new_n917), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(G395));
  XNOR2_X1  g504(.A(G290), .B(G288), .ZN(new_n930));
  XNOR2_X1  g505(.A(G303), .B(G305), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n877), .A2(new_n878), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n634), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n879), .A2(new_n633), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(G299), .B1(new_n610), .B2(new_n605), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n626), .A2(new_n614), .A3(new_n604), .A4(new_n603), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n939), .B(KEYINPUT41), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n934), .A3(new_n935), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n942), .B1(new_n941), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n932), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  INV_X1    g524(.A(new_n932), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n945), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n951), .A3(G868), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT105), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n948), .A2(new_n951), .A3(new_n954), .A4(G868), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n876), .A2(new_n620), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G295));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G331));
  XNOR2_X1  g533(.A(G301), .B(G168), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n933), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n959), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n877), .A2(new_n961), .A3(new_n878), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n943), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n940), .A3(new_n962), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n932), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n926), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n932), .B1(new_n964), .B2(new_n965), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT43), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT106), .B(KEYINPUT43), .C1(new_n967), .C2(new_n968), .ZN(new_n973));
  INV_X1    g548(.A(new_n967), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n939), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n976), .B(new_n963), .C1(new_n943), .C2(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n965), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n950), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n975), .B1(new_n974), .B2(new_n979), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n967), .A2(KEYINPUT43), .A3(new_n968), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT44), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n511), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(G160), .A2(G40), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n764), .B(new_n766), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1996), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n786), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n991), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n995), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(new_n785), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT109), .Z(new_n1000));
  NOR2_X1   g575(.A1(new_n719), .A2(new_n709), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n725), .A2(new_n708), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n991), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  AND2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G290), .A2(G1986), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n991), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT108), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n477), .A2(new_n478), .A3(G138), .A4(new_n468), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n509), .B1(new_n1011), .B2(new_n497), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n1012), .B2(new_n506), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G40), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1016), .B(new_n472), .C1(new_n481), .C2(new_n482), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1010), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT118), .B1(new_n1018), .B2(G2067), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT111), .B(G1384), .C1(new_n1012), .C2(new_n506), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1014), .B1(new_n511), .B2(new_n986), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n766), .A4(new_n1017), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1010), .A2(new_n1026), .A3(new_n1015), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n990), .B1(KEYINPUT50), .B2(new_n987), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1348), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n617), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n611), .A2(new_n616), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n812), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1031), .A2(new_n1033), .A3(new_n1019), .A4(new_n1024), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT60), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1031), .A2(KEYINPUT60), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(new_n1017), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n989), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT120), .B(G1996), .Z(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT58), .B(G1341), .Z(new_n1046));
  AND2_X1   g621(.A1(new_n1018), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1040), .B(new_n554), .C1(new_n1045), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1041), .A2(new_n1017), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1013), .A2(KEYINPUT45), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1044), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1051), .A2(new_n1052), .B1(new_n1018), .B2(new_n1046), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT59), .B1(new_n1053), .B2(new_n631), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1038), .A2(new_n1039), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(KEYINPUT57), .C1(new_n624), .C2(new_n625), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n568), .A2(new_n569), .A3(new_n577), .A4(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1956), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1064), .B2(new_n990), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1051), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1010), .A2(KEYINPUT50), .A3(new_n1015), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1063), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n990), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1061), .B(new_n1067), .C1(new_n1071), .C2(G1956), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1056), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1067), .B1(new_n1071), .B2(G1956), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1061), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(KEYINPUT61), .A3(new_n1072), .ZN(new_n1078));
  AND4_X1   g653(.A1(new_n1036), .A2(new_n1055), .A3(new_n1074), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1037), .A2(new_n617), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1073), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1030), .A2(new_n1077), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(KEYINPUT119), .A3(new_n1072), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n989), .A2(new_n794), .A3(new_n1017), .A4(new_n1041), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n794), .A2(KEYINPUT53), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n987), .B2(new_n988), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n990), .A2(KEYINPUT123), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1017), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .A4(new_n1041), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1017), .B1(new_n1013), .B2(new_n1026), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1089), .B(new_n1095), .C1(new_n1097), .C2(G1961), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G171), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT54), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1089), .B(G301), .C1(new_n1097), .C2(G1961), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n988), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1102), .A2(KEYINPUT122), .A3(new_n1042), .A4(new_n794), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n794), .A3(new_n1042), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1088), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1101), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT124), .B1(new_n1100), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT53), .B1(new_n1051), .B2(new_n794), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1961), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1109), .A2(new_n1110), .A3(G171), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(KEYINPUT53), .A3(new_n1103), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1098), .B2(G171), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1098), .A2(G171), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1089), .B1(new_n1097), .B2(G1961), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1121), .B2(G301), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1108), .A2(new_n1118), .B1(new_n1122), .B2(new_n1115), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT55), .ZN(new_n1125));
  INV_X1    g700(.A(G8), .ZN(new_n1126));
  NOR3_X1   g701(.A1(G166), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1971), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1071), .A2(new_n830), .B1(new_n1131), .B2(new_n1043), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1126), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1071), .A2(new_n830), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1043), .A2(new_n1131), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT116), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1130), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n585), .B(G1976), .C1(new_n587), .C2(new_n589), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT112), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1018), .A2(new_n1141), .A3(G8), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1018), .B2(G8), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT52), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1027), .A2(new_n830), .A3(new_n1028), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1136), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(G8), .A3(new_n1130), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT113), .B(G1976), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT52), .B1(G288), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1140), .B(new_n1150), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT114), .B(G86), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n591), .B1(new_n521), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n593), .A2(new_n528), .ZN(new_n1154));
  OAI21_X1  g729(.A(G1981), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(G305), .B2(G1981), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT115), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1157), .A2(KEYINPUT49), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(KEYINPUT49), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1158), .B(new_n1159), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1145), .A2(new_n1148), .A3(new_n1151), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1139), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(G286), .A2(G8), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1163), .A2(KEYINPUT121), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(KEYINPUT51), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1049), .B1(new_n1166), .B2(new_n988), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1167), .A2(G1966), .B1(new_n1032), .B2(G2084), .ZN(new_n1168));
  OAI211_X1 g743(.A(G8), .B(new_n1165), .C1(new_n1168), .C2(G286), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1027), .A2(new_n800), .A3(new_n1028), .ZN(new_n1170));
  AOI21_X1  g745(.A(G1966), .B1(new_n1102), .B2(new_n1042), .ZN(new_n1171));
  OAI21_X1  g746(.A(G8), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1165), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1172), .A2(new_n1163), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1168), .A2(G8), .A3(G286), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1169), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1123), .A2(new_n1124), .A3(new_n1162), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1120), .ZN(new_n1178));
  AOI21_X1  g753(.A(G301), .B1(new_n1113), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1098), .A2(G171), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1115), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1114), .A2(new_n1117), .A3(new_n1116), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1117), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1160), .A2(new_n1151), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT52), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1020), .A2(new_n1021), .A3(new_n990), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT112), .B1(new_n1187), .B2(new_n1126), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1018), .A2(new_n1141), .A3(G8), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1186), .B1(new_n1190), .B2(new_n1140), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1126), .B(new_n1129), .C1(new_n1136), .C2(new_n1146), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1185), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1135), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(G8), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1129), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1193), .A2(new_n1197), .A3(new_n1176), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT125), .B1(new_n1184), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1086), .B1(new_n1177), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1176), .A2(KEYINPUT62), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1113), .A2(new_n1178), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(G171), .ZN(new_n1205));
  NOR3_X1   g780(.A1(new_n1139), .A2(new_n1161), .A3(new_n1205), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1176), .A2(KEYINPUT62), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1176), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1203), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1130), .B1(new_n1147), .B2(G8), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1168), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1211));
  OR3_X1    g786(.A1(new_n1161), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1168), .A2(G8), .A3(G168), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1139), .A2(new_n1161), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1212), .B1(new_n1214), .B2(KEYINPUT63), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1185), .A2(new_n1191), .A3(new_n1148), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1160), .ZN(new_n1217));
  OR2_X1    g792(.A1(G288), .A2(G1976), .ZN(new_n1218));
  OAI22_X1  g793(.A1(new_n1217), .A2(new_n1218), .B1(G1981), .B2(G305), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1216), .B1(new_n1190), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1209), .A2(new_n1215), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1009), .B1(new_n1200), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT47), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n992), .B(KEYINPUT110), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n786), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n991), .ZN(new_n1226));
  XOR2_X1   g801(.A(new_n998), .B(KEYINPUT46), .Z(new_n1227));
  INV_X1    g802(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1223), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  AOI211_X1 g804(.A(KEYINPUT47), .B(new_n1227), .C1(new_n1225), .C2(new_n991), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1006), .A2(new_n991), .ZN(new_n1231));
  XOR2_X1   g806(.A(new_n1231), .B(KEYINPUT48), .Z(new_n1232));
  OAI22_X1  g807(.A1(new_n1229), .A2(new_n1230), .B1(new_n1004), .B2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1234), .B1(G2067), .B2(new_n764), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1233), .B1(new_n991), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1222), .A2(new_n1236), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g812(.A1(new_n971), .A2(new_n973), .A3(new_n980), .ZN(new_n1239));
  NOR2_X1   g813(.A1(G401), .A2(new_n461), .ZN(new_n1240));
  NAND3_X1  g814(.A1(new_n1240), .A2(new_n686), .A3(new_n704), .ZN(new_n1241));
  XNOR2_X1  g815(.A(new_n1241), .B(KEYINPUT127), .ZN(new_n1242));
  AND3_X1   g816(.A1(new_n1239), .A2(new_n927), .A3(new_n1242), .ZN(G308));
  NAND3_X1  g817(.A1(new_n1239), .A2(new_n927), .A3(new_n1242), .ZN(G225));
endmodule


