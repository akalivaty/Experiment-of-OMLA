//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1206, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n210), .B(new_n211), .C1(new_n202), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G50), .B2(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n209), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G20), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n224), .B(new_n227), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n212), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT67), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  INV_X1    g0043(.A(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT68), .B(G87), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G226), .A2(G1698), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(new_n212), .B2(G1698), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n256), .A2(new_n258), .B1(G33), .B2(G97), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  OAI211_X1 g0060(.A(G1), .B(G13), .C1(new_n254), .C2(new_n260), .ZN(new_n261));
  OR3_X1    g0061(.A1(new_n259), .A2(KEYINPUT73), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n261), .A2(new_n264), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G238), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT73), .B1(new_n259), .B2(new_n261), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n262), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT13), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n262), .A2(new_n272), .A3(new_n268), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G200), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT74), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n228), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n254), .A2(G20), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n280), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  XOR2_X1   g0084(.A(new_n284), .B(KEYINPUT11), .Z(new_n285));
  AOI21_X1  g0085(.A(new_n278), .B1(new_n263), .B2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(KEYINPUT70), .A3(G68), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n288));
  OR3_X1    g0088(.A1(new_n288), .A2(KEYINPUT12), .A3(G68), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(KEYINPUT70), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G68), .ZN(new_n291));
  XOR2_X1   g0091(.A(KEYINPUT75), .B(KEYINPUT12), .Z(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n285), .A2(new_n287), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n271), .A2(G190), .A3(new_n273), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT74), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n274), .A2(new_n296), .A3(G200), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n276), .A2(new_n294), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n286), .A2(KEYINPUT70), .A3(G77), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT71), .Z(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n303));
  INV_X1    g0103(.A(new_n280), .ZN(new_n304));
  XOR2_X1   g0104(.A(KEYINPUT15), .B(G87), .Z(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n290), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n307), .A2(new_n278), .B1(new_n215), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n267), .A2(G244), .ZN(new_n312));
  INV_X1    g0112(.A(G1698), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n256), .A2(G232), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n314), .B(new_n315), .C1(new_n220), .C2(new_n256), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n317));
  AOI211_X1 g0117(.A(new_n266), .B(new_n312), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G190), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n311), .B(new_n319), .C1(new_n320), .C2(new_n318), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(new_n310), .C1(G169), .C2(new_n318), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(new_n274), .B2(G169), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  AOI211_X1 g0128(.A(KEYINPUT14), .B(new_n328), .C1(new_n271), .C2(new_n273), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n274), .A2(new_n322), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n298), .B(new_n325), .C1(new_n331), .C2(new_n294), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(G58), .B(G68), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(G20), .B1(G159), .B2(new_n282), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n252), .A2(G33), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G20), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT78), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n255), .B1(new_n342), .B2(new_n254), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(G20), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n341), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n252), .A2(KEYINPUT76), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT76), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n350), .A3(new_n254), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n337), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(KEYINPUT78), .A3(new_n345), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n340), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n335), .B1(new_n354), .B2(new_n203), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(new_n350), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n253), .B1(new_n358), .B2(G33), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT7), .B1(new_n359), .B2(G20), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n336), .B1(new_n342), .B2(new_n254), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n344), .A3(new_n339), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(G68), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT16), .A3(new_n335), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n363), .A2(KEYINPUT77), .A3(KEYINPUT16), .A4(new_n335), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n357), .A2(new_n278), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n252), .A2(KEYINPUT76), .ZN(new_n370));
  OAI21_X1  g0170(.A(G33), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(G223), .A2(G1698), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n313), .A2(G226), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n371), .A2(new_n336), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n374), .A2(KEYINPUT80), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT80), .B1(new_n374), .B2(new_n375), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n376), .A2(new_n377), .A3(new_n261), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n266), .B1(new_n267), .B2(G232), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n320), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n377), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n374), .A2(KEYINPUT80), .A3(new_n375), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n317), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n379), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n301), .A2(new_n288), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n286), .B2(new_n301), .ZN(new_n389));
  XOR2_X1   g0189(.A(new_n389), .B(KEYINPUT79), .Z(new_n390));
  NAND3_X1  g0190(.A1(new_n368), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n368), .A2(new_n387), .A3(KEYINPUT17), .A4(new_n390), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n366), .A2(new_n278), .A3(new_n367), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n355), .A2(new_n356), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n378), .B2(new_n380), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n384), .A2(G179), .A3(new_n379), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n397), .A2(KEYINPUT18), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT18), .B1(new_n397), .B2(new_n400), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n393), .B(new_n394), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT81), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n266), .B1(new_n267), .B2(G226), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n405), .A2(KEYINPUT69), .ZN(new_n406));
  NOR2_X1   g0206(.A1(G222), .A2(G1698), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n313), .A2(G223), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n256), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n409), .B(new_n317), .C1(G77), .C2(new_n256), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(KEYINPUT69), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G200), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n286), .A2(G50), .ZN(new_n414));
  INV_X1    g0214(.A(new_n288), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n201), .ZN(new_n416));
  INV_X1    g0216(.A(G150), .ZN(new_n417));
  INV_X1    g0217(.A(new_n282), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n301), .A2(new_n304), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(G20), .B2(new_n204), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n414), .B(new_n416), .C1(new_n420), .C2(new_n279), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n421), .A2(KEYINPUT9), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(KEYINPUT9), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n413), .B1(new_n385), .B2(new_n412), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT10), .ZN(new_n425));
  OR3_X1    g0225(.A1(new_n424), .A2(KEYINPUT72), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(KEYINPUT72), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(KEYINPUT72), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n412), .A2(G179), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n412), .A2(new_n328), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n421), .A3(new_n432), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n426), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n393), .A2(new_n394), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n397), .A2(new_n400), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n397), .A2(KEYINPUT18), .A3(new_n400), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT81), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n435), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AND4_X1   g0242(.A1(new_n333), .A2(new_n404), .A3(new_n434), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT5), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G41), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n263), .A2(G45), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n261), .B(G270), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT88), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n254), .B1(new_n348), .B2(new_n350), .ZN(new_n451));
  NOR2_X1   g0251(.A1(G257), .A2(G1698), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n313), .A2(G264), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n451), .A2(new_n253), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G303), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n256), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n317), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n448), .A2(new_n265), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n444), .A3(new_n446), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n339), .C1(G33), .C2(new_n244), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT84), .B(G116), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n278), .B(new_n462), .C1(new_n463), .C2(new_n339), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT20), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n308), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n278), .B1(new_n263), .B2(G33), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n290), .A2(G116), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n460), .A2(new_n471), .A3(G169), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT21), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n460), .A2(new_n471), .A3(KEYINPUT21), .A4(G169), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n460), .A2(new_n322), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n471), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n460), .A2(G200), .ZN(new_n479));
  INV_X1    g0279(.A(new_n471), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n479), .B(new_n480), .C1(new_n385), .C2(new_n460), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n476), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n217), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n371), .A2(new_n339), .A3(new_n336), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n339), .A2(G87), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n483), .B1(new_n338), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n463), .A2(new_n280), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n339), .A2(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT23), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n485), .A2(new_n490), .A3(new_n492), .A4(new_n487), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n279), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n469), .A2(new_n288), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT25), .B1(new_n415), .B2(new_n220), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n415), .A2(KEYINPUT25), .A3(new_n220), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n498), .A2(G107), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n218), .A2(new_n313), .ZN(new_n504));
  INV_X1    g0304(.A(G257), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G1698), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n371), .A2(new_n336), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G294), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n261), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n261), .B1(new_n447), .B2(new_n448), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n221), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n328), .B1(new_n512), .B2(new_n459), .ZN(new_n513));
  INV_X1    g0313(.A(new_n459), .ZN(new_n514));
  NOR4_X1   g0314(.A1(new_n509), .A2(new_n322), .A3(new_n514), .A4(new_n511), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n496), .A2(new_n503), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n507), .A2(new_n508), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n317), .ZN(new_n518));
  INV_X1    g0318(.A(new_n511), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(new_n385), .A3(new_n459), .A4(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n509), .A2(new_n514), .A3(new_n511), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(G200), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n278), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n525), .A3(new_n502), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT89), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n493), .A2(new_n495), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n503), .B1(new_n529), .B2(new_n278), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT89), .B1(new_n530), .B2(new_n522), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n516), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G238), .A2(G1698), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n313), .A2(G244), .ZN(new_n534));
  NOR4_X1   g0334(.A1(new_n451), .A2(new_n253), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n463), .A2(G33), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n317), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT85), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n261), .A2(new_n448), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n540), .A2(new_n218), .B1(new_n265), .B2(new_n448), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n533), .ZN(new_n544));
  INV_X1    g0344(.A(new_n534), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n371), .A2(new_n336), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n261), .B1(new_n546), .B2(new_n536), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT85), .B1(new_n547), .B2(new_n541), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(new_n548), .A3(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n359), .A2(new_n339), .A3(G68), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT19), .B1(new_n280), .B2(G97), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n217), .ZN(new_n553));
  NAND3_X1  g0353(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n339), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n279), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n308), .B2(new_n306), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n498), .A2(G87), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n543), .A2(new_n548), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT87), .B1(new_n561), .B2(G190), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT87), .ZN(new_n563));
  AOI211_X1 g0363(.A(new_n563), .B(new_n385), .C1(new_n543), .C2(new_n548), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n549), .B(new_n560), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n498), .A2(new_n305), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n558), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT86), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n561), .A2(new_n322), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n543), .A2(new_n548), .A3(new_n328), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n558), .A2(new_n571), .A3(new_n566), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n532), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n459), .B1(new_n510), .B2(new_n505), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT83), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(KEYINPUT83), .B(new_n459), .C1(new_n510), .C2(new_n505), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n336), .A2(new_n337), .A3(G250), .A4(G1698), .ZN(new_n582));
  AND2_X1   g0382(.A1(KEYINPUT4), .A2(G244), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n336), .A2(new_n337), .A3(new_n583), .A4(new_n313), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n584), .A3(new_n461), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NOR4_X1   g0386(.A1(new_n451), .A2(new_n216), .A3(G1698), .A4(new_n253), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(KEYINPUT4), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT82), .B1(new_n588), .B2(new_n317), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n371), .A2(G244), .A3(new_n313), .A4(new_n336), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n592), .A2(new_n593), .A3(new_n261), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n581), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n580), .B1(new_n317), .B2(new_n588), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(G200), .B1(new_n596), .B2(G190), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n288), .A2(G97), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n497), .A2(new_n244), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n244), .A2(new_n220), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n603), .B2(new_n552), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n220), .A2(KEYINPUT6), .A3(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n340), .ZN(new_n609));
  AOI211_X1 g0409(.A(new_n341), .B(new_n346), .C1(new_n351), .C2(new_n337), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT78), .B1(new_n352), .B2(new_n345), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n608), .B1(new_n612), .B2(G107), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n599), .B(new_n601), .C1(new_n613), .C2(new_n279), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n597), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n588), .A2(new_n317), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n581), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n328), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n322), .B(new_n581), .C1(new_n589), .C2(new_n594), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n614), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n443), .A2(new_n482), .A3(new_n575), .A4(new_n622), .ZN(G372));
  XNOR2_X1  g0423(.A(new_n538), .B(KEYINPUT90), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n542), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n328), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n569), .A3(new_n567), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT91), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT91), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n626), .A2(new_n629), .A3(new_n569), .A4(new_n567), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n526), .A2(new_n527), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n530), .A2(KEYINPUT89), .A3(new_n522), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n516), .A2(new_n478), .A3(new_n475), .A4(new_n474), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n621), .A3(new_n616), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n625), .A2(G200), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n637), .B(new_n560), .C1(new_n562), .C2(new_n564), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n627), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n631), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n614), .A2(new_n619), .A3(new_n620), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n565), .A2(new_n573), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n638), .A2(new_n644), .A3(new_n641), .A4(new_n627), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n443), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n433), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n331), .A2(new_n294), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT92), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n324), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n324), .A2(new_n651), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n650), .B1(new_n298), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n435), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n440), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n426), .A2(new_n430), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n649), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n648), .A2(new_n659), .ZN(G369));
  NAND2_X1  g0460(.A1(new_n339), .A2(G13), .ZN(new_n661));
  OR3_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .A3(G1), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT27), .B1(new_n661), .B2(G1), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT93), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT93), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n482), .B1(new_n480), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n476), .A2(new_n478), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n471), .A3(new_n669), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n516), .A2(new_n670), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT94), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n634), .B(new_n516), .C1(new_n530), .C2(new_n670), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n672), .A2(new_n670), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n679), .B2(new_n680), .ZN(new_n684));
  INV_X1    g0484(.A(new_n516), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n669), .B(KEYINPUT95), .Z(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n225), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n553), .A2(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n231), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n687), .B1(new_n640), .B2(new_n646), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT26), .B1(new_n639), .B2(new_n621), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n565), .A2(new_n641), .A3(new_n644), .A4(new_n573), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT29), .B(new_n670), .C1(new_n702), .C2(new_n640), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n575), .A2(new_n482), .A3(new_n622), .A4(new_n687), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n477), .A2(new_n596), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n561), .A2(new_n512), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT30), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n512), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n543), .B2(new_n548), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n477), .A3(new_n596), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n521), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n595), .A2(KEYINPUT96), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT96), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n588), .A2(KEYINPUT82), .A3(new_n317), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n593), .B1(new_n592), .B2(new_n261), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n580), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n715), .B1(new_n718), .B2(new_n521), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n714), .A2(new_n719), .A3(new_n322), .A4(new_n625), .ZN(new_n720));
  INV_X1    g0520(.A(new_n460), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n712), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n669), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n704), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n699), .A2(new_n703), .B1(G330), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n696), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n339), .A2(new_n322), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n731), .A2(G190), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G311), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n320), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G20), .A3(G190), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n733), .A2(new_n734), .B1(new_n736), .B2(new_n455), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n731), .A2(new_n320), .A3(G190), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT33), .B(G317), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(G20), .A3(new_n385), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT99), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G283), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G20), .A3(new_n385), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G329), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n339), .B1(new_n748), .B2(G190), .ZN(new_n752));
  INV_X1    g0552(.A(G294), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n338), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n730), .A2(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G200), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n754), .B1(G322), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n740), .A2(new_n747), .A3(new_n751), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n755), .A2(new_n320), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n759), .A2(G326), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n746), .A2(G107), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(G58), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n750), .A2(G159), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT32), .ZN(new_n764));
  INV_X1    g0564(.A(new_n736), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n738), .A2(G68), .B1(G87), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n761), .A2(new_n762), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n752), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n759), .A2(G50), .B1(G97), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n338), .B1(new_n763), .B2(KEYINPUT32), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(new_n215), .C2(new_n733), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n758), .A2(new_n760), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n228), .B1(G20), .B2(new_n328), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n773), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n225), .A2(G355), .A3(new_n256), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n690), .A2(new_n359), .ZN(new_n779));
  INV_X1    g0579(.A(G45), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n250), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n231), .A2(G45), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n778), .B1(G116), .B2(new_n225), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n772), .A2(new_n773), .B1(new_n777), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n661), .B(KEYINPUT98), .Z(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G45), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G1), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n691), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT100), .Z(new_n790));
  INV_X1    g0590(.A(new_n776), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n674), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n677), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n675), .A2(KEYINPUT97), .A3(new_n676), .ZN(new_n794));
  INV_X1    g0594(.A(new_n788), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(KEYINPUT97), .B1(new_n675), .B2(new_n676), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(G396));
  INV_X1    g0598(.A(KEYINPUT102), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n669), .A2(new_n310), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n325), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n310), .B(new_n669), .C1(new_n652), .C2(new_n653), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n321), .A2(new_n324), .A3(new_n800), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(KEYINPUT102), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n697), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n687), .B(new_n805), .C1(new_n640), .C2(new_n646), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT104), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n727), .A2(G330), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n810), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n795), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n806), .A2(new_n774), .ZN(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  INV_X1    g0618(.A(new_n738), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n818), .A2(new_n819), .B1(new_n733), .B2(new_n467), .ZN(new_n820));
  INV_X1    g0620(.A(new_n759), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n821), .A2(new_n455), .B1(new_n220), .B2(new_n736), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n256), .B1(new_n746), .B2(G87), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n756), .A2(G294), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n768), .A2(G97), .B1(new_n750), .B2(G311), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n732), .A2(G159), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n756), .A2(G143), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n831), .B2(new_n821), .C1(new_n417), .C2(new_n819), .ZN(new_n832));
  XNOR2_X1  g0632(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G132), .B2(new_n750), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n746), .A2(G68), .B1(G58), .B2(new_n768), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n361), .B1(new_n832), .B2(new_n833), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n736), .A2(new_n201), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n827), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n773), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n773), .A2(new_n774), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n215), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n817), .A2(new_n788), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT103), .Z(new_n845));
  AND2_X1   g0645(.A1(new_n816), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  INV_X1    g0647(.A(KEYINPUT40), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n363), .A2(new_n335), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n356), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n366), .A2(new_n850), .A3(new_n278), .A4(new_n367), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n667), .B1(new_n851), .B2(new_n390), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n403), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n400), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n854), .A2(new_n667), .B1(new_n390), .B2(new_n851), .ZN(new_n855));
  INV_X1    g0655(.A(new_n391), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n667), .B(KEYINPUT105), .Z(new_n858));
  NAND2_X1  g0658(.A1(new_n397), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n436), .A2(new_n859), .A3(new_n860), .A4(new_n391), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n853), .A2(KEYINPUT38), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT107), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n403), .A2(new_n852), .B1(new_n857), .B2(new_n861), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT107), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n436), .A2(new_n859), .A3(new_n391), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT106), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n860), .B1(new_n859), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n870), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n859), .B1(new_n435), .B2(new_n440), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n848), .B1(new_n868), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n704), .A2(new_n725), .A3(new_n877), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n331), .A2(new_n294), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n670), .A2(new_n294), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n298), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n650), .A2(new_n669), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(new_n883), .A3(new_n805), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n853), .A2(new_n862), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n869), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n863), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n876), .A2(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n443), .A3(new_n878), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n866), .B1(new_n865), .B2(KEYINPUT38), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n875), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n885), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n865), .B(new_n869), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n890), .B1(new_n897), .B2(new_n884), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(G330), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n404), .A2(new_n442), .A3(new_n434), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(G330), .A3(new_n333), .A4(new_n878), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n879), .A2(new_n669), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n875), .B(new_n906), .C1(new_n893), .C2(new_n894), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n440), .A2(new_n858), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n324), .A2(new_n669), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n808), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n883), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n910), .B1(new_n913), .B2(new_n897), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n903), .B(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n443), .A2(new_n699), .A3(new_n703), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n659), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n263), .B2(new_n785), .ZN(new_n920));
  INV_X1    g0720(.A(new_n606), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT35), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n230), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(G116), .C1(new_n922), .C2(new_n921), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT36), .ZN(new_n925));
  OAI21_X1  g0725(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n926), .A2(new_n231), .B1(G50), .B2(new_n203), .ZN(new_n927));
  INV_X1    g0727(.A(G13), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(G1), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n920), .A2(new_n925), .A3(new_n929), .ZN(G367));
  NAND2_X1  g0730(.A1(new_n686), .A2(new_n641), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT110), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n622), .B1(new_n615), .B2(new_n687), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n688), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT45), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n688), .A2(new_n934), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(new_n682), .Z(new_n940));
  XNOR2_X1  g0740(.A(new_n681), .B(new_n683), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n793), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n728), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n728), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n691), .B(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n787), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n934), .A2(new_n684), .ZN(new_n948));
  XOR2_X1   g0748(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n516), .B1(new_n932), .B2(new_n933), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n687), .B1(new_n951), .B2(new_n641), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n670), .A2(new_n560), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n639), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n628), .A2(new_n630), .A3(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g0758(.A(new_n957), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n953), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n961), .B2(new_n953), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n677), .A2(new_n681), .A3(new_n934), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n947), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n777), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n241), .B2(new_n779), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n225), .B2(new_n306), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT112), .Z(new_n970));
  AOI22_X1  g0770(.A1(new_n738), .A2(G294), .B1(G107), .B2(new_n768), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n750), .A2(G317), .ZN(new_n973));
  XNOR2_X1  g0773(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n467), .B2(new_n736), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n745), .A2(new_n244), .ZN(new_n977));
  INV_X1    g0777(.A(new_n756), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n733), .A2(new_n818), .B1(new_n978), .B2(new_n455), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n361), .B1(new_n821), .B2(new_n734), .ZN(new_n980));
  NOR4_X1   g0780(.A1(new_n976), .A2(new_n977), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n765), .A2(G58), .B1(new_n750), .B2(G137), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT114), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n759), .A2(G143), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n768), .A2(G68), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n984), .A2(new_n256), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n746), .A2(G77), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n983), .B2(new_n982), .C1(new_n201), .C2(new_n733), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(G159), .C2(new_n738), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n756), .A2(G150), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT47), .Z(new_n993));
  AOI211_X1 g0793(.A(new_n795), .B(new_n970), .C1(new_n993), .C2(new_n773), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n959), .A2(new_n776), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n966), .A2(new_n996), .ZN(G387));
  NAND2_X1  g0797(.A1(new_n942), .A2(new_n787), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n779), .B1(new_n237), .B2(new_n780), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n225), .A2(new_n256), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n693), .B2(new_n1000), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n301), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT50), .B1(new_n301), .B2(G50), .ZN(new_n1003));
  AOI21_X1  g0803(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n693), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n690), .A2(new_n220), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n967), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n977), .B1(G50), .B2(new_n756), .ZN(new_n1009));
  INV_X1    g0809(.A(G159), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n1010), .B2(new_n821), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT115), .B(G150), .Z(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(new_n750), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n361), .B1(G77), .B2(new_n765), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n732), .A2(G68), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n738), .A2(new_n302), .B1(new_n305), .B2(new_n768), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G303), .A2(new_n732), .B1(new_n738), .B2(G311), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n756), .A2(G317), .ZN(new_n1019));
  XOR2_X1   g0819(.A(KEYINPUT116), .B(G322), .Z(new_n1020));
  NAND2_X1  g0820(.A1(new_n759), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n818), .B2(new_n752), .C1(new_n753), .C2(new_n736), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT49), .Z(new_n1025));
  NAND2_X1  g0825(.A1(new_n746), .A2(new_n463), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n750), .A2(G326), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n361), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1017), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1008), .B1(new_n1029), .B2(new_n773), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1030), .B(new_n788), .C1(new_n681), .C2(new_n791), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n943), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n691), .B1(new_n942), .B2(new_n728), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n998), .B(new_n1031), .C1(new_n1032), .C2(new_n1033), .ZN(G393));
  AOI21_X1  g0834(.A(new_n692), .B1(new_n940), .B2(new_n943), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n944), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n932), .A2(new_n776), .A3(new_n933), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n746), .A2(G87), .B1(G143), .B2(new_n750), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n215), .B2(new_n752), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G150), .A2(new_n759), .B1(new_n756), .B2(G159), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n819), .A2(new_n201), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n359), .B1(new_n203), .B2(new_n736), .C1(new_n733), .C2(new_n301), .ZN(new_n1043));
  NOR4_X1   g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n732), .A2(G294), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n750), .A2(new_n1020), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n761), .A2(new_n338), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G311), .A2(new_n756), .B1(new_n759), .B2(G317), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT52), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n467), .A2(new_n752), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n819), .A2(new_n455), .B1(new_n818), .B2(new_n736), .ZN(new_n1051));
  NOR4_X1   g0851(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n773), .B1(new_n1044), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n779), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n777), .B1(new_n244), .B2(new_n225), .C1(new_n247), .C2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1037), .A2(new_n788), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n787), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n940), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1036), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(G390));
  NAND3_X1  g0860(.A1(new_n907), .A2(new_n908), .A3(new_n774), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n338), .B1(new_n756), .B2(G132), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n1010), .B2(new_n752), .C1(new_n745), .C2(new_n201), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n750), .A2(G125), .ZN(new_n1064));
  INV_X1    g0864(.A(G128), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n821), .B2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT54), .B(G143), .Z(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(new_n732), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n765), .A2(new_n1012), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1068), .B1(KEYINPUT53), .B2(new_n1069), .C1(new_n831), .C2(new_n819), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1063), .B(new_n1070), .C1(KEYINPUT53), .C2(new_n1069), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G107), .A2(new_n738), .B1(new_n756), .B2(G116), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n759), .A2(G283), .B1(new_n765), .B2(G87), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n753), .C2(new_n749), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n338), .B1(new_n215), .B2(new_n752), .C1(new_n745), .C2(new_n203), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(G97), .C2(new_n732), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n773), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n842), .A2(new_n301), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n788), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT118), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1061), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n913), .A2(new_n905), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n907), .A3(new_n908), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n727), .A2(new_n883), .A3(G330), .A4(new_n805), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n670), .B(new_n805), .C1(new_n702), .C2(new_n640), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n911), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n883), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n895), .A2(new_n1091), .A3(new_n905), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1086), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1086), .A2(new_n1092), .B1(G330), .B2(new_n885), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(new_n1057), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n917), .A2(new_n901), .A3(new_n659), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT117), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n917), .A2(new_n901), .A3(new_n659), .A4(KEYINPUT117), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n883), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n811), .B2(new_n806), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n878), .A2(new_n883), .A3(G330), .A4(new_n805), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1102), .A2(new_n1103), .B1(new_n808), .B2(new_n911), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n878), .A2(G330), .A3(new_n805), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1101), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1089), .A2(new_n911), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1106), .A2(new_n1107), .A3(new_n1087), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1099), .B(new_n1100), .C1(new_n1104), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1103), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1086), .A2(new_n1092), .A3(new_n1088), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(new_n692), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1095), .A2(new_n1109), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1084), .B(new_n1096), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(G378));
  NAND2_X1  g0917(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT120), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n915), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n421), .A2(new_n665), .A3(new_n666), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n434), .B(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n891), .B2(G330), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n899), .A2(new_n1124), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n891), .A2(G330), .A3(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n899), .A2(new_n1124), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n1130), .A3(new_n915), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT120), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1118), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1133), .B(new_n1134), .C1(new_n1095), .C2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1119), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT57), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT121), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1119), .A2(new_n1132), .A3(new_n1136), .A4(KEYINPUT57), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1141), .A2(new_n691), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT121), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1137), .A2(new_n1143), .A3(new_n1138), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1124), .A2(new_n774), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n733), .A2(new_n306), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n746), .A2(G58), .B1(G97), .B2(new_n738), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n986), .C1(new_n818), .C2(new_n749), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1147), .B(new_n1149), .C1(G116), .C2(new_n759), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n361), .B(new_n260), .C1(new_n215), .C2(new_n736), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(new_n220), .C2(new_n978), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT58), .Z(new_n1154));
  NAND2_X1  g0954(.A1(new_n765), .A2(new_n1067), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n417), .B2(new_n752), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G137), .B2(new_n732), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G132), .A2(new_n738), .B1(new_n759), .B2(G125), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n1065), .C2(new_n978), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT59), .Z(new_n1160));
  NAND2_X1  g0960(.A1(new_n254), .A2(new_n260), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT119), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n745), .A2(new_n1010), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(G124), .C2(new_n750), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1162), .B(new_n201), .C1(new_n359), .C2(G41), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n773), .B1(new_n1154), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n842), .A2(new_n201), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1146), .A2(new_n788), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1132), .B2(new_n787), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1145), .A2(new_n1172), .ZN(G375));
  NAND2_X1  g0973(.A1(new_n1135), .A2(new_n1118), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1109), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n946), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT122), .Z(new_n1178));
  NOR2_X1   g0978(.A1(new_n1135), .A2(new_n1057), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n736), .A2(new_n244), .B1(new_n455), .B2(new_n749), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT123), .Z(new_n1181));
  OAI221_X1 g0981(.A(new_n988), .B1(new_n220), .B2(new_n733), .C1(new_n753), .C2(new_n821), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G283), .C2(new_n756), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n256), .B1(new_n768), .B2(new_n305), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n467), .C2(new_n819), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT124), .Z(new_n1186));
  NOR2_X1   g0986(.A1(new_n733), .A2(new_n417), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n746), .A2(G58), .B1(G137), .B2(new_n756), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n201), .B2(new_n752), .C1(new_n1065), .C2(new_n749), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n738), .C2(new_n1067), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n759), .A2(G132), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n359), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G159), .B2(new_n765), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n773), .B1(new_n1186), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n795), .B1(new_n1101), .B2(new_n774), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n842), .A2(new_n203), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1179), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1178), .A2(new_n1198), .ZN(G381));
  NOR2_X1   g0999(.A1(G375), .A2(G378), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n947), .A2(new_n965), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n996), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1201), .A2(G390), .A3(new_n1202), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1200), .A2(new_n1203), .A3(new_n846), .A4(new_n1204), .ZN(G407));
  NAND2_X1  g1005(.A1(new_n1200), .A2(new_n668), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(G407), .A2(G213), .A3(new_n1206), .ZN(G409));
  INV_X1    g1007(.A(KEYINPUT126), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT60), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1174), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n691), .A3(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1212), .A2(G384), .A3(new_n1198), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G384), .B1(new_n1212), .B2(new_n1198), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n668), .A2(G213), .A3(G2897), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1216), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1137), .A2(new_n1143), .A3(new_n1138), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1143), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1141), .A2(new_n691), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1172), .ZN(new_n1225));
  OAI21_X1  g1025(.A(G378), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1116), .B(new_n1172), .C1(new_n1176), .C2(new_n1137), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n668), .A2(G213), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1220), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1208), .B1(new_n1231), .B2(KEYINPUT61), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1116), .B1(new_n1145), .B2(new_n1172), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(new_n1229), .ZN(new_n1235));
  OAI211_X1 g1035(.A(KEYINPUT126), .B(new_n1233), .C1(new_n1235), .C2(new_n1220), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1226), .A2(new_n1230), .A3(new_n1215), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT62), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT62), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n1239), .A3(new_n1215), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1232), .A2(new_n1236), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(G390), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(G396), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1243), .A2(new_n1203), .B1(KEYINPUT125), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n966), .A2(new_n996), .A3(new_n1059), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1244), .B(KEYINPUT125), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1242), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1241), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1237), .B1(new_n1231), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1235), .A2(KEYINPUT63), .A3(new_n1215), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1249), .A2(new_n1253), .A3(new_n1233), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(G405));
  INV_X1    g1056(.A(KEYINPUT127), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1245), .A2(new_n1257), .A3(new_n1248), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1246), .A2(new_n1242), .A3(new_n1247), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1244), .A2(KEYINPUT125), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1246), .B2(new_n1242), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT127), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1200), .A2(new_n1234), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1215), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1263), .A2(new_n1215), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1258), .B(new_n1262), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1266), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(new_n1249), .A3(KEYINPUT127), .A4(new_n1264), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(G402));
endmodule


