//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G58), .A3(G68), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G250), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n207), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n214), .B(new_n215), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n221), .A2(new_n222), .B1(new_n223), .B2(new_n207), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G50), .ZN(new_n226));
  INV_X1    g0026(.A(G226), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  OAI22_X1  g0028(.A1(new_n226), .A2(new_n227), .B1(new_n203), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(G116), .B2(G270), .ZN(new_n230));
  AND2_X1   g0030(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G68), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(G238), .ZN(new_n233));
  INV_X1    g0033(.A(G97), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n231), .B1(new_n232), .B2(new_n233), .C1(new_n234), .C2(new_n211), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(new_n208), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n220), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G238), .B(G244), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G150), .ZN(new_n256));
  INV_X1    g0056(.A(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n256), .B1(new_n258), .B2(new_n259), .C1(new_n202), .C2(new_n257), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n264), .A2(new_n257), .A3(G1), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n260), .A2(new_n263), .B1(new_n226), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n263), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G1), .B2(new_n257), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n226), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(G190), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n277), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n216), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT70), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n216), .A2(new_n284), .A3(new_n281), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n280), .B(new_n286), .C1(G77), .C2(new_n276), .ZN(new_n287));
  INV_X1    g0087(.A(G1), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT68), .B(G45), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(G274), .C1(new_n289), .C2(G41), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n281), .A2(KEYINPUT69), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT69), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G33), .A3(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n293), .A3(new_n216), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n288), .B1(G41), .B2(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n287), .B(new_n290), .C1(new_n227), .C2(new_n296), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n269), .A2(new_n270), .B1(new_n271), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n270), .B2(new_n269), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(G200), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n303), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n255), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n259), .A2(new_n306), .B1(new_n257), .B2(new_n203), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT71), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT15), .B(G87), .Z(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n258), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n311), .A2(new_n263), .B1(new_n203), .B2(new_n265), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n268), .A2(new_n203), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n277), .A2(G232), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n276), .B(new_n316), .C1(new_n277), .C2(new_n233), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n286), .C1(G107), .C2(new_n276), .ZN(new_n318));
  INV_X1    g0118(.A(new_n296), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G244), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n320), .A3(new_n290), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n321), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n315), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n297), .A2(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n297), .A2(new_n322), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n269), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n315), .A2(KEYINPUT72), .B1(new_n271), .B2(new_n321), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n305), .A2(new_n327), .A3(new_n330), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT73), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n222), .A2(G1698), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n276), .B(new_n339), .C1(G226), .C2(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n286), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n319), .A2(G238), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n290), .A4(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n283), .A2(new_n285), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n341), .B2(new_n340), .ZN(new_n348));
  INV_X1    g0148(.A(G238), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n290), .B1(new_n296), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT13), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT76), .B1(new_n352), .B2(new_n325), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n346), .A2(new_n351), .A3(new_n354), .A4(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(KEYINPUT75), .ZN(new_n358));
  INV_X1    g0158(.A(new_n352), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n322), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n352), .B(G169), .C1(KEYINPUT75), .C2(new_n357), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n265), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT74), .B1(new_n363), .B2(G68), .ZN(new_n364));
  XOR2_X1   g0164(.A(new_n364), .B(KEYINPUT12), .Z(new_n365));
  OR2_X1    g0165(.A1(new_n268), .A2(new_n232), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n306), .A2(new_n226), .B1(new_n258), .B2(new_n203), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n257), .A2(G68), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n263), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT11), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n359), .A2(new_n333), .ZN(new_n373));
  INV_X1    g0173(.A(new_n371), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n271), .B2(new_n352), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g0178(.A(new_n378), .B(KEYINPUT77), .Z(new_n379));
  NOR2_X1   g0179(.A1(new_n221), .A2(new_n232), .ZN(new_n380));
  NOR2_X1   g0180(.A1(G58), .A2(G68), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G159), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n306), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n384), .B(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n387));
  NOR2_X1   g0187(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n388));
  OAI21_X1  g0188(.A(G33), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n389), .A2(new_n273), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n273), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n257), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n391), .A2(G68), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n386), .A2(new_n395), .A3(KEYINPUT16), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT80), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(new_n393), .C1(new_n276), .C2(G20), .ZN(new_n398));
  AOI21_X1  g0198(.A(G20), .B1(new_n273), .B2(new_n275), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT80), .B1(new_n399), .B2(KEYINPUT7), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n402));
  NAND2_X1  g0202(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n272), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(G20), .B1(new_n404), .B2(new_n275), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT7), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n384), .B1(new_n407), .B2(G68), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n396), .B(new_n263), .C1(new_n408), .C2(KEYINPUT16), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n227), .A2(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n279), .A2(new_n277), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n389), .A2(new_n273), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n272), .B2(new_n223), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n286), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n319), .A2(G232), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n290), .A3(new_n415), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n416), .A2(new_n271), .ZN(new_n417));
  INV_X1    g0217(.A(new_n259), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n265), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n418), .B2(new_n268), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT81), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n416), .A2(G200), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n409), .A2(new_n417), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n409), .A2(new_n421), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n416), .A2(G169), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n416), .A2(new_n325), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n425), .A2(new_n428), .A3(KEYINPUT18), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n379), .A2(new_n424), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n338), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n228), .A2(G1698), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n349), .A2(new_n277), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n389), .A2(new_n273), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G116), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n272), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n286), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G274), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n294), .B(G250), .C1(G1), .C2(new_n442), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n392), .A2(G20), .A3(new_n232), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n223), .A2(new_n234), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n341), .A2(new_n257), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT19), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n258), .A2(new_n234), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(KEYINPUT19), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n263), .B1(new_n448), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n310), .A2(new_n265), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n263), .B(new_n265), .C1(new_n288), .C2(G33), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n309), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n325), .A2(new_n447), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n446), .A2(new_n322), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n363), .B(new_n267), .C1(G1), .C2(new_n272), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n455), .B(new_n456), .C1(new_n223), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(G200), .B2(new_n446), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n447), .A2(G190), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n255), .A2(G77), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n449), .A2(KEYINPUT6), .A3(G97), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n234), .A2(new_n449), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G97), .A2(G107), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n473), .B2(KEYINPUT6), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G20), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n398), .A2(new_n400), .B1(new_n405), .B2(KEYINPUT7), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n469), .B(new_n475), .C1(new_n476), .C2(new_n449), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n477), .A2(new_n263), .B1(new_n234), .B2(new_n265), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n458), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n228), .A2(G1698), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT4), .B1(new_n390), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n481), .A2(KEYINPUT4), .B1(G250), .B2(G1698), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n273), .A2(new_n275), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n286), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n443), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G274), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n294), .A2(new_n490), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G257), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n322), .ZN(new_n496));
  INV_X1    g0296(.A(new_n495), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n325), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n480), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(G190), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n495), .A2(G200), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n500), .A2(new_n478), .A3(new_n479), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n468), .B1(new_n503), .B2(KEYINPUT82), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n294), .A2(new_n490), .A3(G270), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n212), .A2(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n211), .A2(new_n277), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n389), .A2(new_n273), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n485), .A2(G303), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n506), .B1(new_n511), .B2(new_n286), .ZN(new_n512));
  AOI211_X1 g0312(.A(new_n505), .B(new_n322), .C1(new_n512), .C2(new_n492), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n483), .B(new_n257), .C1(G33), .C2(new_n234), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n439), .A2(G20), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n263), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT20), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n514), .A2(KEYINPUT20), .A3(new_n263), .A4(new_n515), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT83), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n261), .A2(new_n262), .B1(G20), .B2(new_n439), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n524), .A2(KEYINPUT83), .A3(new_n514), .A4(KEYINPUT20), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n516), .A2(KEYINPUT84), .A3(new_n517), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n520), .A2(new_n523), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n264), .A2(G1), .ZN(new_n528));
  INV_X1    g0328(.A(new_n515), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n458), .A2(G116), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT85), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n527), .B2(new_n530), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n513), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT86), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n513), .B(KEYINPUT86), .C1(new_n532), .C2(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n512), .A2(new_n492), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n523), .A2(new_n525), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT84), .B1(new_n516), .B2(new_n517), .ZN(new_n540));
  AOI211_X1 g0340(.A(new_n519), .B(KEYINPUT20), .C1(new_n524), .C2(new_n514), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n529), .A2(new_n528), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n463), .B2(new_n439), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT85), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n536), .A2(new_n537), .B1(G179), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n538), .A2(G169), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n545), .B2(new_n546), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n549), .B1(new_n551), .B2(KEYINPUT21), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n322), .B1(new_n512), .B2(new_n492), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n532), .B2(new_n533), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(KEYINPUT87), .A3(new_n505), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n532), .A2(new_n533), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n538), .A2(G200), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n271), .C2(new_n538), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n548), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n493), .A2(G264), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n211), .A2(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n207), .A2(new_n277), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n390), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G294), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n562), .B1(new_n567), .B2(new_n286), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n492), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT89), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n347), .B1(new_n565), .B2(new_n566), .ZN(new_n572));
  INV_X1    g0372(.A(new_n492), .ZN(new_n573));
  NOR4_X1   g0373(.A1(new_n572), .A2(new_n562), .A3(new_n570), .A4(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n575), .A3(new_n271), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(new_n333), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n528), .A2(G20), .A3(new_n449), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n223), .A2(G20), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n389), .A2(new_n273), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT88), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n389), .A2(KEYINPUT88), .A3(new_n273), .A4(new_n585), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(KEYINPUT22), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n276), .A2(new_n591), .A3(new_n585), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n258), .A2(new_n439), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n449), .A2(G20), .ZN(new_n596));
  XOR2_X1   g0396(.A(new_n596), .B(KEYINPUT23), .Z(new_n597));
  AND4_X1   g0397(.A1(new_n584), .A2(new_n593), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n594), .B1(new_n590), .B2(new_n592), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n584), .B1(new_n599), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n263), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n458), .A2(G107), .B1(new_n581), .B2(new_n580), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n578), .A2(new_n583), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n583), .A3(new_n602), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT89), .B1(new_n568), .B2(new_n492), .ZN(new_n605));
  OAI21_X1  g0405(.A(G169), .B1(new_n605), .B2(new_n574), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n568), .A2(G179), .A3(new_n492), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT82), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n499), .A2(new_n502), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n603), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n435), .A2(new_n504), .A3(new_n560), .A4(new_n612), .ZN(G372));
  INV_X1    g0413(.A(new_n305), .ZN(new_n614));
  INV_X1    g0414(.A(new_n433), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n372), .B1(new_n376), .B2(new_n327), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(new_n424), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n330), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g0418(.A(new_n618), .B(KEYINPUT93), .Z(new_n619));
  INV_X1    g0419(.A(new_n435), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n499), .A2(KEYINPUT92), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT90), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n461), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n446), .A2(KEYINPUT90), .A3(new_n322), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT92), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n480), .A2(new_n628), .A3(new_n496), .A4(new_n498), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n621), .A2(new_n622), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT26), .B1(new_n468), .B2(new_n499), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n626), .A2(new_n460), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n609), .A2(new_n548), .A3(new_n556), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n635), .A2(new_n603), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT91), .ZN(new_n637));
  INV_X1    g0437(.A(new_n503), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n627), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n635), .A2(new_n638), .A3(new_n603), .A4(new_n627), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT91), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n634), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n619), .B1(new_n620), .B2(new_n642), .ZN(G369));
  NAND2_X1  g0443(.A1(new_n548), .A2(new_n556), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n264), .A2(G20), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n288), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G343), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT94), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n557), .ZN(new_n653));
  MUX2_X1   g0453(.A(new_n560), .B(new_n644), .S(new_n653), .Z(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n603), .A2(new_n609), .ZN(new_n657));
  INV_X1    g0457(.A(new_n604), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n652), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n609), .B2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n636), .A2(new_n652), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(G399));
  NOR2_X1   g0463(.A1(new_n210), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G1), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n450), .A2(G116), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n666), .A2(new_n667), .B1(new_n218), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n642), .B2(new_n651), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT95), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n635), .A2(new_n467), .A3(new_n638), .A4(new_n603), .ZN(new_n673));
  OR3_X1    g0473(.A1(new_n468), .A2(new_n499), .A3(KEYINPUT26), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n621), .A2(new_n627), .A3(new_n629), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n632), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n652), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT96), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(KEYINPUT96), .A3(new_n652), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT29), .ZN(new_n683));
  INV_X1    g0483(.A(new_n634), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n640), .A2(KEYINPUT91), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n640), .A2(KEYINPUT91), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n652), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT95), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n670), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n672), .A2(new_n683), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n612), .A2(new_n504), .A3(new_n560), .A4(new_n652), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n497), .A2(new_n512), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n607), .A2(new_n446), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n495), .A2(new_n538), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n325), .A3(new_n446), .A4(new_n569), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n693), .A2(KEYINPUT30), .A3(new_n694), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n651), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n692), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n691), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n669), .B1(new_n709), .B2(G1), .ZN(G364));
  AOI21_X1  g0510(.A(new_n666), .B1(G45), .B2(new_n645), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n656), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(G330), .B2(new_n654), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n262), .B1(G20), .B2(new_n322), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n257), .A2(G190), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G179), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n383), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT98), .B(KEYINPUT32), .Z(new_n720));
  AOI21_X1  g0520(.A(new_n257), .B1(new_n716), .B2(G190), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n719), .A2(new_n720), .B1(G97), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n720), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n485), .B1(new_n718), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n325), .A2(G200), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n715), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n723), .B(new_n725), .C1(new_n203), .C2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n715), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n729), .A2(G179), .A3(new_n333), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n449), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n257), .A2(new_n271), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n325), .A2(new_n333), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n732), .B1(G50), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n733), .A2(new_n726), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n325), .A3(G200), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT99), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI221_X1 g0543(.A(new_n737), .B1(new_n221), .B2(new_n738), .C1(new_n743), .C2(new_n223), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n734), .A2(new_n715), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n728), .B(new_n744), .C1(G68), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n730), .A2(G283), .ZN(new_n748));
  INV_X1    g0548(.A(new_n727), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n276), .B1(new_n749), .B2(G311), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n736), .A2(G326), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n722), .A2(G294), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n748), .A2(new_n750), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT33), .B(G317), .Z(new_n754));
  INV_X1    g0554(.A(G322), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n745), .B1(new_n738), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT101), .Z(new_n757));
  INV_X1    g0557(.A(G329), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n717), .B(KEYINPUT100), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n743), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n753), .B(new_n760), .C1(G303), .C2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n714), .B1(new_n747), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n711), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n210), .A2(new_n485), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n765), .A2(G355), .B1(new_n439), .B2(new_n210), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n390), .A2(new_n210), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n768), .B1(new_n218), .B2(new_n289), .C1(new_n250), .C2(new_n442), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n714), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n764), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n773), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n763), .B(new_n775), .C1(new_n654), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n713), .A2(new_n777), .ZN(G396));
  NAND2_X1  g0578(.A1(new_n315), .A2(new_n651), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT104), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n779), .B(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n327), .B1(new_n335), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n327), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n652), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n688), .B(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(new_n707), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n764), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n730), .A2(G87), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n759), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT102), .Z(new_n793));
  NOR2_X1   g0593(.A1(new_n743), .A2(new_n449), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n738), .A2(new_n795), .B1(new_n721), .B2(new_n234), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(KEYINPUT103), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(KEYINPUT103), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n485), .B1(new_n727), .B2(new_n439), .C1(new_n799), .C2(new_n745), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n794), .A2(new_n797), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n793), .B(new_n801), .C1(new_n802), .C2(new_n735), .ZN(new_n803));
  INV_X1    g0603(.A(new_n738), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G143), .A2(new_n804), .B1(new_n746), .B2(G150), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n805), .B1(new_n806), .B2(new_n735), .C1(new_n383), .C2(new_n727), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT34), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n730), .A2(G68), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n743), .A2(new_n226), .B1(new_n810), .B2(new_n759), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G58), .B2(new_n722), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n803), .B1(new_n813), .B2(new_n392), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n714), .A2(new_n771), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(new_n714), .B1(new_n203), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n711), .B(new_n816), .C1(new_n786), .C2(new_n772), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT105), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n789), .A2(new_n818), .ZN(G384));
  NAND4_X1  g0619(.A1(new_n672), .A2(new_n435), .A3(new_n683), .A4(new_n690), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n619), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n687), .A2(new_n652), .A3(new_n786), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n784), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT38), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n386), .A2(new_n395), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT16), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(new_n263), .A3(new_n396), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n421), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n428), .B2(new_n649), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n825), .B1(new_n831), .B2(new_n423), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n425), .A2(new_n649), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n429), .A2(KEYINPUT107), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT107), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n425), .A2(new_n428), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n834), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n423), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n832), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n830), .A2(new_n649), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n433), .B2(new_n424), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n824), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n433), .A2(new_n424), .ZN(new_n845));
  INV_X1    g0645(.A(new_n842), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n425), .A2(new_n428), .A3(new_n836), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n836), .B1(new_n425), .B2(new_n428), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n833), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n840), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n831), .A2(new_n423), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n850), .A2(new_n851), .B1(new_n852), .B2(new_n825), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n847), .A2(new_n853), .A3(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n651), .A2(new_n371), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n372), .A2(new_n377), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT106), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT106), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n372), .A2(new_n377), .A3(new_n859), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n362), .A2(new_n371), .A3(new_n651), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n823), .A2(new_n855), .A3(new_n863), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n844), .A2(new_n854), .A3(KEYINPUT39), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n833), .B1(new_n433), .B2(new_n424), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT108), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n426), .A2(new_n427), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n409), .B2(new_n421), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n868), .B1(new_n839), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n429), .A2(KEYINPUT108), .A3(new_n423), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n833), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n838), .A2(new_n840), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n867), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n854), .B1(new_n876), .B2(KEYINPUT38), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n865), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n372), .A2(new_n651), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n649), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n615), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n864), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n821), .B(new_n883), .Z(new_n884));
  NAND2_X1  g0684(.A1(new_n435), .A2(new_n706), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n785), .B1(new_n861), .B2(new_n862), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n855), .A2(new_n886), .A3(new_n706), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n877), .A2(KEYINPUT40), .A3(new_n706), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n885), .B(new_n891), .Z(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(G330), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n884), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n288), .B2(new_n645), .ZN(new_n895));
  OAI211_X1 g0695(.A(G20), .B(new_n216), .C1(new_n474), .C2(KEYINPUT35), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n439), .B(new_n896), .C1(KEYINPUT35), .C2(new_n474), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT36), .Z(new_n898));
  NOR2_X1   g0698(.A1(new_n201), .A2(new_n232), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n380), .A2(new_n218), .A3(new_n203), .ZN(new_n900));
  OAI211_X1 g0700(.A(G1), .B(new_n264), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(new_n898), .A3(new_n901), .ZN(G367));
  NAND2_X1  g0702(.A1(new_n480), .A2(new_n651), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n638), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT109), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n905), .A2(new_n609), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n651), .B1(new_n906), .B2(new_n499), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n499), .B2(new_n652), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n651), .B1(new_n548), .B2(new_n556), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n657), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT42), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n651), .A2(new_n464), .ZN(new_n915));
  MUX2_X1   g0715(.A(new_n627), .B(new_n632), .S(new_n915), .Z(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(KEYINPUT110), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT110), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n914), .B2(new_n917), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n914), .A2(new_n917), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n919), .A2(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n661), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n908), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT111), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n927), .A2(new_n928), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n664), .B(KEYINPUT41), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT113), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT112), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n657), .A2(new_n909), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n660), .B2(new_n909), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(new_n655), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n709), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT112), .B1(new_n708), .B2(new_n939), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n905), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n662), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT44), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n908), .A2(new_n662), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT45), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(new_n661), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n935), .B1(new_n943), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n925), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n952), .A2(new_n941), .A3(KEYINPUT113), .A4(new_n942), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n934), .B1(new_n954), .B2(new_n709), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n288), .B1(new_n645), .B2(G45), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n932), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n721), .A2(new_n232), .ZN(new_n959));
  INV_X1    g0759(.A(G150), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n731), .A2(new_n203), .B1(new_n960), .B2(new_n738), .ZN(new_n961));
  INV_X1    g0761(.A(new_n717), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n959), .B(new_n961), .C1(G137), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n761), .A2(G58), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n485), .B1(new_n736), .B2(G143), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n746), .A2(G159), .B1(new_n749), .B2(new_n201), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT115), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT116), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT46), .B1(new_n761), .B2(G116), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT114), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n972));
  INV_X1    g0772(.A(G317), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n735), .A2(new_n791), .B1(new_n717), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G294), .B2(new_n746), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n390), .B1(G303), .B2(new_n804), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n730), .A2(G97), .B1(G107), .B2(new_n722), .ZN(new_n977));
  AND4_X1   g0777(.A1(new_n972), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n971), .B(new_n978), .C1(new_n799), .C2(new_n727), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n969), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n764), .B1(new_n981), .B2(new_n714), .ZN(new_n982));
  INV_X1    g0782(.A(new_n768), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n774), .B1(new_n209), .B2(new_n310), .C1(new_n983), .C2(new_n246), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n776), .C2(new_n916), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n958), .A2(new_n985), .ZN(G387));
  OAI211_X1 g0786(.A(new_n943), .B(new_n664), .C1(new_n709), .C2(new_n940), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n983), .B1(new_n243), .B2(new_n289), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n667), .B2(new_n765), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n418), .A2(new_n226), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n667), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n991), .B(new_n442), .C1(KEYINPUT50), .C2(new_n990), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G68), .B2(G77), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n989), .A2(new_n993), .B1(G107), .B2(new_n209), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n764), .B1(new_n994), .B2(new_n774), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G311), .A2(new_n746), .B1(new_n804), .B2(G317), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n802), .B2(new_n727), .C1(new_n755), .C2(new_n735), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT48), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n799), .B2(new_n721), .C1(new_n795), .C2(new_n743), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT49), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n962), .A2(G326), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1000), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n390), .B1(G116), .B2(new_n730), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n745), .A2(new_n259), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n310), .A2(new_n721), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n390), .B1(new_n383), .B2(new_n735), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(G97), .C2(new_n730), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n738), .A2(new_n226), .B1(new_n727), .B2(new_n232), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G150), .B2(new_n962), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(new_n203), .C2(new_n743), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1005), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT117), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n714), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n995), .B1(new_n660), .B2(new_n776), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n939), .B2(new_n956), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n987), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT118), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT118), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n987), .A2(new_n1021), .A3(new_n1018), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(G393));
  NAND2_X1  g0823(.A1(new_n952), .A2(new_n957), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n774), .B1(new_n234), .B2(new_n209), .C1(new_n983), .C2(new_n253), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n201), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n790), .B1(new_n1026), .B2(new_n745), .C1(new_n259), .C2(new_n727), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n392), .B(new_n1027), .C1(G77), .C2(new_n722), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n761), .A2(G68), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n962), .A2(G143), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n735), .A2(new_n960), .B1(new_n738), .B2(new_n383), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT51), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n735), .A2(new_n973), .B1(new_n738), .B2(new_n791), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT52), .Z(new_n1035));
  AOI22_X1  g0835(.A1(G294), .A2(new_n749), .B1(new_n962), .B2(G322), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n439), .B2(new_n721), .C1(new_n802), .C2(new_n745), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n743), .A2(new_n799), .ZN(new_n1038));
  OR4_X1    g0838(.A1(new_n276), .A2(new_n1035), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1033), .B1(new_n732), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n764), .B1(new_n1040), .B2(new_n714), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1025), .B(new_n1041), .C1(new_n908), .C2(new_n776), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1024), .A2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n951), .A2(new_n953), .B1(new_n943), .B2(new_n950), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n664), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(G390));
  NAND3_X1  g0846(.A1(new_n886), .A2(G330), .A3(new_n706), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n642), .A2(new_n651), .A3(new_n785), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n784), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n863), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n879), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n878), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n877), .A2(new_n1052), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n681), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT96), .B1(new_n677), .B2(new_n652), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n782), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n784), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1054), .B1(new_n1058), .B2(new_n863), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1048), .B1(new_n1053), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n435), .A2(G330), .A3(new_n706), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n820), .A2(new_n619), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n877), .A2(new_n866), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n866), .B2(new_n855), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n863), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n822), .B2(new_n784), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1066), .B2(new_n879), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1054), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1050), .B1(new_n682), .B2(new_n782), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n1065), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1070), .A3(new_n1047), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n706), .A2(G330), .A3(new_n786), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1065), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n1047), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n823), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1057), .A2(new_n1073), .A3(new_n784), .A4(new_n1047), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1060), .A2(new_n1062), .A3(new_n1071), .A4(new_n1077), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1077), .A2(new_n619), .A3(new_n820), .A4(new_n1061), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1067), .A2(new_n1070), .A3(new_n1047), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1047), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1078), .A2(new_n1082), .A3(new_n664), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1060), .A2(new_n957), .A3(new_n1071), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT119), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT119), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1060), .A2(new_n1086), .A3(new_n957), .A4(new_n1071), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1064), .A2(new_n771), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G107), .A2(new_n746), .B1(new_n749), .B2(G97), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n439), .B2(new_n738), .C1(new_n799), .C2(new_n735), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G77), .B2(new_n722), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n759), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n761), .A2(G87), .B1(new_n1093), .B2(G294), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1092), .A2(new_n485), .A3(new_n809), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n276), .B1(new_n383), .B2(new_n721), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n736), .A2(G128), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1097), .B1(new_n806), .B2(new_n745), .C1(new_n727), .C2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1096), .B(new_n1099), .C1(new_n201), .C2(new_n730), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n743), .A2(new_n960), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1100), .B(new_n1102), .C1(new_n1103), .C2(new_n759), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n738), .A2(new_n810), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1095), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1106), .A2(new_n714), .B1(new_n259), .B2(new_n815), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1089), .A2(new_n711), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT120), .B1(new_n1088), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT120), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1111), .B(new_n1108), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1083), .B1(new_n1110), .B2(new_n1112), .ZN(G378));
  NAND3_X1  g0913(.A1(new_n889), .A2(new_n890), .A3(G330), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT124), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT55), .Z(new_n1118));
  INV_X1    g0918(.A(new_n330), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n302), .B2(new_n304), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT123), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n269), .A2(new_n649), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n305), .A2(new_n330), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT123), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1118), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1124), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1126), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1116), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT124), .A4(G330), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1066), .A2(new_n855), .B1(new_n878), .B2(new_n879), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n882), .ZN(new_n1137));
  AND4_X1   g0937(.A1(new_n882), .A2(new_n864), .A3(new_n1135), .A4(new_n880), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1135), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n883), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n882), .A3(new_n1135), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1115), .B2(new_n1114), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1139), .A2(new_n957), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n771), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n815), .A2(new_n1026), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G128), .A2(new_n804), .B1(new_n746), .B2(G132), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1103), .B2(new_n735), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G150), .B2(new_n722), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n806), .B2(new_n727), .C1(new_n743), .C2(new_n1098), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT59), .Z(new_n1153));
  AOI21_X1  g0953(.A(G41), .B1(new_n962), .B2(G124), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G33), .B1(new_n730), .B2(G159), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n387), .A2(new_n388), .A3(new_n272), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n226), .B1(new_n1157), .B2(G41), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n746), .A2(G97), .B1(new_n749), .B2(new_n309), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n449), .B2(new_n738), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G41), .B(new_n1160), .C1(G58), .C2(new_n730), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n959), .B1(G116), .B2(new_n736), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT121), .Z(new_n1163));
  AOI22_X1  g0963(.A1(new_n761), .A2(G77), .B1(new_n1093), .B2(G283), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n392), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT58), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1156), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n764), .B1(new_n1167), .B2(new_n714), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1147), .A2(new_n1148), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1146), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1144), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1078), .A2(new_n1062), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1175), .A3(KEYINPUT57), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n664), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1171), .B1(new_n1177), .B2(new_n1178), .ZN(G375));
  NAND3_X1  g0979(.A1(new_n820), .A2(new_n619), .A3(new_n1061), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n933), .A3(new_n1079), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1065), .A2(new_n771), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G294), .A2(new_n736), .B1(new_n749), .B2(G107), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n439), .B2(new_n745), .C1(new_n799), .C2(new_n738), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1186), .A2(new_n276), .A3(new_n1007), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n761), .A2(G97), .B1(new_n1093), .B2(G303), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n203), .C2(new_n731), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n735), .A2(new_n810), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n806), .A2(new_n738), .B1(new_n745), .B2(new_n1098), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n761), .B2(G159), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n392), .B1(G150), .B2(new_n749), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n730), .A2(G58), .B1(G50), .B2(new_n722), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1093), .A2(G128), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1189), .B1(new_n1190), .B2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1197), .A2(new_n714), .B1(new_n232), .B2(new_n815), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1184), .A2(new_n711), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1077), .B2(new_n957), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1183), .A2(new_n1200), .ZN(G381));
  AND3_X1   g1001(.A1(new_n958), .A2(new_n985), .A3(new_n1045), .ZN(new_n1202));
  INV_X1    g1002(.A(G384), .ZN(new_n1203));
  INV_X1    g1003(.A(G381), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G393), .A2(G396), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1180), .B1(new_n1207), .B2(new_n1077), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n665), .B1(new_n1210), .B2(KEYINPUT57), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1178), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1170), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1110), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1088), .A2(KEYINPUT120), .A3(new_n1109), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1083), .A3(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1206), .A2(new_n1217), .ZN(G407));
  AND2_X1   g1018(.A1(new_n1206), .A2(G343), .ZN(new_n1219));
  OAI21_X1  g1019(.A(G213), .B1(new_n1219), .B2(new_n1217), .ZN(G409));
  NAND2_X1  g1020(.A1(G375), .A2(G378), .ZN(new_n1221));
  INV_X1    g1021(.A(G213), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(G343), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1170), .B1(new_n1210), .B2(new_n933), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n1083), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1221), .A2(new_n1224), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n664), .B(new_n1079), .C1(new_n1182), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT60), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1200), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1203), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G384), .B(new_n1200), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT125), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1223), .A2(G2897), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1232), .A2(KEYINPUT125), .A3(new_n1233), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1227), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1221), .A2(new_n1242), .A3(new_n1224), .A4(new_n1226), .ZN(new_n1243));
  XOR2_X1   g1043(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1223), .B1(G375), .B2(G378), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1242), .A3(new_n1226), .A4(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1241), .A2(new_n1245), .A3(new_n1246), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT127), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1238), .B1(new_n1247), .B2(new_n1226), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT61), .B1(new_n1252), .B2(new_n1240), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT127), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1245), .A4(new_n1249), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1045), .B1(new_n958), .B2(new_n985), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1020), .A2(new_n1022), .B1(new_n777), .B2(new_n713), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1202), .A2(new_n1256), .B1(new_n1205), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(G390), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n958), .A2(new_n985), .A3(new_n1045), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1205), .A2(new_n1257), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1258), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1251), .A2(new_n1255), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT61), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1243), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT63), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1241), .A2(KEYINPUT63), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1265), .B(new_n1267), .C1(new_n1266), .C2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1264), .A2(new_n1269), .ZN(G405));
  NAND2_X1  g1070(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(new_n1242), .Z(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(new_n1263), .ZN(G402));
endmodule


