

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767;

  AND2_X1 U369 ( .A1(n349), .A2(n348), .ZN(n640) );
  INV_X1 U370 ( .A(n738), .ZN(n348) );
  AND2_X1 U371 ( .A1(n384), .A2(n421), .ZN(n382) );
  NOR2_X1 U372 ( .A1(n766), .A2(n765), .ZN(n565) );
  NOR2_X1 U373 ( .A1(n706), .A2(n711), .ZN(n387) );
  NOR2_X1 U374 ( .A1(n538), .A2(n537), .ZN(n559) );
  BUF_X1 U375 ( .A(n536), .Z(n699) );
  AND2_X1 U376 ( .A1(n595), .A2(n539), .ZN(n547) );
  XNOR2_X1 U377 ( .A(n481), .B(n431), .ZN(n751) );
  XNOR2_X1 U378 ( .A(G902), .B(KEYINPUT15), .ZN(n616) );
  XNOR2_X1 U379 ( .A(n507), .B(n508), .ZN(n509) );
  INV_X1 U380 ( .A(G146), .ZN(n449) );
  XNOR2_X1 U381 ( .A(G113), .B(KEYINPUT3), .ZN(n378) );
  INV_X1 U382 ( .A(G953), .ZN(n755) );
  XNOR2_X1 U383 ( .A(n638), .B(n350), .ZN(n349) );
  INV_X1 U384 ( .A(n637), .ZN(n350) );
  XNOR2_X2 U385 ( .A(n606), .B(KEYINPUT92), .ZN(n608) );
  AND2_X2 U386 ( .A1(n411), .A2(n410), .ZN(n376) );
  NOR2_X2 U387 ( .A1(n554), .A2(n553), .ZN(n567) );
  NOR2_X2 U388 ( .A1(n558), .A2(n550), .ZN(n675) );
  XNOR2_X2 U389 ( .A(n414), .B(n519), .ZN(n541) );
  NOR2_X1 U390 ( .A1(G953), .A2(G237), .ZN(n471) );
  XOR2_X1 U391 ( .A(n524), .B(n403), .Z(n351) );
  XNOR2_X2 U392 ( .A(n398), .B(n361), .ZN(n644) );
  XNOR2_X2 U393 ( .A(n588), .B(n587), .ZN(n393) );
  XNOR2_X1 U394 ( .A(n404), .B(n470), .ZN(n653) );
  NAND2_X1 U395 ( .A1(n385), .A2(n383), .ZN(n381) );
  AND2_X1 U396 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U397 ( .A1(n397), .A2(n355), .ZN(n588) );
  XNOR2_X1 U398 ( .A(n387), .B(KEYINPUT41), .ZN(n705) );
  NAND2_X1 U399 ( .A1(n408), .A2(n409), .ZN(n375) );
  XNOR2_X1 U400 ( .A(n609), .B(KEYINPUT1), .ZN(n601) );
  XNOR2_X1 U401 ( .A(n479), .B(n478), .ZN(n557) );
  XNOR2_X1 U402 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U403 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U404 ( .A(n510), .B(n464), .ZN(n481) );
  XNOR2_X1 U405 ( .A(n512), .B(G134), .ZN(n459) );
  XNOR2_X1 U406 ( .A(KEYINPUT4), .B(G101), .ZN(n529) );
  XNOR2_X1 U407 ( .A(G104), .B(G122), .ZN(n504) );
  NAND2_X1 U408 ( .A1(n726), .A2(n365), .ZN(n352) );
  AND2_X1 U409 ( .A1(n380), .A2(n353), .ZN(n368) );
  AND2_X1 U410 ( .A1(n767), .A2(KEYINPUT2), .ZN(n353) );
  NAND2_X1 U411 ( .A1(n726), .A2(n365), .ZN(n628) );
  XNOR2_X2 U412 ( .A(n549), .B(KEYINPUT19), .ZN(n583) );
  XNOR2_X2 U413 ( .A(n399), .B(n584), .ZN(n606) );
  NOR2_X2 U414 ( .A1(n583), .A2(n582), .ZN(n399) );
  XNOR2_X2 U415 ( .A(n628), .B(n627), .ZN(n363) );
  XNOR2_X2 U416 ( .A(n352), .B(n627), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n449), .B(G125), .ZN(n510) );
  INV_X1 U418 ( .A(KEYINPUT10), .ZN(n464) );
  NAND2_X1 U419 ( .A1(n678), .A2(n547), .ZN(n501) );
  NOR2_X1 U420 ( .A1(n521), .A2(KEYINPUT87), .ZN(n409) );
  XNOR2_X1 U421 ( .A(n752), .B(n449), .ZN(n531) );
  XNOR2_X1 U422 ( .A(n427), .B(KEYINPUT112), .ZN(n558) );
  XNOR2_X1 U423 ( .A(n430), .B(n429), .ZN(n428) );
  NAND2_X1 U424 ( .A1(n374), .A2(n354), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n448), .B(G131), .ZN(n465) );
  INV_X1 U426 ( .A(KEYINPUT66), .ZN(n448) );
  XNOR2_X1 U427 ( .A(n459), .B(n465), .ZN(n752) );
  NAND2_X1 U428 ( .A1(n601), .A2(n610), .ZN(n440) );
  INV_X1 U429 ( .A(n527), .ZN(n431) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n467) );
  XNOR2_X1 U431 ( .A(G140), .B(KEYINPUT98), .ZN(n466) );
  INV_X1 U432 ( .A(n481), .ZN(n405) );
  XNOR2_X1 U433 ( .A(G143), .B(G113), .ZN(n474) );
  XNOR2_X1 U434 ( .A(G104), .B(G107), .ZN(n526) );
  INV_X1 U435 ( .A(n560), .ZN(n400) );
  XNOR2_X1 U436 ( .A(n691), .B(KEYINPUT88), .ZN(n589) );
  INV_X1 U437 ( .A(KEYINPUT36), .ZN(n403) );
  XNOR2_X1 U438 ( .A(n699), .B(KEYINPUT6), .ZN(n596) );
  XNOR2_X1 U439 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U440 ( .A(G475), .ZN(n476) );
  OR2_X1 U441 ( .A1(n631), .A2(G902), .ZN(n535) );
  NAND2_X1 U442 ( .A1(n351), .A2(n419), .ZN(n423) );
  INV_X1 U443 ( .A(n589), .ZN(n419) );
  INV_X1 U444 ( .A(G237), .ZN(n517) );
  NAND2_X1 U445 ( .A1(n521), .A2(KEYINPUT87), .ZN(n410) );
  XNOR2_X1 U446 ( .A(G137), .B(G116), .ZN(n444) );
  XOR2_X1 U447 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n441) );
  AND2_X1 U448 ( .A1(n422), .A2(n424), .ZN(n421) );
  INV_X1 U449 ( .A(n686), .ZN(n424) );
  AND2_X1 U450 ( .A1(n423), .A2(n568), .ZN(n383) );
  XNOR2_X1 U451 ( .A(KEYINPUT90), .B(KEYINPUT17), .ZN(n508) );
  NAND2_X1 U452 ( .A1(G237), .A2(G234), .ZN(n491) );
  XNOR2_X1 U453 ( .A(n575), .B(KEYINPUT38), .ZN(n709) );
  INV_X1 U454 ( .A(n601), .ZN(n691) );
  INV_X1 U455 ( .A(KEYINPUT28), .ZN(n429) );
  XNOR2_X1 U456 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U457 ( .A(G119), .B(G128), .ZN(n482) );
  XOR2_X1 U458 ( .A(KEYINPUT24), .B(G110), .Z(n483) );
  XNOR2_X1 U459 ( .A(n455), .B(n434), .ZN(n485) );
  INV_X1 U460 ( .A(KEYINPUT8), .ZN(n434) );
  XNOR2_X1 U461 ( .A(n597), .B(KEYINPUT33), .ZN(n715) );
  NOR2_X1 U462 ( .A1(n440), .A2(n596), .ZN(n597) );
  BUF_X1 U463 ( .A(n541), .Z(n575) );
  INV_X1 U464 ( .A(KEYINPUT0), .ZN(n584) );
  INV_X1 U465 ( .A(n440), .ZN(n605) );
  XNOR2_X1 U466 ( .A(n490), .B(n489), .ZN(n595) );
  NOR2_X1 U467 ( .A1(G902), .A2(n637), .ZN(n490) );
  XNOR2_X1 U468 ( .A(n645), .B(n646), .ZN(n647) );
  XNOR2_X1 U469 ( .A(n432), .B(n751), .ZN(n637) );
  XNOR2_X1 U470 ( .A(n435), .B(n433), .ZN(n432) );
  NAND2_X1 U471 ( .A1(n485), .A2(G221), .ZN(n433) );
  XNOR2_X1 U472 ( .A(n484), .B(n356), .ZN(n435) );
  XNOR2_X1 U473 ( .A(n475), .B(n405), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n531), .B(n437), .ZN(n631) );
  XNOR2_X1 U475 ( .A(n439), .B(n438), .ZN(n437) );
  XNOR2_X1 U476 ( .A(n530), .B(n525), .ZN(n439) );
  XNOR2_X1 U477 ( .A(n661), .B(n660), .ZN(n662) );
  AND2_X1 U478 ( .A1(n634), .A2(G953), .ZN(n738) );
  XNOR2_X1 U479 ( .A(n386), .B(KEYINPUT42), .ZN(n766) );
  XNOR2_X1 U480 ( .A(n564), .B(n401), .ZN(n765) );
  INV_X1 U481 ( .A(KEYINPUT40), .ZN(n401) );
  NAND2_X1 U482 ( .A1(n393), .A2(n415), .ZN(n398) );
  AND2_X1 U483 ( .A1(n590), .A2(n596), .ZN(n415) );
  INV_X1 U484 ( .A(KEYINPUT110), .ZN(n395) );
  INV_X1 U485 ( .A(n598), .ZN(n545) );
  INV_X1 U486 ( .A(KEYINPUT105), .ZN(n402) );
  INV_X1 U487 ( .A(n423), .ZN(n683) );
  AND2_X1 U488 ( .A1(n644), .A2(n357), .ZN(n354) );
  AND2_X1 U489 ( .A1(n585), .A2(n689), .ZN(n355) );
  XNOR2_X1 U490 ( .A(KEYINPUT23), .B(KEYINPUT93), .ZN(n356) );
  AND2_X1 U491 ( .A1(n642), .A2(KEYINPUT44), .ZN(n357) );
  AND2_X1 U492 ( .A1(n667), .A2(n614), .ZN(n358) );
  AND2_X1 U493 ( .A1(n721), .A2(n620), .ZN(n359) );
  XNOR2_X1 U494 ( .A(n598), .B(KEYINPUT75), .ZN(n360) );
  XOR2_X1 U495 ( .A(KEYINPUT77), .B(KEYINPUT32), .Z(n361) );
  XNOR2_X1 U496 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n362) );
  XNOR2_X1 U497 ( .A(n531), .B(n450), .ZN(n645) );
  INV_X1 U498 ( .A(n568), .ZN(n425) );
  BUF_X1 U499 ( .A(n721), .Z(n744) );
  AND2_X1 U500 ( .A1(n371), .A2(n372), .ZN(n370) );
  INV_X2 U501 ( .A(KEYINPUT69), .ZN(n377) );
  NAND2_X1 U502 ( .A1(n366), .A2(n626), .ZN(n365) );
  NAND2_X1 U503 ( .A1(n359), .A2(n619), .ZN(n366) );
  XNOR2_X2 U504 ( .A(n367), .B(KEYINPUT72), .ZN(n726) );
  NAND2_X1 U505 ( .A1(n721), .A2(n368), .ZN(n367) );
  XNOR2_X2 U506 ( .A(n412), .B(KEYINPUT45), .ZN(n721) );
  NAND2_X1 U507 ( .A1(n370), .A2(n369), .ZN(n413) );
  NAND2_X1 U508 ( .A1(n643), .A2(n436), .ZN(n371) );
  NAND2_X1 U509 ( .A1(n373), .A2(n436), .ZN(n372) );
  NAND2_X1 U510 ( .A1(n644), .A2(n642), .ZN(n373) );
  INV_X1 U511 ( .A(n643), .ZN(n374) );
  XNOR2_X2 U512 ( .A(n599), .B(KEYINPUT35), .ZN(n643) );
  NAND2_X2 U513 ( .A1(n376), .A2(n375), .ZN(n549) );
  XNOR2_X2 U514 ( .A(n377), .B(G119), .ZN(n379) );
  XNOR2_X2 U515 ( .A(n739), .B(n529), .ZN(n506) );
  XNOR2_X2 U516 ( .A(n379), .B(n378), .ZN(n739) );
  NAND2_X2 U517 ( .A1(n380), .A2(n767), .ZN(n754) );
  AND2_X2 U518 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U519 ( .A1(n426), .A2(n425), .ZN(n384) );
  INV_X1 U520 ( .A(n426), .ZN(n385) );
  NOR2_X1 U521 ( .A1(n558), .A2(n705), .ZN(n386) );
  NAND2_X1 U522 ( .A1(n389), .A2(n388), .ZN(n392) );
  NOR2_X1 U523 ( .A1(n715), .A2(n362), .ZN(n388) );
  INV_X1 U524 ( .A(n608), .ZN(n389) );
  NAND2_X1 U525 ( .A1(n390), .A2(n406), .ZN(n599) );
  NAND2_X1 U526 ( .A1(n608), .A2(n362), .ZN(n391) );
  NAND2_X1 U527 ( .A1(n393), .A2(n596), .ZN(n600) );
  NAND2_X1 U528 ( .A1(n393), .A2(n593), .ZN(n642) );
  INV_X1 U529 ( .A(n606), .ZN(n397) );
  XNOR2_X1 U530 ( .A(n394), .B(KEYINPUT30), .ZN(n538) );
  NAND2_X1 U531 ( .A1(n536), .A2(n708), .ZN(n394) );
  XNOR2_X2 U532 ( .A(n396), .B(n395), .ZN(n764) );
  NAND2_X1 U533 ( .A1(n546), .A2(n545), .ZN(n396) );
  AND2_X1 U534 ( .A1(n407), .A2(n360), .ZN(n406) );
  XNOR2_X1 U535 ( .A(n543), .B(KEYINPUT109), .ZN(n546) );
  NAND2_X1 U536 ( .A1(n413), .A2(n358), .ZN(n412) );
  AND2_X1 U537 ( .A1(n559), .A2(n400), .ZN(n561) );
  XNOR2_X2 U538 ( .A(n563), .B(n402), .ZN(n678) );
  NAND2_X1 U539 ( .A1(n351), .A2(n420), .ZN(n422) );
  NAND2_X1 U540 ( .A1(n715), .A2(n362), .ZN(n407) );
  INV_X1 U541 ( .A(n541), .ZN(n408) );
  NAND2_X1 U542 ( .A1(n541), .A2(KEYINPUT87), .ZN(n411) );
  NAND2_X1 U543 ( .A1(n658), .A2(n616), .ZN(n414) );
  XNOR2_X1 U544 ( .A(n416), .B(KEYINPUT80), .ZN(n554) );
  NAND2_X1 U545 ( .A1(n417), .A2(n418), .ZN(n416) );
  XNOR2_X1 U546 ( .A(n764), .B(KEYINPUT81), .ZN(n417) );
  NAND2_X1 U547 ( .A1(n552), .A2(KEYINPUT47), .ZN(n418) );
  NAND2_X1 U548 ( .A1(n675), .A2(n551), .ZN(n552) );
  NOR2_X1 U549 ( .A1(n589), .A2(n568), .ZN(n420) );
  NAND2_X1 U550 ( .A1(n567), .A2(n566), .ZN(n426) );
  NAND2_X1 U551 ( .A1(n428), .A2(n548), .ZN(n427) );
  NAND2_X1 U552 ( .A1(n547), .A2(n699), .ZN(n430) );
  INV_X1 U553 ( .A(KEYINPUT44), .ZN(n436) );
  XNOR2_X1 U554 ( .A(n527), .B(n526), .ZN(n438) );
  NOR2_X1 U555 ( .A1(n595), .A2(n594), .ZN(n610) );
  NOR2_X2 U556 ( .A1(n555), .A2(n557), .ZN(n563) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n443) );
  XNOR2_X1 U558 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U559 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U560 ( .A(n488), .B(n487), .ZN(n489) );
  BUF_X1 U561 ( .A(n658), .Z(n661) );
  NAND2_X1 U562 ( .A1(n471), .A2(G210), .ZN(n442) );
  XNOR2_X1 U563 ( .A(n442), .B(n441), .ZN(n446) );
  XNOR2_X1 U564 ( .A(n506), .B(n447), .ZN(n450) );
  XNOR2_X2 U565 ( .A(G143), .B(G128), .ZN(n512) );
  INV_X1 U566 ( .A(G902), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n645), .A2(n518), .ZN(n452) );
  XOR2_X1 U568 ( .A(KEYINPUT97), .B(G472), .Z(n451) );
  XNOR2_X2 U569 ( .A(n452), .B(n451), .ZN(n536) );
  XNOR2_X1 U570 ( .A(KEYINPUT103), .B(G478), .ZN(n463) );
  XOR2_X1 U571 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n454) );
  XNOR2_X1 U572 ( .A(G122), .B(KEYINPUT7), .ZN(n453) );
  XNOR2_X1 U573 ( .A(n454), .B(n453), .ZN(n457) );
  NAND2_X1 U574 ( .A1(G234), .A2(n755), .ZN(n455) );
  NAND2_X1 U575 ( .A1(G217), .A2(n485), .ZN(n456) );
  XNOR2_X1 U576 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X2 U577 ( .A(G107), .B(G116), .ZN(n503) );
  XNOR2_X1 U578 ( .A(n503), .B(KEYINPUT101), .ZN(n458) );
  XNOR2_X1 U579 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U580 ( .A(n461), .B(n460), .ZN(n734) );
  NOR2_X1 U581 ( .A1(G902), .A2(n734), .ZN(n462) );
  XNOR2_X1 U582 ( .A(n463), .B(n462), .ZN(n555) );
  XNOR2_X1 U583 ( .A(n465), .B(KEYINPUT12), .ZN(n469) );
  XNOR2_X1 U584 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U585 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U586 ( .A1(G214), .A2(n471), .ZN(n472) );
  XNOR2_X1 U587 ( .A(n472), .B(n504), .ZN(n473) );
  XOR2_X1 U588 ( .A(n474), .B(n473), .Z(n475) );
  NOR2_X1 U589 ( .A1(G902), .A2(n653), .ZN(n479) );
  XNOR2_X1 U590 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n477) );
  INV_X1 U591 ( .A(G140), .ZN(n480) );
  XNOR2_X1 U592 ( .A(n480), .B(G137), .ZN(n527) );
  NAND2_X1 U593 ( .A1(n616), .A2(G234), .ZN(n486) );
  XNOR2_X1 U594 ( .A(n486), .B(KEYINPUT20), .ZN(n497) );
  NAND2_X1 U595 ( .A1(n497), .A2(G217), .ZN(n488) );
  XOR2_X1 U596 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n487) );
  XNOR2_X1 U597 ( .A(n491), .B(KEYINPUT14), .ZN(n493) );
  NAND2_X1 U598 ( .A1(G952), .A2(n493), .ZN(n720) );
  NOR2_X1 U599 ( .A1(n720), .A2(G953), .ZN(n492) );
  XNOR2_X1 U600 ( .A(n492), .B(KEYINPUT91), .ZN(n581) );
  NAND2_X1 U601 ( .A1(G902), .A2(n493), .ZN(n578) );
  NOR2_X1 U602 ( .A1(G900), .A2(n578), .ZN(n494) );
  NAND2_X1 U603 ( .A1(G953), .A2(n494), .ZN(n495) );
  NAND2_X1 U604 ( .A1(n581), .A2(n495), .ZN(n496) );
  XNOR2_X1 U605 ( .A(n496), .B(KEYINPUT78), .ZN(n500) );
  NAND2_X1 U606 ( .A1(G221), .A2(n497), .ZN(n499) );
  INV_X1 U607 ( .A(KEYINPUT21), .ZN(n498) );
  XNOR2_X1 U608 ( .A(n499), .B(n498), .ZN(n689) );
  AND2_X1 U609 ( .A1(n500), .A2(n689), .ZN(n539) );
  NOR2_X2 U610 ( .A1(n596), .A2(n501), .ZN(n570) );
  XNOR2_X1 U611 ( .A(KEYINPUT113), .B(n570), .ZN(n523) );
  XNOR2_X1 U612 ( .A(G110), .B(KEYINPUT16), .ZN(n502) );
  XNOR2_X1 U613 ( .A(n503), .B(n502), .ZN(n505) );
  XNOR2_X1 U614 ( .A(n505), .B(n504), .ZN(n741) );
  XNOR2_X1 U615 ( .A(n506), .B(n741), .ZN(n516) );
  NAND2_X1 U616 ( .A1(n755), .A2(G224), .ZN(n507) );
  XNOR2_X1 U617 ( .A(n510), .B(n509), .ZN(n514) );
  XNOR2_X1 U618 ( .A(KEYINPUT18), .B(KEYINPUT74), .ZN(n511) );
  XNOR2_X1 U619 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U620 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U621 ( .A(n516), .B(n515), .ZN(n658) );
  NAND2_X1 U622 ( .A1(n518), .A2(n517), .ZN(n520) );
  NAND2_X1 U623 ( .A1(n520), .A2(G210), .ZN(n519) );
  NAND2_X1 U624 ( .A1(n520), .A2(G214), .ZN(n708) );
  INV_X1 U625 ( .A(n708), .ZN(n521) );
  INV_X1 U626 ( .A(n549), .ZN(n522) );
  NOR2_X1 U627 ( .A1(n523), .A2(n522), .ZN(n524) );
  AND2_X1 U628 ( .A1(n755), .A2(G227), .ZN(n525) );
  XNOR2_X1 U629 ( .A(G110), .B(KEYINPUT73), .ZN(n528) );
  XNOR2_X1 U630 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U631 ( .A(KEYINPUT68), .B(G469), .ZN(n533) );
  INV_X1 U632 ( .A(KEYINPUT67), .ZN(n532) );
  XNOR2_X1 U633 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X2 U634 ( .A(n535), .B(n534), .ZN(n609) );
  INV_X1 U635 ( .A(n609), .ZN(n537) );
  INV_X1 U636 ( .A(n539), .ZN(n540) );
  OR2_X1 U637 ( .A1(n595), .A2(n540), .ZN(n560) );
  NOR2_X1 U638 ( .A1(n560), .A2(n575), .ZN(n542) );
  NAND2_X1 U639 ( .A1(n559), .A2(n542), .ZN(n543) );
  INV_X1 U640 ( .A(n557), .ZN(n544) );
  NAND2_X1 U641 ( .A1(n544), .A2(n555), .ZN(n598) );
  XOR2_X1 U642 ( .A(KEYINPUT111), .B(n609), .Z(n548) );
  BUF_X1 U643 ( .A(n583), .Z(n550) );
  AND2_X1 U644 ( .A1(n555), .A2(n557), .ZN(n680) );
  NOR2_X1 U645 ( .A1(n563), .A2(n680), .ZN(n707) );
  INV_X1 U646 ( .A(n707), .ZN(n551) );
  NOR2_X1 U647 ( .A1(n552), .A2(KEYINPUT47), .ZN(n553) );
  INV_X1 U648 ( .A(n555), .ZN(n556) );
  NAND2_X1 U649 ( .A1(n557), .A2(n556), .ZN(n711) );
  NAND2_X1 U650 ( .A1(n709), .A2(n708), .ZN(n706) );
  NAND2_X1 U651 ( .A1(n561), .A2(n709), .ZN(n562) );
  XNOR2_X1 U652 ( .A(KEYINPUT39), .B(n562), .ZN(n569) );
  NAND2_X1 U653 ( .A1(n569), .A2(n563), .ZN(n564) );
  XNOR2_X1 U654 ( .A(n565), .B(KEYINPUT46), .ZN(n566) );
  XNOR2_X1 U655 ( .A(KEYINPUT48), .B(KEYINPUT85), .ZN(n568) );
  AND2_X1 U656 ( .A1(n680), .A2(n569), .ZN(n686) );
  NAND2_X1 U657 ( .A1(n570), .A2(n708), .ZN(n571) );
  XOR2_X1 U658 ( .A(KEYINPUT106), .B(n571), .Z(n572) );
  NAND2_X1 U659 ( .A1(n572), .A2(n691), .ZN(n574) );
  XOR2_X1 U660 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n573) );
  XNOR2_X1 U661 ( .A(n574), .B(n573), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U663 ( .A(n577), .B(KEYINPUT108), .ZN(n767) );
  INV_X1 U664 ( .A(n578), .ZN(n579) );
  NOR2_X1 U665 ( .A1(G898), .A2(n755), .ZN(n742) );
  NAND2_X1 U666 ( .A1(n579), .A2(n742), .ZN(n580) );
  AND2_X1 U667 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U668 ( .A(n711), .ZN(n585) );
  INV_X1 U669 ( .A(KEYINPUT70), .ZN(n586) );
  XNOR2_X1 U670 ( .A(n586), .B(KEYINPUT22), .ZN(n587) );
  XOR2_X1 U671 ( .A(KEYINPUT104), .B(n595), .Z(n688) );
  NOR2_X1 U672 ( .A1(n688), .A2(n589), .ZN(n590) );
  INV_X1 U673 ( .A(n699), .ZN(n591) );
  NAND2_X1 U674 ( .A1(n591), .A2(n595), .ZN(n592) );
  NOR2_X1 U675 ( .A1(n592), .A2(n601), .ZN(n593) );
  INV_X1 U676 ( .A(n689), .ZN(n594) );
  INV_X1 U677 ( .A(n610), .ZN(n692) );
  XOR2_X1 U678 ( .A(KEYINPUT86), .B(n600), .Z(n604) );
  INV_X1 U679 ( .A(n688), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n667) );
  NAND2_X1 U682 ( .A1(n605), .A2(n699), .ZN(n701) );
  NOR2_X1 U683 ( .A1(n606), .A2(n701), .ZN(n607) );
  XOR2_X1 U684 ( .A(KEYINPUT31), .B(n607), .Z(n681) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  OR2_X1 U686 ( .A1(n611), .A2(n699), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n608), .A2(n612), .ZN(n669) );
  NOR2_X1 U688 ( .A1(n681), .A2(n669), .ZN(n613) );
  OR2_X1 U689 ( .A1(n613), .A2(n707), .ZN(n614) );
  AND2_X1 U690 ( .A1(KEYINPUT2), .A2(KEYINPUT83), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n622) );
  INV_X1 U692 ( .A(n622), .ZN(n618) );
  INV_X1 U693 ( .A(n616), .ZN(n617) );
  OR2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n754), .B(KEYINPUT71), .ZN(n619) );
  INV_X1 U696 ( .A(n620), .ZN(n625) );
  INV_X1 U697 ( .A(KEYINPUT83), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n621), .A2(KEYINPUT2), .ZN(n623) );
  AND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U701 ( .A(KEYINPUT64), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n364), .A2(G469), .ZN(n633) );
  XNOR2_X1 U703 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n629) );
  XNOR2_X1 U704 ( .A(n629), .B(KEYINPUT57), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(n635) );
  INV_X1 U706 ( .A(G952), .ZN(n634) );
  NOR2_X2 U707 ( .A1(n635), .A2(n738), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n636), .B(KEYINPUT124), .ZN(G54) );
  NAND2_X1 U709 ( .A1(n363), .A2(G217), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n640), .B(KEYINPUT126), .ZN(G66) );
  XOR2_X1 U711 ( .A(G110), .B(KEYINPUT115), .Z(n641) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(G12) );
  XOR2_X1 U713 ( .A(n643), .B(G122), .Z(G24) );
  XNOR2_X1 U714 ( .A(n644), .B(G119), .ZN(G21) );
  NAND2_X1 U715 ( .A1(n363), .A2(G472), .ZN(n648) );
  XOR2_X1 U716 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n646) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X2 U718 ( .A1(n649), .A2(n738), .ZN(n651) );
  XNOR2_X1 U719 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(G57) );
  NAND2_X1 U721 ( .A1(n364), .A2(G475), .ZN(n655) );
  XNOR2_X1 U722 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U724 ( .A1(n656), .A2(n738), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U726 ( .A1(n364), .A2(G210), .ZN(n663) );
  XNOR2_X1 U727 ( .A(KEYINPUT79), .B(KEYINPUT54), .ZN(n659) );
  XOR2_X1 U728 ( .A(n659), .B(KEYINPUT55), .Z(n660) );
  XNOR2_X1 U729 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X2 U730 ( .A1(n664), .A2(n738), .ZN(n666) );
  XNOR2_X1 U731 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n665) );
  XNOR2_X1 U732 ( .A(n666), .B(n665), .ZN(G51) );
  XNOR2_X1 U733 ( .A(G101), .B(n667), .ZN(G3) );
  NAND2_X1 U734 ( .A1(n678), .A2(n669), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(G104), .ZN(G6) );
  XOR2_X1 U736 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n671) );
  NAND2_X1 U737 ( .A1(n669), .A2(n680), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(G107), .B(n672), .ZN(G9) );
  XOR2_X1 U740 ( .A(G128), .B(KEYINPUT29), .Z(n674) );
  NAND2_X1 U741 ( .A1(n675), .A2(n680), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(G30) );
  XOR2_X1 U743 ( .A(G146), .B(KEYINPUT117), .Z(n677) );
  NAND2_X1 U744 ( .A1(n675), .A2(n678), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n677), .B(n676), .ZN(G48) );
  NAND2_X1 U746 ( .A1(n678), .A2(n681), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n679), .B(G113), .ZN(G15) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(G116), .ZN(G18) );
  XNOR2_X1 U750 ( .A(n683), .B(KEYINPUT118), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n684), .B(KEYINPUT37), .ZN(n685) );
  XNOR2_X1 U752 ( .A(G125), .B(n685), .ZN(G27) );
  XOR2_X1 U753 ( .A(G134), .B(n686), .Z(G36) );
  XOR2_X1 U754 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n733) );
  NOR2_X1 U755 ( .A1(n705), .A2(n715), .ZN(n687) );
  NOR2_X1 U756 ( .A1(n687), .A2(G953), .ZN(n731) );
  NOR2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U758 ( .A(KEYINPUT49), .B(n690), .ZN(n697) );
  NAND2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT120), .B(KEYINPUT50), .Z(n693) );
  XNOR2_X1 U761 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U762 ( .A(KEYINPUT119), .B(n695), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U765 ( .A(n700), .B(KEYINPUT121), .ZN(n702) );
  NAND2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(n703), .ZN(n704) );
  NOR2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n713) );
  NOR2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U772 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U775 ( .A(n718), .B(KEYINPUT52), .ZN(n719) );
  NOR2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n729) );
  NOR2_X1 U777 ( .A1(n744), .A2(KEYINPUT2), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n722), .B(KEYINPUT82), .ZN(n725) );
  INV_X1 U779 ( .A(n754), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n723), .A2(KEYINPUT2), .ZN(n724) );
  NOR2_X1 U781 ( .A1(n725), .A2(n724), .ZN(n727) );
  AND2_X1 U782 ( .A1(n726), .A2(n727), .ZN(n728) );
  NOR2_X1 U783 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U784 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n733), .B(n732), .ZN(G75) );
  NAND2_X1 U786 ( .A1(n363), .A2(G478), .ZN(n736) );
  XOR2_X1 U787 ( .A(KEYINPUT125), .B(n734), .Z(n735) );
  XNOR2_X1 U788 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U789 ( .A1(n738), .A2(n737), .ZN(G63) );
  XOR2_X1 U790 ( .A(n739), .B(G101), .Z(n740) );
  XOR2_X1 U791 ( .A(n741), .B(n740), .Z(n743) );
  NOR2_X1 U792 ( .A1(n743), .A2(n742), .ZN(n750) );
  NAND2_X1 U793 ( .A1(n744), .A2(n755), .ZN(n748) );
  NAND2_X1 U794 ( .A1(G953), .A2(G224), .ZN(n745) );
  XNOR2_X1 U795 ( .A(KEYINPUT61), .B(n745), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n746), .A2(G898), .ZN(n747) );
  NAND2_X1 U797 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U798 ( .A(n750), .B(n749), .ZN(G69) );
  XNOR2_X1 U799 ( .A(n751), .B(KEYINPUT4), .ZN(n753) );
  XNOR2_X1 U800 ( .A(n752), .B(n753), .ZN(n757) );
  XNOR2_X1 U801 ( .A(n754), .B(n757), .ZN(n756) );
  NAND2_X1 U802 ( .A1(n756), .A2(n755), .ZN(n762) );
  XNOR2_X1 U803 ( .A(n757), .B(G227), .ZN(n758) );
  NAND2_X1 U804 ( .A1(n758), .A2(G900), .ZN(n759) );
  XOR2_X1 U805 ( .A(KEYINPUT127), .B(n759), .Z(n760) );
  NAND2_X1 U806 ( .A1(G953), .A2(n760), .ZN(n761) );
  NAND2_X1 U807 ( .A1(n762), .A2(n761), .ZN(G72) );
  XOR2_X1 U808 ( .A(G143), .B(KEYINPUT116), .Z(n763) );
  XNOR2_X1 U809 ( .A(n764), .B(n763), .ZN(G45) );
  XOR2_X1 U810 ( .A(G131), .B(n765), .Z(G33) );
  XOR2_X1 U811 ( .A(n766), .B(G137), .Z(G39) );
  XNOR2_X1 U812 ( .A(G140), .B(n767), .ZN(G42) );
endmodule

