//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n209), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  INV_X1    g0021(.A(KEYINPUT1), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n226), .A2(new_n207), .A3(new_n227), .ZN(new_n228));
  NOR4_X1   g0028(.A1(new_n213), .A2(new_n223), .A3(new_n224), .A4(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G68), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  OAI21_X1  g0049(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(new_n250), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(G226), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(new_n260), .B2(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI211_X1 g0063(.A(new_n252), .B(new_n256), .C1(new_n263), .C2(new_n253), .ZN(new_n264));
  INV_X1    g0064(.A(G179), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT69), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n227), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(new_n273), .B1(new_n202), .B2(new_n269), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n271), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n274), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n267), .B(new_n284), .C1(G169), .C2(new_n264), .ZN(new_n285));
  INV_X1    g0085(.A(G200), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n264), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n264), .A2(G190), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n284), .B(KEYINPUT9), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT10), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT10), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n287), .A2(new_n292), .A3(new_n289), .A4(new_n288), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT3), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(G232), .A4(G1698), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(G226), .A4(new_n258), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G97), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n253), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n252), .B1(new_n255), .B2(G238), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT13), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n302), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G200), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n278), .A2(G77), .ZN(new_n310));
  INV_X1    g0110(.A(new_n280), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n310), .B1(new_n207), .B2(G68), .C1(new_n202), .C2(new_n311), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n312), .A2(KEYINPUT11), .A3(new_n271), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT11), .B1(new_n312), .B2(new_n271), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n283), .B1(G1), .B2(new_n207), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT12), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n269), .B2(new_n244), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n315), .A2(new_n244), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n313), .A2(new_n314), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n309), .B(new_n320), .C1(new_n321), .C2(new_n308), .ZN(new_n322));
  INV_X1    g0122(.A(G238), .ZN(new_n323));
  INV_X1    g0123(.A(G107), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n261), .A2(new_n323), .B1(new_n324), .B2(new_n257), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n296), .A2(new_n297), .ZN(new_n326));
  INV_X1    g0126(.A(G232), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n326), .A2(new_n327), .A3(G1698), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n253), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n252), .B1(new_n255), .B2(G244), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n276), .A2(new_n280), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n283), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n269), .A2(new_n260), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n315), .B2(new_n260), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n332), .A2(G169), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n331), .A2(G179), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n337), .A2(new_n339), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n331), .B2(new_n321), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(G200), .B2(new_n331), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n285), .A2(new_n294), .A3(new_n322), .A4(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n252), .B1(new_n255), .B2(G232), .ZN(new_n348));
  INV_X1    g0148(.A(new_n296), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT70), .A2(G33), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT70), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n352), .B2(KEYINPUT3), .ZN(new_n353));
  MUX2_X1   g0153(.A(G223), .B(G226), .S(G1698), .Z(new_n354));
  AOI22_X1  g0154(.A1(new_n353), .A2(new_n354), .B1(G33), .B2(G87), .ZN(new_n355));
  INV_X1    g0155(.A(new_n227), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G41), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(G190), .B(new_n348), .C1(new_n355), .C2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n277), .ZN(new_n361));
  NAND2_X1  g0161(.A1(KEYINPUT70), .A2(G33), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(KEYINPUT3), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n354), .A2(new_n363), .A3(new_n296), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n358), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n358), .A2(new_n250), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n367), .A2(new_n327), .B1(new_n251), .B2(new_n250), .ZN(new_n368));
  OAI21_X1  g0168(.A(G200), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  INV_X1    g0171(.A(G159), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n311), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n280), .A2(KEYINPUT71), .A3(G159), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G58), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n244), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n377), .B2(new_n201), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(G20), .B1(new_n363), .B2(new_n296), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n353), .A2(KEYINPUT7), .A3(G20), .ZN(new_n383));
  OAI211_X1 g0183(.A(KEYINPUT16), .B(new_n379), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT16), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n381), .A2(G20), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT3), .B1(new_n361), .B2(new_n362), .ZN(new_n387));
  INV_X1    g0187(.A(new_n297), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n381), .B1(new_n257), .B2(G20), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n244), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n375), .A2(new_n378), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n385), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n384), .A2(new_n393), .A3(new_n271), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n315), .A2(new_n276), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n275), .A2(new_n268), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n370), .A2(new_n394), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n394), .A2(new_n399), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT73), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n265), .B(new_n348), .C1(new_n355), .C2(new_n358), .ZN(new_n404));
  INV_X1    g0204(.A(G169), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n366), .B2(new_n368), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n403), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  INV_X1    g0211(.A(new_n409), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n407), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n402), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n401), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n307), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n306), .B1(new_n302), .B2(new_n303), .ZN(new_n418));
  OAI21_X1  g0218(.A(G169), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n308), .A2(new_n421), .A3(G169), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n305), .A2(G179), .A3(new_n307), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n320), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n347), .A2(new_n416), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G41), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n429), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT75), .B1(new_n429), .B2(KEYINPUT5), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n251), .B1(new_n356), .B2(new_n357), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n206), .B(G45), .C1(new_n429), .C2(KEYINPUT5), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT74), .ZN(new_n435));
  INV_X1    g0235(.A(G45), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(G1), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT74), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT5), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G41), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n432), .A2(new_n433), .A3(new_n435), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT75), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n439), .B2(G41), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n429), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n437), .A4(new_n440), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(G270), .A3(new_n358), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(G264), .A2(G1698), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n363), .A2(new_n296), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n326), .A2(G303), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT81), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n353), .A2(new_n454), .A3(G257), .A4(new_n258), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n363), .A2(G257), .A3(new_n258), .A4(new_n296), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n453), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n449), .B1(new_n458), .B2(new_n358), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n268), .A2(G116), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n206), .A2(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n283), .A2(new_n268), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n463), .B2(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n207), .C1(G33), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G20), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n271), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT20), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n405), .B1(new_n464), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n459), .A2(KEYINPUT21), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n459), .A2(KEYINPUT82), .A3(KEYINPUT21), .A4(new_n473), .ZN(new_n477));
  INV_X1    g0277(.A(new_n453), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n448), .B1(new_n481), .B2(new_n253), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n464), .A2(new_n472), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(G179), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT83), .B(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(G169), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n476), .A2(new_n477), .A3(new_n484), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n483), .B1(new_n459), .B2(G200), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(G190), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n446), .A2(G264), .A3(new_n358), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT84), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n446), .A2(KEYINPUT84), .A3(G264), .A4(new_n358), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n363), .A2(new_n296), .ZN(new_n497));
  INV_X1    g0297(.A(G250), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n258), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G257), .B2(new_n258), .ZN(new_n500));
  INV_X1    g0300(.A(G294), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n497), .A2(new_n500), .B1(new_n501), .B2(new_n352), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n495), .A2(new_n496), .B1(new_n502), .B2(new_n253), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n405), .B1(new_n503), .B2(new_n442), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n495), .A2(new_n496), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n253), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(new_n442), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n504), .A2(KEYINPUT85), .B1(new_n507), .B2(G179), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT85), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n507), .B2(new_n405), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT25), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n268), .B2(G107), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n268), .A2(new_n512), .A3(G107), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n463), .A2(G107), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n207), .B(G116), .C1(new_n350), .C2(new_n351), .ZN(new_n518));
  OR3_X1    g0318(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G87), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(G20), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT22), .B1(new_n257), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n522), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n363), .A2(new_n207), .A3(new_n296), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n521), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n529), .B(KEYINPUT24), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n517), .B1(new_n530), .B2(new_n271), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n505), .A2(new_n442), .A3(new_n506), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT24), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n524), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n538), .B2(new_n528), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n271), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n503), .A2(G190), .A3(new_n442), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n540), .A2(new_n541), .A3(new_n516), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n511), .A2(new_n532), .B1(new_n534), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n363), .A2(G244), .A3(G1698), .A4(new_n296), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n363), .A2(G238), .A3(new_n258), .A4(new_n296), .ZN(new_n545));
  OAI21_X1  g0345(.A(G116), .B1(new_n350), .B2(new_n351), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n253), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n358), .B(G250), .C1(G1), .C2(new_n436), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n437), .A2(G274), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT80), .B1(new_n553), .B2(new_n321), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(G200), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n547), .B2(new_n253), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT80), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(G190), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n334), .A2(new_n268), .ZN(new_n559));
  OR2_X1    g0359(.A1(KEYINPUT78), .A2(G87), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT78), .A2(G87), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n207), .B1(new_n300), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n563), .A2(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n363), .A2(new_n207), .A3(G68), .A4(new_n296), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n559), .B1(new_n569), .B2(new_n271), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n463), .A2(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n554), .A2(new_n555), .A3(new_n558), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(G169), .B1(new_n548), .B2(new_n552), .ZN(new_n575));
  AOI211_X1 g0375(.A(G179), .B(new_n551), .C1(new_n547), .C2(new_n253), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT77), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n569), .A2(new_n271), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n462), .A2(new_n333), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n559), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n570), .A2(KEYINPUT79), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n548), .A2(new_n265), .A3(new_n552), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT77), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n587), .B(new_n588), .C1(G169), .C2(new_n556), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n577), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n446), .A2(G257), .A3(new_n358), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n442), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(KEYINPUT4), .A2(G244), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n296), .A2(new_n297), .A3(new_n593), .A4(new_n258), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n296), .A2(new_n297), .A3(G250), .A4(G1698), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n465), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT4), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n363), .A2(G244), .A3(new_n258), .A4(new_n296), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n592), .B(new_n265), .C1(new_n599), .C2(new_n358), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT76), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n442), .A2(new_n591), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n597), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n594), .A2(new_n595), .A3(new_n465), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n605), .B2(new_n253), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT76), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n265), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n358), .B1(new_n603), .B2(new_n604), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n405), .B1(new_n609), .B2(new_n602), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n324), .B1(new_n389), .B2(new_n390), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT6), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n612), .A2(new_n466), .A3(G107), .ZN(new_n613));
  XNOR2_X1  g0413(.A(G97), .B(G107), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n615), .A2(new_n207), .B1(new_n260), .B2(new_n311), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n271), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n269), .A2(new_n466), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n463), .A2(G97), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n601), .A2(new_n608), .A3(new_n610), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n618), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n389), .A2(new_n390), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G107), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n614), .A2(new_n612), .ZN(new_n625));
  INV_X1    g0425(.A(new_n613), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n622), .B1(new_n629), .B2(new_n271), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n606), .A2(G190), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n630), .B(new_n631), .C1(new_n286), .C2(new_n606), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n574), .A2(new_n590), .A3(new_n621), .A4(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n428), .A2(new_n492), .A3(new_n543), .A4(new_n633), .ZN(G372));
  AND2_X1   g0434(.A1(new_n411), .A2(new_n415), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n322), .ZN(new_n637));
  INV_X1    g0437(.A(new_n342), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n426), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n636), .B1(new_n639), .B2(new_n401), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT88), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n294), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n291), .A2(KEYINPUT88), .A3(new_n293), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n285), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n534), .A2(new_n540), .A3(new_n541), .A4(new_n516), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n621), .A2(new_n632), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n558), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n557), .B1(new_n556), .B2(G190), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n650), .A2(new_n651), .A3(new_n572), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n547), .A2(KEYINPUT86), .A3(new_n253), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT86), .B1(new_n547), .B2(new_n253), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n552), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G200), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n576), .B1(new_n584), .B2(new_n585), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n405), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n652), .A2(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n531), .B1(new_n508), .B2(new_n510), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n649), .B(new_n659), .C1(new_n488), .C2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT87), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n610), .B1(new_n600), .B2(KEYINPUT76), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n607), .B1(new_n606), .B2(new_n265), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n601), .A2(new_n608), .A3(KEYINPUT87), .A4(new_n610), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n665), .A2(new_n620), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n659), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT86), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n548), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n547), .A2(KEYINPUT86), .A3(new_n253), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(G169), .B1(new_n673), .B2(new_n552), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT79), .B1(new_n570), .B2(new_n580), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n283), .B1(new_n567), .B2(new_n568), .ZN(new_n676));
  NOR4_X1   g0476(.A1(new_n676), .A2(new_n579), .A3(new_n583), .A4(new_n559), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n587), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n621), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n590), .A3(new_n574), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n681), .B2(KEYINPUT26), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n661), .A2(new_n669), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n428), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n647), .A2(new_n684), .ZN(G369));
  NAND3_X1  g0485(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G343), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n543), .B1(new_n531), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n660), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  INV_X1    g0494(.A(new_n691), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n483), .A2(new_n695), .ZN(new_n696));
  MUX2_X1   g0496(.A(new_n488), .B(new_n492), .S(new_n696), .Z(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n697), .A3(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n660), .A2(new_n691), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n488), .A2(new_n691), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n543), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n210), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G1), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n563), .A2(G116), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(new_n226), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n683), .A2(new_n711), .A3(new_n691), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n649), .A2(new_n659), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n488), .A2(new_n660), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n665), .A2(new_n620), .A3(new_n666), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n554), .A2(new_n558), .A3(new_n573), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n286), .B1(new_n673), .B2(new_n552), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n674), .B2(new_n678), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT26), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n679), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n680), .A2(new_n590), .A3(new_n668), .A4(new_n574), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n715), .B1(new_n723), .B2(KEYINPUT91), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n720), .A2(new_n725), .A3(new_n721), .A4(new_n722), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n695), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n712), .B1(new_n727), .B2(new_n711), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n492), .A2(new_n633), .A3(new_n543), .A4(new_n691), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT90), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n655), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n265), .B1(new_n609), .B2(new_n602), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n507), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(KEYINPUT90), .B(new_n552), .C1(new_n653), .C2(new_n654), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n731), .A2(new_n733), .A3(new_n459), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n605), .A2(new_n253), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n503), .A2(new_n736), .A3(new_n556), .A4(new_n592), .ZN(new_n737));
  OAI211_X1 g0537(.A(G179), .B(new_n449), .C1(new_n458), .C2(new_n358), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT89), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT89), .B(new_n741), .C1(new_n737), .C2(new_n738), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n735), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n695), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n729), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n728), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n710), .B1(new_n751), .B2(G1), .ZN(G364));
  AND2_X1   g0552(.A1(new_n207), .A2(G13), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n206), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n705), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n697), .B2(G330), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G330), .B2(new_n697), .ZN(new_n758));
  INV_X1    g0558(.A(new_n756), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n227), .B1(G20), .B2(new_n405), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n207), .B1(new_n762), .B2(G190), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n466), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n207), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n762), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G159), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n207), .A2(new_n265), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n771), .A2(G190), .A3(new_n286), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n764), .B(new_n769), .C1(G68), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n286), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G20), .A3(G190), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n560), .B2(new_n562), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n765), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n326), .B(new_n776), .C1(G107), .C2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n780), .A2(KEYINPUT95), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(KEYINPUT95), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G50), .ZN(new_n785));
  AOI21_X1  g0585(.A(G200), .B1(new_n771), .B2(KEYINPUT94), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(KEYINPUT94), .B2(new_n771), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n321), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(G190), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G58), .A2(new_n788), .B1(new_n789), .B2(G77), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n773), .A2(new_n779), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G311), .A2(new_n789), .B1(new_n788), .B2(G322), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n784), .A2(G326), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n777), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G303), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n326), .B1(new_n775), .B2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n795), .B(new_n797), .C1(G329), .C2(new_n767), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  INV_X1    g0599(.A(new_n763), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n772), .A2(new_n799), .B1(G294), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n792), .A2(new_n793), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n761), .B1(new_n791), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G13), .A2(G33), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT93), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n760), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n248), .A2(new_n436), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n704), .A2(new_n353), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n226), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(new_n436), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n810), .B1(new_n814), .B2(KEYINPUT92), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(KEYINPUT92), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n704), .A2(new_n326), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G355), .B1(new_n468), .B2(new_n704), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n759), .B(new_n803), .C1(new_n809), .C2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n697), .B2(new_n807), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n758), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT96), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  NAND2_X1  g0624(.A1(new_n683), .A2(new_n691), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n342), .A2(new_n691), .ZN(new_n826));
  INV_X1    g0626(.A(new_n343), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n345), .B1(new_n827), .B2(new_n695), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n828), .B2(new_n342), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n829), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n683), .A2(new_n691), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n756), .B1(new_n833), .B2(new_n749), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n749), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n760), .A2(new_n804), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n759), .B1(new_n260), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n775), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G107), .B1(new_n767), .B2(G311), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n778), .A2(G87), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n326), .A3(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n764), .B(new_n841), .C1(G283), .C2(new_n772), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G294), .A2(new_n788), .B1(new_n784), .B2(G303), .ZN(new_n843));
  INV_X1    g0643(.A(new_n789), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n842), .B(new_n843), .C1(new_n468), .C2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n784), .A2(G137), .B1(G150), .B2(new_n772), .ZN(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  INV_X1    g0647(.A(new_n788), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n846), .B1(new_n847), .B2(new_n848), .C1(new_n372), .C2(new_n844), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n775), .A2(new_n202), .B1(new_n777), .B2(new_n244), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n353), .B1(new_n376), .B2(new_n763), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(G132), .C2(new_n767), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n849), .B2(new_n850), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n845), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT97), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n837), .B1(new_n805), .B2(new_n831), .C1(new_n857), .C2(new_n761), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n835), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  OR2_X1    g0660(.A1(new_n627), .A2(KEYINPUT35), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n627), .A2(KEYINPUT35), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n227), .A2(new_n207), .A3(new_n468), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT36), .Z(new_n865));
  OR3_X1    g0665(.A1(new_n226), .A2(new_n260), .A3(new_n377), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n206), .B(G13), .C1(new_n866), .C2(new_n243), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n385), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n271), .A3(new_n384), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n399), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n413), .B2(new_n690), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n870), .B1(new_n875), .B2(new_n400), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n370), .A2(new_n394), .A3(new_n399), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n402), .B2(new_n413), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n402), .A2(new_n690), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(KEYINPUT99), .A3(new_n870), .A4(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n410), .A2(new_n879), .A3(new_n870), .A4(new_n400), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT99), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n876), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n874), .A2(new_n690), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n635), .B2(new_n401), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n410), .A2(new_n400), .A3(new_n879), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n881), .A2(new_n882), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n881), .A2(new_n882), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n416), .A2(new_n402), .A3(new_n690), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n869), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n426), .A2(KEYINPUT98), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT98), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n424), .A2(new_n898), .A3(new_n425), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n691), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n887), .B1(new_n884), .B2(new_n886), .ZN(new_n903));
  INV_X1    g0703(.A(new_n876), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n891), .B2(new_n892), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n416), .A2(new_n690), .A3(new_n874), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT38), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n903), .A2(new_n907), .A3(KEYINPUT39), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n896), .A2(new_n902), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n425), .A2(new_n695), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n637), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n897), .A2(new_n912), .A3(new_n899), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n424), .A2(new_n911), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n832), .B2(new_n826), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n903), .A2(new_n907), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n917), .A2(new_n918), .B1(new_n636), .B2(new_n689), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT101), .ZN(new_n921));
  INV_X1    g0721(.A(new_n712), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n668), .B1(new_n667), .B2(new_n659), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n722), .A2(new_n721), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT91), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n661), .A3(new_n726), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n691), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n927), .B2(KEYINPUT29), .ZN(new_n928));
  INV_X1    g0728(.A(new_n428), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT100), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT100), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n711), .B1(new_n926), .B2(new_n691), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n931), .B(new_n428), .C1(new_n932), .C2(new_n922), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n646), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n921), .B(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n829), .B1(new_n913), .B2(new_n914), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n748), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n918), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n748), .A2(new_n937), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n880), .A2(new_n883), .B1(KEYINPUT37), .B2(new_n889), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n879), .B1(new_n635), .B2(new_n401), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n887), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n940), .B1(new_n907), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n939), .B1(new_n944), .B2(new_n936), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n428), .A2(new_n748), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(G330), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n935), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n206), .B2(new_n753), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n935), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n868), .B1(new_n951), .B2(new_n952), .ZN(G367));
  NOR2_X1   g0753(.A1(new_n630), .A2(new_n691), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n665), .A2(new_n666), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT102), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n621), .A2(new_n632), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(new_n956), .C1(new_n957), .C2(new_n954), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n956), .B2(new_n955), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT42), .B1(new_n959), .B2(new_n702), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n621), .B1(new_n959), .B2(new_n693), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(KEYINPUT103), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n691), .B1(new_n961), .B2(KEYINPUT103), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT104), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n959), .A2(new_n702), .A3(KEYINPUT42), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n964), .B2(KEYINPUT104), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n572), .A2(new_n695), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n659), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n721), .B2(new_n968), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n965), .A2(new_n967), .B1(KEYINPUT43), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n698), .A2(new_n959), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT105), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n976), .A2(KEYINPUT43), .A3(new_n970), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(KEYINPUT43), .B2(new_n970), .ZN(new_n978));
  XNOR2_X1  g0778(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n705), .B(new_n979), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n702), .A2(new_n699), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n959), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT44), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n982), .A2(new_n959), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT45), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n984), .A2(new_n698), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n698), .B1(new_n984), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n702), .B1(new_n694), .B2(new_n701), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n697), .A2(G330), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n751), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n751), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n981), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n754), .B(KEYINPUT107), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n977), .A2(new_n978), .A3(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n809), .B1(new_n210), .B2(new_n333), .C1(new_n236), .C2(new_n812), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1002), .A2(new_n756), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G283), .A2(new_n789), .B1(new_n784), .B2(G311), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n775), .A2(new_n468), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT46), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n772), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1007), .A2(new_n501), .B1(new_n763), .B2(new_n324), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n497), .B1(new_n466), .B2(new_n777), .C1(new_n1009), .C2(new_n766), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1004), .B(new_n1011), .C1(new_n796), .C2(new_n848), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G50), .A2(new_n789), .B1(new_n784), .B2(G143), .ZN(new_n1013));
  INV_X1    g0813(.A(G150), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1013), .B1(new_n1014), .B2(new_n848), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(KEYINPUT108), .B(G137), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n775), .A2(new_n376), .B1(new_n766), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT109), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n257), .B1(new_n777), .B2(new_n260), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G159), .B2(new_n772), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(new_n244), .C2(new_n763), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1012), .B1(new_n1015), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT47), .Z(new_n1023));
  OAI221_X1 g0823(.A(new_n1003), .B1(new_n970), .B2(new_n807), .C1(new_n761), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1001), .A2(new_n1024), .ZN(G387));
  AOI22_X1  g0825(.A1(new_n817), .A2(new_n708), .B1(new_n324), .B2(new_n704), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n708), .B(KEYINPUT110), .Z(new_n1027));
  OAI21_X1  g0827(.A(new_n436), .B1(new_n244), .B2(new_n260), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n276), .A2(new_n202), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(KEYINPUT50), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(KEYINPUT50), .B2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n811), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT111), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1032), .A2(new_n1033), .B1(new_n436), .B2(new_n233), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1036), .A2(new_n809), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G50), .A2(new_n788), .B1(new_n789), .B2(G68), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n775), .A2(new_n260), .B1(new_n777), .B2(new_n466), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G150), .B2(new_n767), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n353), .B1(new_n333), .B2(new_n763), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n276), .B2(new_n772), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n784), .A2(G159), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n838), .A2(G294), .B1(new_n800), .B2(G283), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G317), .A2(new_n788), .B1(new_n784), .B2(G322), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n789), .A2(G303), .B1(G311), .B2(new_n772), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT112), .Z(new_n1051));
  NAND2_X1  g0851(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(KEYINPUT49), .A3(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n778), .A2(G116), .B1(new_n767), .B2(G326), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n497), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT49), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1044), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n759), .B(new_n1037), .C1(new_n1057), .C2(new_n760), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n694), .A2(new_n807), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n999), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1058), .A2(new_n1059), .B1(new_n994), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n995), .A2(new_n705), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n751), .A2(new_n994), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(G393));
  NAND2_X1  g0864(.A1(new_n959), .A2(new_n808), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n809), .B1(new_n466), .B2(new_n210), .C1(new_n242), .C2(new_n812), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT113), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n756), .A3(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n848), .A2(new_n372), .B1(new_n1014), .B2(new_n783), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n840), .B1(new_n244), .B2(new_n775), .C1(new_n847), .C2(new_n766), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n353), .B1(new_n260), .B2(new_n763), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n844), .A2(new_n275), .B1(new_n202), .B2(new_n1007), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT114), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1073), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1072), .B(new_n1077), .C1(new_n1076), .C2(new_n1075), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT115), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G311), .A2(new_n788), .B1(new_n784), .B2(G317), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  OAI22_X1  g0883(.A1(new_n1007), .A2(new_n796), .B1(new_n763), .B2(new_n468), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n838), .A2(G283), .B1(new_n767), .B2(G322), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1085), .B(new_n326), .C1(new_n324), .C2(new_n777), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(G294), .C2(new_n789), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1080), .A2(new_n1081), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1070), .B1(new_n1089), .B2(new_n760), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n989), .A2(new_n1060), .B1(new_n1065), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n990), .A2(new_n995), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n705), .B1(new_n990), .B2(new_n995), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(G390));
  NAND2_X1  g0895(.A1(new_n750), .A2(new_n937), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n943), .A2(new_n907), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n901), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n828), .A2(new_n342), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n826), .B1(new_n927), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1099), .B1(new_n1101), .B2(new_n915), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n832), .A2(new_n826), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n915), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n896), .A2(new_n908), .B1(new_n1104), .B2(new_n901), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1097), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n902), .B1(new_n943), .B2(new_n907), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1100), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n727), .A2(new_n1108), .B1(new_n342), .B2(new_n691), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1109), .B2(new_n916), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n896), .A2(new_n908), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1104), .A2(new_n901), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n1113), .A3(new_n1096), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1111), .A2(new_n804), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n836), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n756), .B1(new_n276), .B2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G116), .A2(new_n788), .B1(new_n784), .B2(G283), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1007), .A2(new_n324), .B1(new_n763), .B2(new_n260), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n326), .B1(new_n777), .B2(new_n244), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n775), .A2(new_n522), .B1(new_n766), .B2(new_n501), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1119), .B(new_n1123), .C1(new_n466), .C2(new_n844), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1016), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n789), .A2(new_n1126), .B1(new_n772), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT117), .Z(new_n1129));
  AOI22_X1  g0929(.A1(G132), .A2(new_n788), .B1(new_n784), .B2(G128), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n257), .B1(new_n777), .B2(new_n202), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G125), .B2(new_n767), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n838), .A2(G150), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1133), .A2(KEYINPUT53), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1133), .A2(KEYINPUT53), .B1(G159), .B2(new_n800), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1130), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1124), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1118), .B1(new_n1137), .B2(new_n760), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1115), .A2(new_n1060), .B1(new_n1116), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n929), .A2(new_n749), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n646), .B(new_n1140), .C1(new_n930), .C2(new_n933), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1103), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n916), .B1(new_n749), .B2(new_n829), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1096), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1096), .A2(new_n1143), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1109), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n706), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1115), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1150), .A2(KEYINPUT116), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT116), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1139), .B1(new_n1152), .B2(new_n1153), .ZN(G378));
  NAND2_X1  g0954(.A1(new_n644), .A2(new_n285), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n284), .A2(new_n690), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n643), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT88), .B1(new_n291), .B2(new_n293), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n285), .B(new_n1156), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1158), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1162), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1161), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1156), .B1(new_n644), .B2(new_n285), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n940), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n936), .B1(new_n1098), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n748), .A2(new_n937), .A3(new_n936), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n907), .B2(new_n903), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1168), .B(G330), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1168), .B1(new_n945), .B2(G330), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n920), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT119), .ZN(new_n1177));
  OAI21_X1  g0977(.A(G330), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1168), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n920), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1173), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1176), .A2(new_n1177), .A3(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(KEYINPUT119), .A4(new_n1173), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n1060), .A3(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n772), .A2(G97), .B1(G68), .B2(new_n800), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n353), .A2(G41), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n778), .A2(G58), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n838), .A2(G77), .B1(new_n767), .B2(G283), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n848), .A2(new_n324), .B1(new_n468), .B2(new_n783), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n334), .C2(new_n789), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1193));
  INV_X1    g0993(.A(new_n1187), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G50), .B1(new_n277), .B2(new_n429), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1192), .A2(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n838), .A2(new_n1126), .B1(new_n800), .B2(G150), .ZN(new_n1197));
  INV_X1    g0997(.A(G132), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1007), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n789), .A2(G137), .ZN(new_n1200));
  INV_X1    g1000(.A(G128), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n848), .B2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1199), .B(new_n1202), .C1(G125), .C2(new_n784), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n778), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1196), .B1(new_n1193), .B2(new_n1192), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n760), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n759), .B1(new_n202), .B2(new_n836), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n1168), .C2(new_n805), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1185), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1140), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n933), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n931), .B1(new_n728), .B2(new_n428), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n647), .B(new_n1215), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1115), .B2(new_n1147), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1180), .A2(new_n1181), .A3(new_n1173), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1181), .B1(new_n1180), .B2(new_n1173), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n705), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1141), .B1(new_n1149), .B2(new_n1146), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1223), .B1(new_n1227), .B2(KEYINPUT120), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT120), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1225), .A2(new_n1229), .A3(new_n1226), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1214), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(G375));
  OAI22_X1  g1032(.A1(new_n775), .A2(new_n372), .B1(new_n766), .B2(new_n1201), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT122), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n1198), .B2(new_n783), .C1(new_n844), .C2(new_n1014), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n788), .A2(new_n1127), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n497), .B1(G58), .B2(new_n778), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT121), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n772), .A2(new_n1126), .B1(G50), .B2(new_n800), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(KEYINPUT121), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n324), .A2(new_n844), .B1(new_n848), .B2(new_n794), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n775), .A2(new_n466), .B1(new_n766), .B2(new_n796), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n257), .B(new_n1243), .C1(G77), .C2(new_n778), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n772), .A2(G116), .B1(new_n334), .B2(new_n800), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n501), .C2(new_n783), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1235), .A2(new_n1241), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n760), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1248), .B(new_n756), .C1(G68), .C2(new_n1117), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n916), .B2(new_n804), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1147), .B2(new_n1060), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1148), .A2(new_n981), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(G381));
  INV_X1    g1054(.A(G390), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n859), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G396), .A2(new_n1256), .A3(G393), .A4(G381), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1139), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1231), .A2(new_n1260), .ZN(new_n1261));
  OR3_X1    g1061(.A1(new_n1257), .A2(G387), .A3(new_n1261), .ZN(G407));
  OAI211_X1 g1062(.A(G407), .B(G213), .C1(G343), .C2(new_n1261), .ZN(G409));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(G2897), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1218), .A2(KEYINPUT60), .A3(new_n1146), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT123), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1218), .A2(new_n1270), .A3(KEYINPUT60), .A4(new_n1146), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n706), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1269), .A2(new_n1271), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(G384), .A3(new_n1251), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1275), .B2(new_n1251), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(new_n1251), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n859), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT125), .B1(new_n1282), .B2(new_n1276), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1267), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1276), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G2897), .B(new_n1266), .C1(new_n1285), .C2(new_n1279), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1227), .A2(KEYINPUT120), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1223), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1230), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1214), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(G378), .A3(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1225), .A2(new_n980), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1060), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1294), .A2(new_n1213), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1259), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1266), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1264), .B1(new_n1287), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT126), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1301), .B(new_n1264), .C1(new_n1287), .C2(new_n1298), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1296), .B1(new_n1231), .B2(G378), .ZN(new_n1303));
  NOR4_X1   g1103(.A1(new_n1303), .A2(KEYINPUT62), .A3(new_n1266), .A4(new_n1285), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1298), .B2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1300), .A2(new_n1302), .A3(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(G393), .B(new_n823), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1001), .A2(new_n1024), .A3(G390), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G390), .B1(new_n1001), .B2(new_n1024), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1311), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1314), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1309), .A2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(KEYINPUT61), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1303), .A2(new_n1266), .A3(new_n1285), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1321), .A2(KEYINPUT63), .ZN(new_n1322));
  OAI21_X1  g1122(.A(KEYINPUT124), .B1(new_n1303), .B2(new_n1266), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT124), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1298), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1323), .A2(new_n1325), .A3(new_n1284), .A4(new_n1286), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1321), .A2(KEYINPUT63), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1320), .A2(new_n1322), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1319), .A2(new_n1328), .ZN(G405));
  INV_X1    g1129(.A(KEYINPUT127), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1292), .B1(new_n1330), .B2(new_n1285), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1231), .A2(new_n1259), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1333), .B1(KEYINPUT127), .B2(new_n1306), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1330), .B(new_n1285), .C1(new_n1331), .C2(new_n1332), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1318), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1336), .B(new_n1337), .ZN(G402));
endmodule


