//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT23), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n203), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(KEYINPUT23), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT24), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n219), .A2(new_n220), .A3(G190gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n209), .B(new_n213), .C1(new_n218), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n225), .B2(new_n207), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n215), .A2(new_n217), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n203), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT27), .B(G183gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(KEYINPUT28), .A3(new_n228), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT27), .B1(new_n219), .B2(new_n220), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(G190gat), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(new_n238), .B2(KEYINPUT28), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n204), .A2(new_n205), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(KEYINPUT26), .B2(new_n208), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n210), .A2(new_n242), .A3(new_n212), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n241), .A2(new_n243), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n239), .A2(KEYINPUT66), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT66), .B1(new_n239), .B2(new_n244), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n232), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n248), .A2(KEYINPUT1), .ZN(new_n249));
  XOR2_X1   g048(.A(G127gat), .B(G134gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n233), .A2(KEYINPUT28), .A3(new_n228), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT27), .ZN(new_n255));
  OR2_X1    g054(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n228), .B1(new_n258), .B2(new_n236), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n243), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n214), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n253), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n239), .A2(KEYINPUT66), .A3(new_n244), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n231), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n249), .B(new_n250), .Z(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G227gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n202), .B1(new_n273), .B2(KEYINPUT34), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n264), .A2(new_n265), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n267), .B1(new_n275), .B2(new_n232), .ZN(new_n276));
  AOI211_X1 g075(.A(new_n251), .B(new_n231), .C1(new_n264), .C2(new_n265), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT34), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(KEYINPUT70), .A3(new_n279), .A4(new_n272), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(KEYINPUT34), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n274), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n272), .B1(new_n252), .B2(new_n268), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT67), .B1(new_n283), .B2(KEYINPUT33), .ZN(new_n284));
  XNOR2_X1  g083(.A(G15gat), .B(G43gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G71gat), .B(G99gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n271), .B1(new_n276), .B2(new_n277), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(KEYINPUT32), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT33), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n284), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n291), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n294), .B2(new_n287), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(KEYINPUT32), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n288), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n282), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n282), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n289), .A3(new_n292), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n299), .A4(new_n300), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(KEYINPUT71), .B(new_n282), .C1(new_n293), .C2(new_n301), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n311), .A2(G141gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(G141gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G155gat), .ZN(new_n315));
  INV_X1    g114(.A(G162gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT78), .B(G141gat), .Z(new_n321));
  AOI21_X1  g120(.A(new_n312), .B1(new_n321), .B2(G148gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n317), .B1(new_n310), .B2(new_n318), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n267), .A2(new_n325), .A3(KEYINPUT4), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(new_n251), .B2(new_n324), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n320), .B(new_n331), .C1(new_n322), .C2(new_n323), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n251), .A3(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n326), .A2(new_n327), .A3(new_n329), .A4(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n251), .B(new_n324), .ZN(new_n337));
  INV_X1    g136(.A(new_n327), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n334), .A2(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT6), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n335), .A2(new_n339), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n346), .B1(new_n350), .B2(new_n341), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT6), .A4(new_n347), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT29), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n247), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n239), .A2(new_n244), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n232), .A2(new_n359), .A3(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n362));
  INV_X1    g161(.A(G197gat), .ZN(new_n363));
  INV_X1    g162(.A(G204gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n367));
  NAND2_X1  g166(.A1(G211gat), .A2(G218gat), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT75), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G211gat), .B(G218gat), .Z(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(new_n369), .B2(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n367), .ZN(new_n374));
  NOR2_X1   g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375));
  AND2_X1   g174(.A1(G197gat), .A2(G204gat), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n374), .B(KEYINPUT74), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n371), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n370), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(KEYINPUT75), .A3(new_n377), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n380), .B1(new_n379), .B2(new_n384), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n362), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n381), .B2(new_n372), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(new_n377), .B2(new_n383), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n376), .A2(new_n375), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n382), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AND4_X1   g192(.A1(KEYINPUT75), .A2(new_n393), .A3(new_n377), .A4(new_n372), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT76), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT77), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n361), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n266), .A2(new_n356), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n232), .A2(new_n359), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n357), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  NOR2_X1   g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n404), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n398), .B2(new_n361), .ZN(new_n413));
  INV_X1    g212(.A(new_n408), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(KEYINPUT30), .A3(new_n414), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n355), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n419), .B(KEYINPUT79), .Z(new_n420));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n332), .A2(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n400), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n369), .A2(new_n370), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n381), .A2(new_n372), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n325), .B1(new_n331), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n420), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n387), .A2(new_n397), .A3(new_n422), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n379), .A2(new_n421), .A3(new_n384), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n331), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n419), .B1(new_n432), .B2(new_n324), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n429), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n429), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n428), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G22gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n438));
  INV_X1    g237(.A(G22gat), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(new_n428), .C1(new_n434), .C2(new_n435), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n437), .B2(new_n440), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n443));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n441), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n446), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n440), .B2(KEYINPUT81), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n433), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT80), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n430), .A3(new_n433), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n439), .B1(new_n454), .B2(new_n428), .ZN(new_n455));
  INV_X1    g254(.A(new_n440), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT82), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n450), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n309), .B(new_n418), .C1(new_n448), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT72), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n302), .A2(new_n305), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n301), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n465), .A2(KEYINPUT72), .A3(new_n303), .A4(new_n304), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n464), .A2(KEYINPUT87), .A3(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n413), .A2(new_n414), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n473), .A2(new_n409), .A3(new_n410), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n472), .B(new_n354), .C1(new_n474), .C2(new_n416), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n450), .A3(new_n458), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n447), .B1(new_n441), .B2(new_n442), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n461), .A2(new_n462), .B1(new_n471), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n477), .A2(new_n476), .B1(new_n307), .B2(new_n308), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n472), .B1(new_n480), .B2(new_n418), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT88), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT83), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n448), .B2(new_n459), .ZN(new_n484));
  INV_X1    g283(.A(new_n418), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n477), .A2(KEYINPUT83), .A3(new_n476), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n474), .A2(new_n416), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n326), .A2(new_n333), .A3(new_n329), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n338), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(KEYINPUT39), .C1(new_n338), .C2(new_n337), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n491), .B(new_n346), .C1(KEYINPUT39), .C2(new_n490), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n492), .A2(new_n493), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n488), .A2(new_n348), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n413), .A2(KEYINPUT37), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n414), .B1(new_n413), .B2(KEYINPUT37), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT38), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT86), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n498), .A2(KEYINPUT38), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n361), .A2(new_n398), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n401), .A2(new_n400), .A3(new_n403), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n505), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(KEYINPUT84), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n503), .A2(new_n506), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT37), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n354), .A2(new_n473), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n513), .B(KEYINPUT38), .C1(new_n497), .C2(new_n498), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n500), .A2(new_n511), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n496), .B(new_n515), .C1(new_n448), .C2(new_n459), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n487), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n464), .A2(new_n518), .A3(new_n466), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n309), .A2(KEYINPUT36), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n479), .A2(new_n482), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(G1gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT95), .ZN(new_n531));
  INV_X1    g330(.A(new_n528), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(KEYINPUT94), .B2(new_n526), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n526), .A2(KEYINPUT94), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G43gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(G50gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT92), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n537), .B2(G50gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(new_n537), .A3(G50gat), .ZN(new_n543));
  INV_X1    g342(.A(G50gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(KEYINPUT91), .A3(G43gat), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n539), .A2(new_n541), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n550));
  INV_X1    g349(.A(G36gat), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n550), .A2(KEYINPUT93), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT93), .B1(new_n550), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n538), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n537), .A2(G50gat), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n555), .A2(new_n556), .A3(new_n547), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT90), .B(G29gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(G36gat), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n548), .A2(new_n554), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n550), .A2(new_n551), .ZN(new_n562));
  INV_X1    g361(.A(new_n560), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n562), .B(new_n557), .C1(new_n563), .C2(new_n549), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT17), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n536), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n565), .B1(new_n531), .B2(new_n535), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n574), .A2(KEYINPUT18), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(KEYINPUT18), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT96), .B1(new_n536), .B2(new_n566), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(new_n571), .Z(new_n578));
  XOR2_X1   g377(.A(new_n573), .B(KEYINPUT13), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT89), .B(G197gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(KEYINPUT11), .B(G169gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT12), .Z(new_n587));
  OR2_X1    g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n581), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT99), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT41), .ZN(new_n595));
  XOR2_X1   g394(.A(G134gat), .B(G162gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT101), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n599), .A2(new_n600), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G99gat), .B(G106gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n567), .A3(new_n569), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n607), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n610), .A2(new_n565), .B1(KEYINPUT41), .B2(new_n594), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT102), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n614), .ZN(new_n616));
  AOI211_X1 g415(.A(new_n597), .B(new_n615), .C1(KEYINPUT104), .C2(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(KEYINPUT104), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n619));
  INV_X1    g418(.A(new_n616), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n597), .B1(new_n620), .B2(new_n615), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n617), .A2(new_n618), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n621), .A2(new_n619), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(KEYINPUT9), .ZN(new_n627));
  NOR2_X1   g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  OAI22_X1  g427(.A1(new_n627), .A2(KEYINPUT97), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G57gat), .B(G64gat), .Z(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(KEYINPUT9), .B2(new_n626), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G127gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n632), .B(KEYINPUT98), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n536), .B1(new_n639), .B2(new_n633), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G155gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n624), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT105), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n608), .B(new_n632), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(KEYINPUT10), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n639), .A2(new_n608), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(G230gat), .ZN(new_n655));
  OAI22_X1  g454(.A1(new_n652), .A2(new_n654), .B1(new_n655), .B2(new_n270), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n270), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n650), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n524), .A2(new_n591), .A3(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n669), .A2(KEYINPUT106), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(KEYINPUT106), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n354), .B(KEYINPUT107), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  INV_X1    g475(.A(new_n488), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n529), .B2(new_n678), .ZN(new_n681));
  MUX2_X1   g480(.A(new_n680), .B(new_n681), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g481(.A(new_n471), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n672), .A2(G15gat), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n672), .B2(new_n523), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1326gat));
  NAND2_X1  g485(.A1(new_n484), .A2(new_n486), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT108), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NOR2_X1   g491(.A1(new_n524), .A2(new_n624), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n591), .A2(new_n667), .A3(new_n648), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n674), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n695), .A2(new_n559), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT45), .Z(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n524), .B2(new_n624), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n523), .A2(new_n487), .A3(new_n516), .ZN(new_n701));
  INV_X1    g500(.A(new_n482), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n471), .A2(new_n478), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(KEYINPUT88), .B2(new_n481), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n701), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n624), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(KEYINPUT44), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n700), .A2(new_n707), .A3(new_n694), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n700), .A2(new_n707), .A3(KEYINPUT109), .A4(new_n694), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n559), .B1(new_n712), .B2(new_n696), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n713), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n695), .A2(G36gat), .A3(new_n677), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n712), .B2(new_n677), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G36gat), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n712), .A2(new_n717), .A3(new_n677), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(G1329gat));
  OAI21_X1  g520(.A(G43gat), .B1(new_n708), .B2(new_n523), .ZN(new_n722));
  INV_X1    g521(.A(new_n695), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n537), .A3(new_n471), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n724), .A3(KEYINPUT47), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT112), .Z(new_n726));
  OAI21_X1  g525(.A(G43gat), .B1(new_n712), .B2(new_n523), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT47), .B1(new_n727), .B2(new_n724), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n726), .B1(new_n730), .B2(new_n731), .ZN(G1330gat));
  NOR3_X1   g531(.A1(new_n695), .A2(G50gat), .A3(new_n687), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n448), .A2(new_n459), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G50gat), .B1(new_n708), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(KEYINPUT48), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n710), .A2(new_n688), .A3(new_n711), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G50gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n734), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT113), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n733), .B1(new_n739), .B2(G50gat), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT48), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n738), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT114), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n738), .B(new_n749), .C1(new_n743), .C2(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1331gat));
  INV_X1    g550(.A(new_n667), .ZN(new_n752));
  OR4_X1    g551(.A1(new_n524), .A2(new_n590), .A3(new_n650), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n696), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g554(.A(new_n753), .B(KEYINPUT115), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n757));
  INV_X1    g556(.A(G64gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n488), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT116), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n758), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1333gat));
  INV_X1    g562(.A(new_n523), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n756), .A2(G71gat), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n753), .A2(new_n683), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(G71gat), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n756), .A2(new_n688), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g569(.A1(new_n700), .A2(new_n707), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n752), .A2(new_n590), .A3(new_n648), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n696), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n590), .A2(new_n648), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n776));
  NAND3_X1  g575(.A1(new_n693), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n693), .A2(new_n775), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT117), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n674), .A2(new_n667), .A3(new_n599), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n774), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n773), .B2(new_n677), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n667), .A2(new_n600), .A3(new_n488), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n773), .B2(new_n523), .ZN(new_n789));
  OR3_X1    g588(.A1(new_n683), .A2(G99gat), .A3(new_n752), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n782), .B2(new_n790), .ZN(G1338gat));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n736), .A2(G106gat), .A3(new_n752), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT53), .B1(new_n781), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G106gat), .B1(new_n773), .B2(new_n736), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n795), .A2(new_n793), .A3(new_n796), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n794), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n771), .A2(new_n688), .A3(new_n772), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n799), .A2(KEYINPUT118), .B1(G106gat), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  OAI221_X1 g603(.A(new_n792), .B1(new_n797), .B2(new_n798), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n798), .A2(new_n797), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n800), .B2(new_n802), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT120), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1339gat));
  OR2_X1    g608(.A1(new_n668), .A2(new_n590), .ZN(new_n810));
  INV_X1    g609(.A(new_n648), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n578), .A2(new_n579), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n572), .A2(new_n573), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n586), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n588), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n752), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n663), .B1(new_n656), .B2(KEYINPUT54), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n652), .A2(new_n654), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n657), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n656), .A2(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n821), .A2(KEYINPUT55), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n664), .B1(new_n821), .B2(KEYINPUT55), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n816), .B1(new_n824), .B2(new_n590), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n706), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n706), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n815), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n811), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n810), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n688), .A3(new_n683), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n696), .A2(new_n488), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(G113gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(new_n834), .A3(new_n591), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n810), .A2(new_n829), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n836), .A2(new_n480), .A3(new_n832), .ZN(new_n837));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n590), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n835), .A2(new_n838), .ZN(G1340gat));
  OAI21_X1  g638(.A(G120gat), .B1(new_n833), .B2(new_n752), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT121), .Z(new_n841));
  INV_X1    g640(.A(G120gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n842), .A3(new_n667), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n833), .B2(new_n811), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n637), .A3(new_n648), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  INV_X1    g646(.A(G134gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n837), .A2(new_n848), .A3(new_n706), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT56), .Z(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n833), .B2(new_n624), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1343gat));
  INV_X1    g651(.A(new_n816), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n823), .B(new_n590), .C1(new_n821), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n706), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n811), .B1(new_n828), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n810), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT57), .A3(new_n688), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n836), .A2(new_n735), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n859), .B1(new_n861), .B2(KEYINPUT57), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n523), .A2(new_n832), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n590), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n321), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT58), .B1(new_n866), .B2(KEYINPUT123), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(new_n863), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(G141gat), .A3(new_n591), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n867), .B(new_n870), .ZN(G1344gat));
  INV_X1    g670(.A(new_n868), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n311), .A3(new_n667), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT124), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n862), .A2(new_n863), .ZN(new_n875));
  AOI211_X1 g674(.A(KEYINPUT59), .B(new_n311), .C1(new_n875), .C2(new_n667), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n827), .A2(KEYINPUT125), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n815), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n827), .A2(KEYINPUT125), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n856), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n810), .B1(new_n881), .B2(new_n648), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n687), .A2(KEYINPUT57), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n860), .A2(KEYINPUT57), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n667), .A3(new_n863), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n877), .B1(new_n885), .B2(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n874), .B1(new_n876), .B2(new_n886), .ZN(G1345gat));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n315), .A3(new_n648), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n875), .A2(new_n648), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n315), .ZN(G1346gat));
  AOI21_X1  g689(.A(G162gat), .B1(new_n872), .B2(new_n706), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n624), .A2(new_n316), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n875), .B2(new_n892), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n674), .A2(new_n677), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n831), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n204), .A3(new_n591), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n836), .A2(new_n480), .A3(new_n894), .ZN(new_n897));
  AOI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n590), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n896), .A2(new_n898), .ZN(G1348gat));
  OAI21_X1  g698(.A(G176gat), .B1(new_n895), .B2(new_n752), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n205), .A3(new_n667), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1349gat));
  OAI22_X1  g701(.A1(new_n895), .A2(new_n811), .B1(new_n220), .B2(new_n219), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n233), .A3(new_n648), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n895), .B2(new_n624), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT61), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n897), .A2(new_n228), .A3(new_n706), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1351gat));
  AND2_X1   g709(.A1(new_n523), .A2(new_n894), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n861), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n590), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n884), .A2(new_n911), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n591), .A2(new_n363), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1352gat));
  NAND3_X1  g716(.A1(new_n912), .A2(new_n364), .A3(new_n667), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G204gat), .B1(new_n914), .B2(new_n752), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n921), .B(new_n922), .C1(KEYINPUT62), .C2(new_n918), .ZN(G1353gat));
  INV_X1    g722(.A(G211gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n912), .A2(new_n924), .A3(new_n648), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n915), .A2(new_n648), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n926), .B2(G211gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1354gat));
  AOI21_X1  g728(.A(G218gat), .B1(new_n912), .B2(new_n706), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n706), .A2(G218gat), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT127), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n915), .B2(new_n932), .ZN(G1355gat));
endmodule


