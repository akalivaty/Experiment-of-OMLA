//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT68), .A3(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n190), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n200), .B2(new_n193), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n193), .B1(new_n189), .B2(new_n191), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT2), .B(G113), .Z(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G104), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(G107), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n209), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n208), .A2(G107), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n206), .A2(new_n207), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n196), .A2(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n221));
  INV_X1    g035(.A(new_n219), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT81), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n203), .A2(new_n204), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n203), .A2(KEYINPUT5), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n201), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n220), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G110), .B(G122), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT8), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n229), .A2(KEYINPUT82), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT82), .B1(new_n229), .B2(new_n231), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n222), .A2(new_n202), .A3(new_n205), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n209), .A2(new_n212), .A3(new_n214), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G101), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n203), .A2(new_n204), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n224), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n234), .B(new_n230), .C1(new_n239), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G125), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G143), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT66), .A3(new_n249), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT65), .B1(new_n245), .B2(G143), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n247), .A3(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n246), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT0), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT64), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(KEYINPUT0), .B2(G128), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n249), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n244), .B1(new_n255), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n253), .A2(new_n269), .A3(G128), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n256), .A2(new_n258), .B1(G143), .B2(new_n245), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n262), .B1(new_n246), .B2(KEYINPUT1), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n270), .B(new_n244), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G224), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(G953), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT7), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n268), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n263), .A2(new_n265), .ZN(new_n281));
  INV_X1    g095(.A(new_n249), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n252), .B(new_n254), .C1(new_n283), .C2(new_n271), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G125), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n278), .B1(new_n285), .B2(new_n273), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n243), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n232), .A2(new_n233), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT83), .B1(new_n288), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n233), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n229), .A2(KEYINPUT82), .A3(new_n231), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n234), .B1(new_n239), .B2(new_n242), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n285), .A2(new_n273), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n279), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n285), .A2(new_n273), .A3(new_n278), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n293), .A2(new_n230), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n230), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n292), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT6), .A3(new_n243), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n294), .A2(new_n276), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n285), .A2(new_n273), .A3(new_n277), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT6), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n292), .A2(new_n308), .A3(new_n302), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT80), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n304), .A2(new_n307), .A3(new_n312), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n289), .A2(new_n301), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G210), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n289), .A2(new_n314), .A3(new_n301), .A4(new_n316), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G214), .B1(G237), .B2(G902), .ZN(new_n321));
  INV_X1    g135(.A(G221), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT9), .B(G234), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(new_n324), .B2(new_n300), .ZN(new_n325));
  INV_X1    g139(.A(G469), .ZN(new_n326));
  AND4_X1   g140(.A1(new_n269), .A2(new_n246), .A3(new_n248), .A4(G128), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n328), .A2(G128), .B1(new_n246), .B2(new_n248), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n215), .B(new_n218), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(new_n222), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT11), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT67), .ZN(new_n334));
  INV_X1    g148(.A(G134), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G137), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(KEYINPUT67), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n339));
  INV_X1    g153(.A(G137), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT11), .A4(G134), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(G137), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G131), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(KEYINPUT11), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n339), .A2(KEYINPUT11), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n340), .A2(G134), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G131), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n342), .A4(new_n341), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n332), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT12), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  INV_X1    g168(.A(G953), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(G227), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n354), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n241), .A2(new_n255), .A3(new_n237), .A4(new_n267), .ZN(new_n359));
  INV_X1    g173(.A(new_n351), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n222), .A2(new_n331), .A3(KEYINPUT10), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n330), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT12), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n332), .A2(new_n365), .A3(new_n351), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n353), .A2(new_n358), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n359), .A2(new_n361), .A3(new_n363), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n351), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n358), .B1(new_n369), .B2(new_n364), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI211_X1 g186(.A(KEYINPUT78), .B(new_n358), .C1(new_n369), .C2(new_n364), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n326), .B(new_n300), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n353), .A2(new_n364), .A3(new_n366), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n357), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n369), .A2(new_n358), .A3(new_n364), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(G469), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(G469), .A2(G902), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n325), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n320), .A2(new_n321), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n272), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n327), .B1(new_n260), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n349), .B1(new_n347), .B2(new_n342), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n350), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n385), .B1(new_n388), .B2(KEYINPUT69), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT69), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n350), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  INV_X1    g205(.A(new_n284), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n389), .A2(new_n391), .B1(new_n392), .B2(new_n351), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n224), .A2(new_n238), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT70), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n338), .A2(new_n343), .A3(G131), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT69), .B1(new_n396), .B2(new_n386), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n331), .A3(new_n391), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n351), .A2(new_n267), .A3(new_n255), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(KEYINPUT70), .A3(new_n394), .A4(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n394), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n398), .B2(new_n399), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n331), .A2(new_n350), .A3(new_n387), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n399), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n403), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(G237), .A2(G953), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G210), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT27), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G101), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n398), .A2(new_n394), .A3(new_n399), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT70), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n399), .A2(new_n406), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n403), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n422), .A3(new_n400), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT28), .B1(new_n393), .B2(new_n394), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n416), .B(new_n417), .C1(new_n428), .C2(new_n415), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n420), .B(new_n400), .C1(new_n394), .C2(new_n393), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n430), .B2(KEYINPUT28), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n415), .A2(new_n417), .ZN(new_n432));
  AOI21_X1  g246(.A(G902), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G472), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT32), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n428), .A2(new_n415), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n408), .A2(new_n414), .A3(new_n420), .A4(new_n400), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT31), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n402), .A2(KEYINPUT31), .A3(new_n414), .A4(new_n408), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G472), .A2(G902), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n436), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  AOI211_X1 g260(.A(KEYINPUT32), .B(new_n446), .C1(new_n437), .C2(new_n442), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n435), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G217), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(G234), .B2(new_n300), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT72), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT72), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT23), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n452), .A2(new_n454), .B1(new_n188), .B2(G128), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT73), .B1(new_n188), .B2(G128), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n262), .A3(G119), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n262), .A2(G119), .ZN(new_n460));
  OAI22_X1  g274(.A1(new_n455), .A2(new_n459), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G119), .B(G128), .ZN(new_n462));
  XOR2_X1   g276(.A(KEYINPUT24), .B(G110), .Z(new_n463));
  OAI22_X1  g277(.A1(new_n461), .A2(G110), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT75), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n244), .A3(G140), .ZN(new_n466));
  INV_X1    g280(.A(G140), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n244), .A2(G140), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(KEYINPUT16), .B(new_n466), .C1(new_n470), .C2(new_n465), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT16), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G146), .ZN(new_n475));
  XNOR2_X1  g289(.A(G125), .B(G140), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n245), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n464), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT74), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n461), .A2(new_n479), .A3(G110), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n461), .B2(G110), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n463), .A2(new_n462), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n471), .A2(new_n245), .A3(new_n473), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n245), .B1(new_n471), .B2(new_n473), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n478), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT76), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT76), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n478), .C1(new_n482), .C2(new_n486), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT22), .B(G137), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n355), .A2(G221), .A3(G234), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n493), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(KEYINPUT76), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT25), .B1(new_n497), .B2(new_n300), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n499), .B(G902), .C1(new_n494), .C2(new_n496), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n450), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n450), .A2(G902), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT77), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(G475), .A2(G902), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n471), .A2(new_n245), .A3(new_n473), .ZN(new_n507));
  INV_X1    g321(.A(G237), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n355), .A3(G214), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n247), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n410), .A2(G143), .A3(G214), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT17), .A3(G131), .ZN(new_n513));
  INV_X1    g327(.A(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(G143), .B1(new_n410), .B2(G214), .ZN(new_n515));
  OAI21_X1  g329(.A(G131), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n349), .A3(new_n511), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n475), .A2(new_n507), .A3(new_n513), .A4(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G113), .B(G122), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(new_n208), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n476), .A2(KEYINPUT75), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n466), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n477), .B1(new_n524), .B2(new_n245), .ZN(new_n525));
  AND2_X1   g339(.A1(KEYINPUT18), .A2(G131), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n512), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n512), .A2(new_n526), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n520), .A2(new_n522), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n474), .A2(G146), .B1(new_n516), .B2(new_n518), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT19), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n523), .B2(new_n466), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n476), .A2(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n245), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n522), .B1(new_n536), .B2(new_n529), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n506), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT20), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n520), .A2(new_n522), .A3(new_n529), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n527), .A2(new_n528), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n525), .A2(new_n541), .B1(new_n531), .B2(new_n535), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n542), .B2(new_n522), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n506), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n520), .A2(new_n529), .ZN(new_n547));
  INV_X1    g361(.A(new_n522), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(KEYINPUT85), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT85), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n540), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n522), .B1(new_n520), .B2(new_n529), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n300), .B(new_n549), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT84), .B(G475), .Z(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n262), .A2(G143), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT13), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n335), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G128), .B(G143), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT86), .B1(new_n190), .B2(G122), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT86), .ZN(new_n564));
  INV_X1    g378(.A(G122), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(G116), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n190), .A2(G122), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n211), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n211), .B1(new_n567), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n568), .B(KEYINPUT14), .ZN(new_n573));
  INV_X1    g387(.A(new_n567), .ZN(new_n574));
  OAI21_X1  g388(.A(G107), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n561), .B(new_n335), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n323), .A2(new_n449), .A3(G953), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n572), .B2(new_n577), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n300), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G478), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT15), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI221_X1 g399(.A(new_n300), .B1(KEYINPUT15), .B2(new_n583), .C1(new_n580), .C2(new_n581), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G952), .ZN(new_n588));
  AOI211_X1 g402(.A(G953), .B(new_n588), .C1(G234), .C2(G237), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n300), .B(new_n355), .C1(G234), .C2(G237), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT21), .B(G898), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n557), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n383), .A2(new_n448), .A3(new_n505), .A4(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  OAI21_X1  g409(.A(KEYINPUT33), .B1(new_n580), .B2(new_n581), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n572), .A2(new_n577), .ZN(new_n597));
  INV_X1    g411(.A(new_n578), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n579), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n583), .A2(G902), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT89), .B(G478), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n602), .A2(new_n603), .B1(new_n582), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n557), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n592), .ZN(new_n609));
  INV_X1    g423(.A(new_n321), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n318), .B2(new_n319), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(KEYINPUT88), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT88), .ZN(new_n613));
  AOI211_X1 g427(.A(new_n613), .B(new_n610), .C1(new_n318), .C2(new_n319), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n609), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n443), .B(new_n300), .C1(KEYINPUT87), .C2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(KEYINPUT87), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n415), .A2(new_n428), .B1(new_n440), .B2(new_n441), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(G902), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n381), .A2(new_n501), .A3(new_n504), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n320), .A2(new_n321), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n613), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n611), .A2(KEYINPUT88), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT91), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n556), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n553), .A2(KEYINPUT91), .A3(new_n555), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n539), .A2(KEYINPUT90), .A3(new_n545), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT90), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n538), .A2(new_n637), .A3(KEYINPUT20), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n587), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n635), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n592), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n641), .A2(KEYINPUT92), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT92), .B1(new_n641), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n631), .A2(new_n623), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NOR2_X1   g462(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT94), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT93), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(new_n487), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n487), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n503), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n501), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n593), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n621), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n383), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n589), .B1(new_n590), .B2(new_n661), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n635), .A2(new_n639), .A3(new_n640), .A4(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n663), .A2(new_n381), .A3(new_n655), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(new_n448), .C1(new_n612), .C2(new_n614), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  XOR2_X1   g480(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n320), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n557), .A2(new_n587), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n668), .A2(new_n610), .A3(new_n655), .A4(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT96), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT32), .B1(new_n619), .B2(new_n446), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n440), .A2(new_n441), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n414), .B1(new_n425), .B2(new_n427), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n436), .B(new_n444), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(G902), .B1(new_n409), .B2(new_n414), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n430), .A2(new_n414), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n616), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n671), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  AOI211_X1 g495(.A(KEYINPUT96), .B(new_n679), .C1(new_n672), .C2(new_n675), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n670), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n662), .B(KEYINPUT39), .Z(new_n686));
  AND2_X1   g500(.A1(new_n381), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT97), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n247), .ZN(G45));
  NOR2_X1   g506(.A1(new_n608), .A2(new_n662), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n655), .A2(new_n381), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n695), .B(new_n448), .C1(new_n612), .C2(new_n614), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  AOI22_X1  g511(.A1(new_n672), .A2(new_n675), .B1(G472), .B2(new_n434), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n501), .A2(new_n504), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n300), .B1(new_n372), .B2(new_n373), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  INV_X1    g516(.A(new_n325), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n374), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT98), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n702), .A2(KEYINPUT98), .A3(new_n703), .A4(new_n374), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n631), .A2(new_n700), .A3(new_n609), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n631), .A2(new_n700), .A3(new_n645), .A4(new_n708), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT99), .B(G116), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G18));
  NOR2_X1   g528(.A1(new_n698), .A2(new_n656), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n631), .A2(new_n708), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  XNOR2_X1  g531(.A(new_n669), .B(KEYINPUT100), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n431), .A2(new_n414), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n444), .B1(new_n673), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n619), .B2(G902), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n505), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n706), .A2(new_n642), .A3(new_n707), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n631), .A2(new_n719), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  AND4_X1   g541(.A1(new_n655), .A2(new_n722), .A3(new_n693), .A4(new_n721), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(new_n708), .C1(new_n612), .C2(new_n614), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  NAND3_X1  g544(.A1(new_n318), .A2(new_n321), .A3(new_n319), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n375), .A2(KEYINPUT101), .A3(new_n357), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT101), .B1(new_n375), .B2(new_n357), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n377), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n374), .B(new_n379), .C1(new_n734), .C2(new_n326), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n703), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n448), .A2(new_n737), .A3(new_n505), .A4(new_n693), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(KEYINPUT102), .A3(KEYINPUT42), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT42), .B1(new_n738), .B2(KEYINPUT102), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NAND4_X1  g556(.A1(new_n448), .A2(new_n737), .A3(new_n505), .A4(new_n663), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n734), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n376), .A2(new_n377), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n326), .B1(new_n747), .B2(new_n745), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n379), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n750), .A2(KEYINPUT46), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(KEYINPUT103), .A3(KEYINPUT46), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n379), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n751), .A2(new_n374), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n703), .A3(new_n686), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n731), .ZN(new_n760));
  INV_X1    g574(.A(new_n557), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT43), .A3(new_n607), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n606), .A2(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n606), .A2(KEYINPUT105), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n765), .A2(KEYINPUT106), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT106), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n621), .A3(new_n655), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n760), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n759), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  AND4_X1   g589(.A1(new_n699), .A2(new_n698), .A3(new_n693), .A4(new_n760), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT108), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n756), .A2(new_n703), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n756), .A2(new_n703), .B1(KEYINPUT107), .B2(new_n781), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n777), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT109), .B(G140), .Z(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G42));
  NAND3_X1  g599(.A1(new_n607), .A2(new_n321), .A3(new_n703), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n699), .A2(new_n557), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n702), .A2(new_n374), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT110), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n789), .B2(KEYINPUT49), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(KEYINPUT49), .B2(new_n789), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n683), .A3(new_n668), .ZN(new_n792));
  INV_X1    g606(.A(new_n723), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n769), .A2(new_n589), .A3(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n780), .A2(new_n782), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n789), .A2(new_n703), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n731), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n708), .A2(new_n589), .A3(new_n760), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n683), .A2(new_n505), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n557), .A3(new_n607), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n668), .A2(new_n610), .A3(new_n708), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n794), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n802), .A2(new_n804), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n798), .A2(new_n769), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n722), .A2(new_n655), .A3(new_n721), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OR4_X1    g624(.A1(new_n800), .A2(new_n806), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n797), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT51), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT115), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n736), .A2(new_n655), .A3(new_n662), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n681), .B2(new_n682), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n719), .B1(new_n612), .B2(new_n614), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n729), .A2(new_n665), .A3(new_n696), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n718), .B1(new_n629), .B2(new_n630), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n823), .B(new_n817), .C1(new_n682), .C2(new_n681), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n631), .B(new_n448), .C1(new_n664), .C2(new_n695), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(KEYINPUT52), .A3(new_n729), .A4(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n621), .ZN(new_n828));
  INV_X1    g642(.A(new_n608), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n610), .B(new_n592), .C1(new_n318), .C2(new_n319), .ZN(new_n830));
  INV_X1    g644(.A(new_n622), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n594), .A2(new_n832), .A3(new_n658), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n448), .A2(new_n708), .A3(new_n505), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n615), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n298), .A2(new_n300), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n837), .A2(KEYINPUT83), .B1(new_n311), .B2(new_n313), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n316), .B1(new_n838), .B2(new_n301), .ZN(new_n839));
  INV_X1    g653(.A(new_n319), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n321), .B(new_n642), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n557), .A2(new_n640), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n836), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n611), .A2(KEYINPUT111), .A3(new_n642), .A4(new_n842), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n844), .A2(new_n623), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n833), .A2(new_n835), .A3(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n712), .A2(new_n716), .A3(new_n726), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n728), .A2(new_n737), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n743), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n662), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n585), .A2(new_n586), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n636), .A2(new_n852), .A3(new_n638), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n635), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n450), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n490), .A2(new_n493), .ZN(new_n856));
  OAI221_X1 g670(.A(new_n483), .B1(new_n484), .B2(new_n485), .C1(new_n480), .C2(new_n481), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n489), .B1(new_n857), .B2(new_n478), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n496), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n300), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n499), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n497), .A2(KEYINPUT25), .A3(new_n300), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n855), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n654), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n854), .B(new_n381), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n448), .A2(new_n867), .A3(new_n868), .A4(new_n760), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n448), .A2(new_n867), .A3(new_n760), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT112), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n850), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n847), .A2(new_n848), .A3(new_n741), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n827), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n738), .A2(KEYINPUT102), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT42), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n871), .A2(new_n869), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n738), .A2(KEYINPUT102), .A3(KEYINPUT42), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n743), .A2(new_n849), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n712), .A2(new_n716), .A3(new_n726), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n621), .A2(new_n608), .A3(new_n622), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n884), .A2(new_n830), .B1(new_n657), .B2(new_n383), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n844), .A2(new_n623), .A3(new_n845), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n709), .A2(new_n885), .A3(new_n594), .A4(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n882), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n822), .A2(new_n826), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n815), .B1(new_n875), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n874), .B1(new_n827), .B2(new_n873), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(KEYINPUT53), .A3(new_n889), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(KEYINPUT54), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n794), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n631), .A3(new_n708), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n897), .A2(G952), .A3(new_n355), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n798), .A2(new_n700), .A3(new_n769), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT48), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n898), .B(new_n900), .C1(new_n608), .C2(new_n799), .ZN(new_n901));
  INV_X1    g715(.A(new_n812), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n814), .A2(new_n895), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n792), .B1(new_n905), .B2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n355), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n892), .A2(new_n893), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n300), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT56), .B1(new_n912), .B2(G210), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n304), .A2(new_n309), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n307), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT55), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n909), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT116), .B1(new_n910), .B2(G902), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n919), .B(new_n300), .C1(new_n892), .C2(new_n893), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n317), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n916), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n922), .B2(new_n924), .ZN(G51));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n379), .B(KEYINPUT57), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n891), .A2(new_n894), .A3(new_n927), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n372), .A2(new_n373), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n928), .A2(KEYINPUT117), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT117), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n918), .A2(new_n920), .A3(new_n749), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n926), .B1(new_n933), .B2(new_n908), .ZN(new_n934));
  INV_X1    g748(.A(new_n932), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n928), .A2(new_n929), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(KEYINPUT118), .B(new_n909), .C1(new_n939), .C2(new_n930), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n934), .A2(new_n940), .ZN(G54));
  NAND3_X1  g755(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n942), .B(new_n540), .C1(new_n522), .C2(new_n542), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .A4(new_n543), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n943), .A2(new_n909), .A3(new_n944), .ZN(G60));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT59), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n891), .A2(new_n894), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n602), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n908), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n911), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n955), .A2(new_n652), .A3(new_n653), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n909), .B1(new_n955), .B2(new_n497), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n958));
  OAI22_X1  g772(.A1(new_n956), .A2(new_n957), .B1(KEYINPUT119), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT119), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G66));
  NOR3_X1   g775(.A1(new_n591), .A2(new_n275), .A3(new_n355), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n887), .A2(new_n883), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n355), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n914), .B1(G898), .B2(new_n355), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(G69));
  AOI21_X1  g780(.A(new_n355), .B1(G227), .B2(G900), .ZN(new_n967));
  INV_X1    g781(.A(new_n821), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n783), .A2(new_n968), .A3(new_n743), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n774), .A2(new_n741), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n759), .A2(new_n700), .A3(new_n823), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n741), .A3(new_n774), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT126), .B1(new_n975), .B2(new_n969), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n355), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n533), .A2(new_n534), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT120), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT121), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n405), .A2(new_n407), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(new_n982));
  NAND2_X1  g796(.A1(G900), .A2(G953), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n977), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n691), .A2(KEYINPUT62), .A3(new_n821), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT122), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n843), .A2(new_n608), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT123), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n700), .A2(new_n988), .A3(new_n687), .A4(new_n760), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n774), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n774), .A2(new_n992), .A3(new_n989), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT62), .B1(new_n691), .B2(new_n821), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n783), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n986), .A2(new_n991), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n982), .B1(new_n996), .B2(new_n355), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n984), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n967), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n997), .A2(new_n998), .ZN(new_n1003));
  INV_X1    g817(.A(new_n967), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1003), .A2(new_n1004), .A3(new_n1000), .A4(new_n984), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(new_n409), .A2(new_n414), .ZN(new_n1007));
  OR3_X1    g821(.A1(new_n996), .A2(new_n883), .A3(new_n887), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT63), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT127), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1007), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n974), .A2(new_n963), .A3(new_n976), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n414), .B(new_n409), .C1(new_n1013), .C2(new_n1011), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n1010), .B(new_n911), .C1(new_n438), .C2(new_n416), .ZN(new_n1015));
  NOR4_X1   g829(.A1(new_n1012), .A2(new_n1014), .A3(new_n908), .A4(new_n1015), .ZN(G57));
endmodule


