//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(G125), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n464), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n466), .A2(G137), .A3(new_n468), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n468), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n470), .A2(new_n471), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(new_n468), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n468), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT70), .Z(G162));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n470), .B2(new_n471), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n470), .B2(new_n471), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n502), .B(new_n505), .C1(new_n471), .C2(new_n470), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n500), .B1(new_n504), .B2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n517), .B1(new_n514), .B2(KEYINPUT5), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n512), .A2(KEYINPUT72), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n516), .A2(new_n520), .A3(G88), .A4(new_n508), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n510), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n516), .A2(new_n520), .A3(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT73), .Z(new_n526));
  AOI21_X1  g101(.A(new_n523), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n516), .A2(new_n520), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n516), .A2(new_n520), .A3(KEYINPUT74), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n531), .A2(G63), .A3(G651), .A4(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n516), .A2(new_n520), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G89), .A3(new_n508), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n509), .A2(G51), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  AND2_X1   g116(.A1(new_n534), .A2(new_n508), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G90), .B1(G52), .B2(new_n509), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n516), .A2(new_n520), .A3(KEYINPUT74), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT74), .B1(new_n516), .B2(new_n520), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n546), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n543), .B1(new_n547), .B2(new_n523), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n509), .A2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n534), .A2(new_n508), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n531), .A2(G56), .A3(new_n532), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g132(.A(KEYINPUT75), .B(new_n554), .C1(new_n557), .C2(new_n523), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n523), .B1(new_n555), .B2(new_n556), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(new_n553), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND4_X1  g143(.A1(new_n516), .A2(new_n520), .A3(G91), .A4(new_n508), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n516), .A2(new_n520), .A3(G65), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n508), .A2(G53), .A3(G543), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n570), .A2(new_n574), .A3(new_n576), .A4(new_n577), .ZN(G299));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n509), .A2(G49), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n516), .A2(new_n520), .A3(G87), .A4(new_n508), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n544), .B2(new_n545), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n582), .B1(new_n584), .B2(G651), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n509), .A2(G48), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n516), .A2(new_n520), .A3(G86), .A4(new_n508), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n516), .A2(new_n520), .A3(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT77), .Z(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n591), .B1(new_n595), .B2(G651), .ZN(new_n596));
  AOI211_X1 g171(.A(KEYINPUT78), .B(new_n523), .C1(new_n592), .C2(new_n594), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n546), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n523), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n509), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n551), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n529), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n516), .A2(new_n520), .A3(G92), .A4(new_n508), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G171), .B2(new_n614), .ZN(G284));
  OAI21_X1  g191(.A(new_n615), .B1(G171), .B2(new_n614), .ZN(G321));
  NOR2_X1   g192(.A1(G286), .A2(new_n614), .ZN(new_n618));
  XNOR2_X1  g193(.A(G299), .B(KEYINPUT79), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n614), .ZN(G297));
  AOI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n614), .ZN(G280));
  AND2_X1   g196(.A1(new_n609), .A2(new_n612), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT80), .Z(G148));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n563), .B2(G868), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n466), .A2(new_n478), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT81), .B(G2100), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n484), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n486), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n468), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n635), .A3(new_n641), .ZN(G156));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2430), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT82), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n654), .ZN(G401));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2096), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  AND2_X1   g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT84), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n672), .A2(new_n679), .A3(new_n675), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1981), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(KEYINPUT103), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G26), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT28), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n484), .A2(G140), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n486), .A2(G128), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n468), .A2(G116), .ZN(new_n696));
  OAI21_X1  g271(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n694), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n693), .B1(new_n702), .B2(G29), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT94), .ZN(new_n704));
  INV_X1    g279(.A(G2067), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G19), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n563), .B2(new_n707), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1341), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(G20), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT23), .ZN(new_n712));
  AND4_X1   g287(.A1(new_n576), .A2(new_n570), .A3(new_n574), .A4(new_n577), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n707), .ZN(new_n714));
  INV_X1    g289(.A(G1956), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n691), .A2(G35), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G162), .B2(new_n691), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT29), .B(G2090), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n622), .A2(G16), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G4), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT92), .B(G1348), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n720), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AND4_X1   g301(.A1(new_n706), .A2(new_n710), .A3(new_n716), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT102), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT26), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G129), .B2(new_n486), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n478), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT96), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G29), .B2(G32), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT97), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT97), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n736), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G33), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n466), .A2(G127), .ZN(new_n746));
  NAND2_X1  g321(.A1(G115), .A2(G2104), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n468), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n745), .B(new_n748), .C1(G139), .C2(new_n484), .ZN(new_n749));
  MUX2_X1   g324(.A(new_n743), .B(new_n749), .S(G29), .Z(new_n750));
  INV_X1    g325(.A(G2072), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT31), .B(G11), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n691), .B1(new_n754), .B2(G28), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(KEYINPUT99), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(G28), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n755), .B2(KEYINPUT99), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n753), .B1(new_n756), .B2(new_n758), .C1(new_n640), .C2(new_n691), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n750), .B2(new_n751), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n752), .B(new_n760), .C1(new_n736), .C2(new_n737), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT24), .B(G34), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(new_n691), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT95), .Z(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n481), .B2(new_n691), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G16), .A2(G21), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G168), .B2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT98), .B(G1966), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n691), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n691), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT100), .B(G2078), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT101), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n742), .A2(new_n768), .A3(new_n772), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n707), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n707), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1961), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n728), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n778), .A2(KEYINPUT102), .A3(new_n782), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n690), .B(new_n727), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n727), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(KEYINPUT103), .ZN(new_n788));
  NOR2_X1   g363(.A1(G25), .A2(G29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n484), .A2(G131), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n486), .A2(G119), .ZN(new_n791));
  OR2_X1    g366(.A1(G95), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(G29), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT35), .B(G1991), .Z(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT85), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n604), .A2(G16), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G16), .B2(G24), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT86), .B(G1986), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT87), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G305), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n707), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G6), .B2(new_n707), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT32), .B(G1981), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n707), .A2(G23), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n585), .B2(new_n707), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT33), .B(G1976), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n707), .A2(G22), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT89), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G166), .B2(new_n707), .ZN(new_n820));
  INV_X1    g395(.A(G1971), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n809), .A2(new_n811), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n817), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n817), .A2(new_n827), .A3(new_n824), .A4(new_n825), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n803), .A2(KEYINPUT87), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n806), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(KEYINPUT91), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n833), .A2(KEYINPUT91), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n786), .A2(new_n788), .B1(new_n835), .B2(new_n836), .ZN(G311));
  NAND2_X1  g412(.A1(new_n788), .A2(new_n786), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n836), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(G150));
  NAND2_X1  g415(.A1(new_n542), .A2(G93), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n509), .A2(G55), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n546), .A2(G67), .ZN(new_n844));
  INV_X1    g419(.A(G80), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n845), .B2(new_n514), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n843), .B1(new_n846), .B2(G651), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT105), .B(G860), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n546), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n842), .B(new_n841), .C1(new_n851), .C2(new_n523), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n562), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n554), .B1(new_n557), .B2(new_n523), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n613), .A2(new_n623), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT106), .Z(new_n863));
  OAI21_X1  g438(.A(new_n848), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n850), .B1(new_n863), .B2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n481), .B(new_n640), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(G162), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n504), .A2(new_n506), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n492), .B1(new_n494), .B2(G2105), .ZN(new_n870));
  OR2_X1    g445(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n871));
  NAND2_X1  g446(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n497), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n496), .A2(new_n499), .A3(KEYINPUT107), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n702), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n795), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n486), .A2(G130), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n468), .A2(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(G142), .B2(new_n484), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT108), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n631), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n878), .A2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n749), .A2(new_n733), .ZN(new_n888));
  INV_X1    g463(.A(new_n734), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(new_n749), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n886), .B2(new_n887), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n867), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n878), .B(new_n885), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n890), .ZN(new_n898));
  INV_X1    g473(.A(new_n867), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n892), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(new_n852), .A2(new_n614), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n622), .A2(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n713), .A2(new_n613), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT41), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n905), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n626), .B(KEYINPUT109), .Z(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(new_n857), .ZN(new_n912));
  MUX2_X1   g487(.A(new_n909), .B(new_n910), .S(new_n912), .Z(new_n913));
  NAND2_X1  g488(.A1(G290), .A2(new_n807), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n604), .A2(G305), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G303), .B(new_n585), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT42), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n913), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n903), .B1(new_n920), .B2(new_n614), .ZN(G295));
  OAI21_X1  g496(.A(new_n903), .B1(new_n920), .B2(new_n614), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  XNOR2_X1  g498(.A(G301), .B(G168), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n847), .B1(new_n561), .B2(new_n558), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n855), .ZN(new_n926));
  XNOR2_X1  g501(.A(G301), .B(G286), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n853), .A3(new_n856), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n910), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n906), .A2(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n906), .A2(KEYINPUT110), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n908), .A3(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(KEYINPUT111), .A3(new_n928), .A4(new_n926), .ZN(new_n936));
  INV_X1    g511(.A(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n908), .B1(new_n906), .B2(KEYINPUT110), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n926), .B(new_n928), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n904), .A2(new_n905), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n926), .B2(new_n928), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT112), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n932), .A2(new_n936), .A3(new_n941), .A4(new_n944), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n916), .B(new_n917), .Z(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n926), .A2(new_n909), .A3(new_n928), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n918), .A2(new_n930), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n950), .A2(new_n896), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n930), .A2(new_n949), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n946), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n948), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n923), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n941), .A2(new_n936), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n943), .B(new_n931), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n918), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n950), .A2(new_n896), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT43), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n955), .A2(new_n948), .A3(new_n896), .A4(new_n950), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT113), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n948), .B1(new_n947), .B2(new_n951), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n957), .B1(new_n965), .B2(new_n969), .ZN(G397));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n876), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT114), .B(KEYINPUT45), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n477), .A2(G40), .A3(new_n479), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n474), .B1(new_n473), .B2(G2105), .ZN(new_n977));
  AOI211_X1 g552(.A(KEYINPUT69), .B(new_n468), .C1(new_n472), .C2(new_n464), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n702), .A2(G2067), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n700), .A2(new_n705), .A3(new_n701), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n983), .B2(new_n733), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT126), .Z(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  INV_X1    g565(.A(new_n983), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n733), .A2(G1996), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n991), .B(new_n992), .C1(G1996), .C2(new_n889), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n794), .B(new_n797), .Z(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n980), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OR3_X1    g572(.A1(G290), .A2(new_n996), .A3(G1986), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(KEYINPUT48), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(KEYINPUT48), .B2(new_n999), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n795), .A2(new_n797), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n982), .B1(new_n993), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n980), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n990), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT60), .ZN(new_n1006));
  INV_X1    g581(.A(new_n723), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n466), .A2(new_n498), .B1(new_n493), .B2(new_n495), .ZN(new_n1009));
  INV_X1    g584(.A(new_n506), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n505), .B1(new_n466), .B2(new_n502), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1008), .B1(new_n1012), .B2(new_n971), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(new_n979), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n876), .A2(new_n1008), .A3(new_n971), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1007), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n972), .A2(new_n979), .A3(G2067), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1006), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n477), .A2(G40), .A3(new_n479), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n469), .B2(new_n475), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1015), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n723), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1017), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT60), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1025), .A3(new_n622), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n974), .B1(G164), .B2(G1384), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n986), .A4(new_n1021), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT58), .B(G1341), .Z(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n972), .B2(new_n979), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT119), .B(new_n1027), .C1(new_n1034), .C2(new_n562), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT60), .A3(new_n613), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1026), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n972), .A2(KEYINPUT50), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1012), .A2(new_n1008), .A3(new_n971), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT116), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1012), .A2(new_n1042), .A3(new_n1008), .A4(new_n971), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1039), .A2(new_n1041), .A3(new_n1021), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n715), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1028), .A2(new_n1029), .A3(new_n1021), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n523), .B1(new_n571), .B2(new_n572), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(new_n576), .C1(KEYINPUT117), .C2(KEYINPUT57), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT117), .A4(new_n577), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n1057));
  NAND3_X1  g632(.A1(G299), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(KEYINPUT118), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1050), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1044), .A2(new_n715), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n1059), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1045), .A2(new_n1059), .A3(new_n1049), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1059), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n563), .A2(new_n1071), .A3(new_n1033), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT119), .B1(new_n1034), .B2(new_n562), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(KEYINPUT59), .A3(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1038), .A2(new_n1067), .A3(new_n1070), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n622), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1068), .A2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(new_n1063), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1012), .A2(new_n971), .A3(new_n973), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1021), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT45), .B1(new_n876), .B2(new_n971), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT120), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n1086));
  NOR4_X1   g661(.A1(new_n1081), .A2(new_n1082), .A3(new_n1086), .A4(G2078), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT121), .B(G1961), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1022), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1028), .A2(new_n1029), .A3(new_n1084), .A4(new_n1021), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1092), .A2(KEYINPUT122), .A3(new_n1088), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT122), .B1(new_n1092), .B2(new_n1088), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(G171), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g671(.A(new_n1088), .B(G2078), .C1(new_n473), .C2(G2105), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n975), .A2(new_n976), .A3(new_n1028), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1092), .A2(new_n1088), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1092), .A2(KEYINPUT122), .A3(new_n1088), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1100), .A2(new_n1105), .A3(G301), .A4(new_n1091), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT54), .B1(new_n1096), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n522), .B2(new_n527), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n973), .B1(new_n1012), .B2(new_n971), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(new_n979), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1971), .B1(new_n1112), .B2(new_n1028), .ZN(new_n1113));
  INV_X1    g688(.A(G2090), .ZN(new_n1114));
  AND4_X1   g689(.A1(new_n1114), .A2(new_n1015), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1110), .B(G8), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G8), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n979), .B1(new_n972), .B2(KEYINPUT50), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(new_n1114), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1046), .A2(new_n821), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1116), .B1(new_n1121), .B2(new_n1110), .ZN(new_n1122));
  INV_X1    g697(.A(G1981), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(new_n590), .C1(new_n596), .C2(new_n597), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n523), .B1(new_n592), .B2(new_n594), .ZN(new_n1125));
  OAI21_X1  g700(.A(G1981), .B1(new_n589), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT49), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(KEYINPUT49), .A3(new_n1126), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n876), .A2(new_n971), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1117), .B1(new_n1131), .B2(new_n1021), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n585), .B2(G1976), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n585), .A2(G1976), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1976), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1138), .B(new_n582), .C1(new_n584), .C2(G651), .ZN(new_n1139));
  OAI21_X1  g714(.A(G8), .B1(new_n972), .B2(new_n979), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1134), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1133), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1122), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n771), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1015), .A2(new_n1019), .A3(new_n766), .A4(new_n1021), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(G168), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(G8), .ZN(new_n1148));
  AOI21_X1  g723(.A(G168), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT51), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(new_n1151), .A3(G8), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1144), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1107), .A2(new_n1154), .ZN(new_n1155));
  OR3_X1    g730(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1156), .A2(G301), .A3(new_n1105), .A4(new_n1091), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1098), .B(KEYINPUT123), .ZN(new_n1158));
  OAI21_X1  g733(.A(G171), .B1(new_n1095), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(KEYINPUT54), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1157), .A2(new_n1159), .A3(new_n1162), .A4(KEYINPUT54), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1079), .A2(new_n1155), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1166), .A2(G8), .A3(G168), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(KEYINPUT63), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1110), .B2(new_n1121), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1143), .B1(new_n1169), .B2(new_n1116), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1143), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1110), .ZN(new_n1173));
  OAI21_X1  g748(.A(G8), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1167), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1171), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1132), .B(KEYINPUT115), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1133), .A2(new_n1138), .A3(new_n585), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n1124), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1170), .A2(new_n1176), .A3(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1164), .A2(new_n1165), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1165), .B1(new_n1164), .B2(new_n1180), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1153), .A2(KEYINPUT62), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1096), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n1144), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1153), .A2(KEYINPUT62), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1181), .A2(new_n1182), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n604), .B(G1986), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n996), .B1(new_n995), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1005), .B1(new_n1188), .B2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g766(.A(new_n961), .B1(new_n954), .B2(new_n946), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n952), .B1(new_n948), .B2(new_n1193), .ZN(new_n1194));
  NOR3_X1   g768(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1195));
  XOR2_X1   g769(.A(new_n1195), .B(KEYINPUT127), .Z(new_n1196));
  NOR2_X1   g770(.A1(new_n1196), .A2(G229), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n1194), .A2(new_n901), .A3(new_n1197), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


