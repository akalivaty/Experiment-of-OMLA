//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1214, new_n1215,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT69), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n459), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n464));
  NAND4_X1  g039(.A1(new_n462), .A2(G137), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n459), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n461), .A2(new_n473), .A3(G125), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n461), .A2(new_n473), .A3(new_n476), .A4(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n469), .A2(new_n471), .B1(G2105), .B2(new_n478), .ZN(G160));
  AND2_X1   g054(.A1(new_n462), .A2(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  OR3_X1    g057(.A1(new_n481), .A2(KEYINPUT71), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n480), .A2(new_n463), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT71), .B1(new_n481), .B2(new_n482), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n483), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n490), .B(new_n491), .ZN(G162));
  NAND2_X1  g067(.A1(new_n461), .A2(new_n473), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n463), .A3(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n462), .A2(G138), .A3(new_n463), .A4(new_n464), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n462), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n498), .A2(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n504), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT74), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(new_n517), .A3(G651), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n507), .A2(new_n509), .B1(new_n506), .B2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G88), .B1(G50), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n516), .A2(new_n518), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  AND2_X1   g102(.A1(new_n522), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n528), .A2(new_n533), .ZN(G168));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n521), .A2(new_n535), .B1(new_n536), .B2(new_n523), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n519), .A2(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR3_X1    g116(.A1(new_n537), .A2(new_n541), .A3(KEYINPUT75), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT75), .B1(new_n537), .B2(new_n541), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G171));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n521), .A2(new_n545), .B1(new_n546), .B2(new_n523), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n550), .B2(new_n538), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n512), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n554), .A2(KEYINPUT76), .A3(G651), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n548), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n512), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n522), .A2(G91), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n523), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n520), .A2(new_n571), .A3(G53), .A4(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n567), .A2(new_n568), .A3(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  NAND2_X1  g151(.A1(new_n524), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n519), .A2(G87), .A3(new_n520), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n524), .A2(G48), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n538), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n519), .A2(G86), .A3(new_n520), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n512), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(KEYINPUT78), .A3(G651), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n522), .A2(G85), .B1(G47), .B2(new_n524), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n512), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n538), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g178(.A(KEYINPUT80), .B(new_n599), .C1(new_n512), .C2(new_n600), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n606));
  NAND3_X1  g181(.A1(new_n522), .A2(G92), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n606), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n521), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n524), .A2(G54), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n605), .A2(KEYINPUT81), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT81), .B1(new_n605), .B2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n598), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n598), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  XNOR2_X1  g194(.A(G299), .B(KEYINPUT82), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n556), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n615), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n625), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT83), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g205(.A(new_n481), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n485), .A2(G135), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n638), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT13), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2446), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n654), .A2(G2443), .ZN(new_n655));
  INV_X1    g230(.A(G2443), .ZN(new_n656));
  NAND4_X1  g231(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n656), .A4(new_n653), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n648), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(G2443), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n657), .A3(new_n647), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1341), .B(G1348), .Z(new_n663));
  AOI21_X1  g238(.A(KEYINPUT86), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n659), .A2(new_n665), .A3(new_n661), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G14), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(KEYINPUT86), .A3(new_n663), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  OR3_X1    g250(.A1(new_n674), .A2(KEYINPUT87), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(KEYINPUT87), .B1(new_n674), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n673), .B(KEYINPUT17), .Z(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n677), .C1(new_n671), .C2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n675), .A3(new_n671), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n672), .A2(new_n675), .A3(new_n673), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT18), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n690), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n689), .B(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n699), .A2(new_n695), .A3(new_n691), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n690), .B2(new_n694), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n699), .A2(KEYINPUT20), .A3(new_n693), .A4(new_n692), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n701), .A2(new_n702), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G1991), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n704), .A2(new_n705), .A3(new_n700), .A4(new_n697), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT88), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n707), .B1(new_n706), .B2(new_n709), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n688), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n712), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n714), .A2(G1996), .A3(new_n710), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1981), .B(G1986), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n717), .B1(new_n713), .B2(new_n715), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n687), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n713), .A2(new_n715), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(new_n716), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n723), .A2(new_n686), .A3(new_n718), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(G229));
  NAND2_X1  g300(.A1(G162), .A2(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G29), .B2(G35), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT29), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT100), .ZN(new_n729));
  INV_X1    g304(.A(G2090), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT89), .B(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G20), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G299), .B2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1956), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n485), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n466), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n631), .A2(KEYINPUT97), .A3(G129), .ZN(new_n746));
  AOI21_X1  g321(.A(KEYINPUT97), .B1(new_n631), .B2(G129), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n740), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G32), .B(new_n748), .S(G29), .Z(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  OAI21_X1  g325(.A(new_n739), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n636), .A2(G29), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT98), .Z(new_n753));
  NAND2_X1  g328(.A1(G168), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G16), .B2(G21), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT31), .B(G11), .Z(new_n759));
  INV_X1    g334(.A(G28), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT99), .B1(new_n760), .B2(KEYINPUT30), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(KEYINPUT30), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n760), .A2(KEYINPUT99), .A3(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n757), .A2(new_n758), .A3(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n751), .A2(new_n753), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G33), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n466), .A2(G103), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT95), .Z(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT25), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n485), .A2(G139), .ZN(new_n773));
  NAND2_X1  g348(.A1(G115), .A2(G2104), .ZN(new_n774));
  INV_X1    g349(.A(G127), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n493), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G2105), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n771), .A2(KEYINPUT25), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n772), .A2(new_n773), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n769), .B1(new_n780), .B2(new_n768), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G2072), .Z(new_n782));
  NOR2_X1   g357(.A1(G27), .A2(G29), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G164), .B2(G29), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G2078), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(G2078), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n749), .B2(new_n750), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n767), .A2(new_n782), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n789));
  INV_X1    g364(.A(G26), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G29), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(G29), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n480), .A2(G128), .A3(G2105), .ZN(new_n793));
  OR2_X1    g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n795));
  INV_X1    g370(.A(G140), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n793), .B(new_n795), .C1(new_n484), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n792), .B1(new_n797), .B2(G29), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n791), .B1(new_n798), .B2(new_n789), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(G2067), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT24), .B(G34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(new_n768), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT96), .ZN(new_n803));
  INV_X1    g378(.A(G160), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n768), .ZN(new_n805));
  INV_X1    g380(.A(G2084), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n799), .A2(G2067), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n800), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G5), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G171), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1961), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n734), .A2(G19), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n557), .B2(new_n734), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT94), .B(G1341), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  NOR4_X1   g392(.A1(new_n788), .A2(new_n810), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G16), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G4), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n616), .B2(new_n819), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT93), .B(G1348), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n728), .B2(new_n730), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n733), .A2(new_n818), .A3(new_n824), .ZN(new_n825));
  MUX2_X1   g400(.A(G290), .B(G24), .S(new_n734), .Z(new_n826));
  XOR2_X1   g401(.A(KEYINPUT90), .B(G1986), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n768), .A2(G25), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n631), .A2(G119), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n485), .A2(G131), .ZN(new_n831));
  OR2_X1    g406(.A1(G95), .A2(G2105), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n829), .B1(new_n835), .B2(new_n768), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT35), .B(G1991), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n819), .A2(G6), .ZN(new_n840));
  INV_X1    g415(.A(G305), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(new_n819), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT32), .B(G1981), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(G16), .A2(G23), .ZN(new_n847));
  INV_X1    g422(.A(G288), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(G16), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT33), .B(G1976), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n845), .A2(new_n846), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n734), .A2(G22), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(G166), .B2(new_n734), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G1971), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n828), .B(new_n839), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(KEYINPUT92), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n860), .A2(new_n862), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n825), .B1(new_n863), .B2(new_n864), .ZN(G311));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n863), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n866), .A2(new_n733), .A3(new_n818), .A4(new_n824), .ZN(G150));
  NOR2_X1   g442(.A1(new_n615), .A2(new_n623), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT39), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n868), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(G80), .A2(G543), .ZN(new_n872));
  INV_X1    g447(.A(G67), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n512), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G651), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n510), .A2(G93), .A3(new_n511), .A4(new_n520), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  XNOR2_X1  g452(.A(KEYINPUT103), .B(G55), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n520), .A2(new_n878), .A3(G543), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(new_n876), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n875), .B(KEYINPUT105), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n556), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n881), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n887), .A2(new_n888), .B1(G651), .B2(new_n874), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n554), .A2(G651), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n547), .B1(new_n890), .B2(new_n549), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n889), .A2(new_n891), .A3(KEYINPUT105), .A4(new_n555), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n871), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n871), .A2(new_n893), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n894), .A2(new_n895), .A3(G860), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT106), .Z(new_n897));
  NAND2_X1  g472(.A1(new_n882), .A2(G860), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT37), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(G145));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n797), .B(G164), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n748), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(new_n779), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(new_n748), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n748), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n780), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n640), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n480), .A2(G130), .A3(G2105), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n480), .A2(G142), .A3(new_n463), .ZN(new_n911));
  OR2_X1    g486(.A1(G106), .A2(G2105), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n912), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT107), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n910), .A2(new_n911), .A3(new_n916), .A4(new_n913), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n834), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n834), .B1(new_n915), .B2(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n909), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n915), .A2(new_n917), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n835), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n918), .A3(new_n640), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n904), .A2(new_n908), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n903), .A2(new_n779), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n906), .A2(new_n780), .A3(new_n907), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n927), .A2(new_n928), .B1(new_n924), .B2(new_n921), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n901), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n636), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n490), .A2(new_n491), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n490), .A2(new_n491), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n932), .A2(new_n804), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n804), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G162), .A2(G160), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n804), .A3(new_n933), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n636), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n927), .A2(new_n924), .A3(new_n928), .A4(new_n921), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(new_n941), .B2(KEYINPUT108), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n930), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n925), .B1(new_n904), .B2(new_n908), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n941), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n945), .B2(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g523(.A1(G290), .A2(G288), .ZN(new_n949));
  NOR2_X1   g524(.A1(G290), .A2(G288), .ZN(new_n950));
  OAI21_X1  g525(.A(G166), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OR2_X1    g526(.A1(G290), .A2(G288), .ZN(new_n952));
  NAND2_X1  g527(.A1(G290), .A2(G288), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(G303), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G305), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n954), .A3(new_n841), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n958), .B(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT109), .B(G299), .C1(new_n605), .C2(new_n612), .ZN(new_n961));
  NAND2_X1  g536(.A1(G299), .A2(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n603), .A2(new_n604), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n567), .A2(new_n568), .A3(new_n965), .A4(new_n573), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n961), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT41), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n961), .A2(new_n967), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT111), .B(KEYINPUT41), .Z(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n627), .A2(new_n893), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n627), .A2(new_n893), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n971), .B(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n960), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n983), .A2(KEYINPUT112), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n977), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n958), .B(KEYINPUT42), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n983), .B2(KEYINPUT112), .ZN(new_n988));
  OAI21_X1  g563(.A(G868), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n882), .A2(new_n625), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(G295));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n990), .ZN(G331));
  XNOR2_X1  g567(.A(KEYINPUT113), .B(KEYINPUT43), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n886), .A2(G171), .A3(new_n892), .ZN(new_n994));
  AOI21_X1  g569(.A(G171), .B1(new_n886), .B2(new_n892), .ZN(new_n995));
  OAI21_X1  g570(.A(G286), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n893), .A2(G301), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n886), .A2(G171), .A3(new_n892), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(G168), .A3(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n996), .A2(new_n999), .A3(new_n968), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n996), .A2(new_n999), .B1(new_n973), .B2(new_n970), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n958), .A2(KEYINPUT114), .ZN(new_n1003));
  AOI21_X1  g578(.A(G37), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT114), .B(new_n958), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n993), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G37), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n971), .A2(new_n972), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(KEYINPUT41), .B2(new_n971), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n994), .A2(new_n995), .A3(G286), .ZN(new_n1010));
  AOI21_X1  g585(.A(G168), .B1(new_n997), .B2(new_n998), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n980), .A2(new_n999), .A3(new_n996), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n958), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n974), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n996), .A2(new_n999), .A3(new_n968), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n957), .A3(new_n956), .A4(new_n1016), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n1007), .A2(new_n1014), .A3(new_n1017), .A4(new_n993), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1006), .A2(new_n1018), .A3(KEYINPUT44), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1004), .A2(new_n1005), .A3(new_n993), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(new_n1017), .A3(new_n1007), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT43), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1019), .B1(KEYINPUT44), .B2(new_n1023), .ZN(G397));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n498), .B2(new_n502), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n478), .A2(G2105), .ZN(new_n1030));
  INV_X1    g605(.A(new_n471), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n470), .B1(new_n465), .B2(new_n467), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1030), .B(G40), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n797), .B(G2067), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(new_n748), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1034), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(G1996), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1038), .B2(KEYINPUT46), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(KEYINPUT46), .B2(new_n1038), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT47), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n748), .B(new_n688), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1035), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n835), .A2(new_n838), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n834), .A2(new_n837), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1037), .A2(G1986), .A3(G290), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1047), .A2(new_n1037), .B1(KEYINPUT48), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(KEYINPUT48), .B2(new_n1048), .ZN(new_n1050));
  XOR2_X1   g625(.A(new_n1044), .B(KEYINPUT126), .Z(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1051), .A2(new_n1052), .B1(G2067), .B2(new_n797), .ZN(new_n1053));
  AOI211_X1 g628(.A(new_n1041), .B(new_n1050), .C1(new_n1034), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G303), .A2(G8), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT45), .B(new_n1025), .C1(new_n498), .C2(new_n502), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(new_n1033), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1026), .A2(new_n1061), .A3(new_n1028), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1029), .A2(KEYINPUT116), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1971), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n1025), .C1(new_n498), .C2(new_n502), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1067), .A2(G40), .A3(G160), .A4(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(G2090), .ZN(new_n1071));
  OAI211_X1 g646(.A(G8), .B(new_n1057), .C1(new_n1066), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT117), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1074), .A2(G1971), .B1(G2090), .B2(new_n1070), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(G8), .A4(new_n1057), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1057), .B1(new_n1075), .B2(G8), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  OAI221_X1 g655(.A(G8), .B1(new_n1080), .B2(G288), .C1(new_n1033), .C2(new_n1026), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1082), .B(new_n1083), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1033), .A2(new_n1026), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1089), .A2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(new_n585), .ZN(new_n1091));
  OAI21_X1  g666(.A(G1981), .B1(new_n583), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT120), .ZN(new_n1093));
  INV_X1    g668(.A(G1981), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n584), .A2(new_n1094), .A3(new_n586), .A4(new_n587), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(G1981), .C1(new_n583), .C2(new_n1091), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1093), .A2(new_n1095), .A3(KEYINPUT49), .A4(new_n1097), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1090), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1081), .A2(KEYINPUT52), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1087), .A2(new_n1086), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT119), .B1(new_n1104), .B2(new_n1081), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1088), .A2(new_n1102), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1079), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1033), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT45), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1026), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1108), .B(new_n1110), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n756), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1033), .B1(KEYINPUT50), .B2(new_n1026), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n806), .A3(new_n1069), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G8), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(G286), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1078), .A2(new_n1107), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT63), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1078), .A2(new_n1107), .A3(new_n1120), .A4(new_n1117), .ZN(new_n1121));
  AND4_X1   g696(.A1(new_n1103), .A2(new_n1088), .A3(new_n1102), .A4(new_n1105), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1073), .A2(new_n1122), .A3(new_n1077), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1102), .A2(new_n1080), .A3(new_n848), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1095), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1090), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1119), .A2(new_n1121), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(G8), .C1(new_n1115), .C2(G286), .ZN(new_n1130));
  NAND2_X1  g705(.A1(G286), .A2(G8), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g709(.A(KEYINPUT124), .B(new_n1131), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1130), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1116), .A2(KEYINPUT51), .A3(new_n1131), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT62), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1132), .B(new_n1133), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n1137), .A4(new_n1130), .ZN(new_n1142));
  INV_X1    g717(.A(G2078), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n1074), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1113), .A2(KEYINPUT121), .A3(new_n1069), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1070), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1961), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1143), .A2(KEYINPUT53), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1111), .B2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1151), .A2(G171), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1139), .A2(new_n1142), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT56), .B(G2072), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1060), .A2(new_n1063), .A3(new_n1062), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(G1956), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1070), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(G299), .B(KEYINPUT57), .Z(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n822), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1089), .A2(G2067), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1155), .A2(new_n1159), .A3(new_n1157), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n616), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1155), .A2(new_n1159), .A3(new_n1157), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1159), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT123), .ZN(new_n1172));
  NAND2_X1  g747(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1060), .A2(new_n1063), .A3(new_n688), .A4(new_n1062), .ZN(new_n1175));
  XOR2_X1   g750(.A(KEYINPUT58), .B(G1341), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n1089), .A2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n556), .B(new_n1174), .C1(new_n1175), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1173), .B1(new_n1179), .B2(new_n557), .ZN(new_n1180));
  OAI22_X1  g755(.A1(new_n1170), .A2(new_n1172), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1161), .A2(new_n1165), .A3(new_n1172), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1171), .A2(KEYINPUT123), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n613), .A2(KEYINPUT60), .A3(new_n614), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1164), .A2(new_n1187), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1162), .A2(new_n1186), .A3(new_n1163), .ZN(new_n1189));
  OAI22_X1  g764(.A1(new_n1188), .A2(new_n1189), .B1(KEYINPUT60), .B2(new_n616), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1167), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(G171), .B(KEYINPUT54), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1151), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1060), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1029), .A2(KEYINPUT53), .A3(new_n1143), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1149), .B(new_n1192), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1194), .B(new_n1197), .C1(new_n1138), .C2(new_n1136), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1153), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1078), .A2(new_n1107), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1128), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  XOR2_X1   g778(.A(G290), .B(G1986), .Z(new_n1204));
  AOI21_X1  g779(.A(new_n1037), .B1(new_n1047), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1054), .B1(new_n1203), .B2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(G319), .ZN(new_n1208));
  OR2_X1    g782(.A1(G227), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g783(.A(new_n1209), .B1(new_n668), .B2(new_n669), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n721), .A2(new_n724), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1211), .B1(new_n943), .B2(new_n946), .ZN(new_n1212));
  OAI21_X1  g786(.A(new_n1212), .B1(new_n1006), .B2(new_n1018), .ZN(G225));
  NAND2_X1  g787(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1214));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n1215));
  OAI211_X1 g789(.A(new_n1212), .B(new_n1215), .C1(new_n1006), .C2(new_n1018), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1214), .A2(new_n1216), .ZN(G308));
endmodule


