//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1306, new_n1307, new_n1308, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G250), .B1(G257), .B2(G264), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n217), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT64), .Z(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n219), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n213), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G50), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n206), .B1(new_n201), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT66), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n257), .A2(new_n259), .B1(G150), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n251), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n213), .A3(new_n249), .ZN(new_n264));
  OAI21_X1  g0064(.A(G50), .B1(new_n206), .B2(G1), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n264), .A2(new_n265), .B1(G50), .B2(new_n263), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT70), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NOR4_X1   g0071(.A1(new_n262), .A2(new_n269), .A3(new_n271), .A4(new_n266), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G222), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G223), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n279), .B(new_n280), .C1(G77), .C2(new_n275), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  OAI211_X1 g0084(.A(G1), .B(G13), .C1(new_n258), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n285), .A3(G274), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n282), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G226), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n281), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G190), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n280), .A2(new_n293), .A3(new_n282), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(G226), .B2(new_n288), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n281), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT71), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n292), .A2(new_n298), .B1(G200), .B2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n271), .B1(new_n262), .B2(new_n266), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n274), .A2(new_n299), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(G200), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n291), .B1(new_n290), .B2(G190), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n296), .A2(KEYINPUT71), .A3(new_n297), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n301), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT70), .B1(new_n267), .B2(KEYINPUT9), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n272), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT10), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n267), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n290), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n311), .B(new_n313), .C1(G169), .C2(new_n290), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT79), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n294), .B1(G232), .B2(new_n288), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT77), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT3), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(G33), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(G33), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n258), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(G223), .A2(G1698), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(G226), .B2(new_n277), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n323), .A2(new_n325), .B1(new_n258), .B2(new_n223), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n280), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n317), .A2(new_n297), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(G200), .B1(new_n317), .B2(new_n327), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n316), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n317), .A2(new_n327), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n317), .A2(new_n327), .A3(new_n297), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(KEYINPUT79), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n321), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(new_n206), .C1(KEYINPUT78), .C2(KEYINPUT7), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n275), .B2(G20), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n221), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G58), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n221), .ZN(new_n345));
  OAI21_X1  g0145(.A(G20), .B1(new_n345), .B2(new_n201), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n260), .A2(G159), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n337), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n348), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n323), .A2(new_n351), .A3(new_n206), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G68), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n323), .B2(new_n206), .ZN(new_n354));
  OAI211_X1 g0154(.A(KEYINPUT16), .B(new_n350), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n349), .A2(new_n355), .A3(new_n250), .ZN(new_n356));
  INV_X1    g0156(.A(new_n264), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n206), .A2(G1), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n256), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n263), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n357), .A2(new_n359), .B1(new_n360), .B2(new_n256), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n336), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT17), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n356), .A2(new_n361), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n331), .A2(G169), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n317), .A2(new_n327), .A3(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT18), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n366), .A2(new_n372), .A3(new_n369), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n336), .A2(new_n362), .A3(KEYINPUT17), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n365), .A2(new_n371), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n264), .A2(new_n221), .A3(new_n358), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n360), .A2(new_n221), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT12), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT76), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(KEYINPUT76), .A3(new_n380), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n260), .A2(G50), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT74), .ZN(new_n386));
  INV_X1    g0186(.A(new_n259), .ZN(new_n387));
  INV_X1    g0187(.A(G77), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n387), .A2(new_n388), .B1(new_n206), .B2(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n250), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT11), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n383), .A2(new_n384), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n237), .A2(G1698), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n275), .B(new_n395), .C1(G226), .C2(G1698), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G97), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n280), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n286), .B1(new_n287), .B2(new_n222), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n394), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n285), .B1(new_n396), .B2(new_n397), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n403), .A2(new_n400), .A3(KEYINPUT13), .ZN(new_n404));
  OAI21_X1  g0204(.A(G200), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(new_n401), .A3(new_n394), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT73), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n399), .A2(new_n401), .A3(KEYINPUT73), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n394), .A2(KEYINPUT72), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n410), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n399), .A2(new_n401), .A3(KEYINPUT73), .A4(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n408), .A2(new_n411), .A3(G190), .A4(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n393), .A2(new_n405), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(G169), .B1(new_n402), .B2(new_n404), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT14), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n408), .A2(new_n411), .A3(G179), .A4(new_n413), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(G169), .C1(new_n402), .C2(new_n404), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n392), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n294), .B1(G244), .B2(new_n288), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n338), .A2(new_n321), .A3(G238), .A4(G1698), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT68), .B(G107), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n275), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n277), .A2(G232), .ZN(new_n427));
  OR3_X1    g0227(.A1(new_n339), .A2(KEYINPUT67), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT67), .B1(new_n339), .B2(new_n427), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n423), .B1(new_n430), .B2(new_n285), .ZN(new_n431));
  INV_X1    g0231(.A(G169), .ZN(new_n432));
  INV_X1    g0232(.A(new_n260), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n256), .A2(new_n433), .B1(new_n206), .B2(new_n388), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT15), .B(G87), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n387), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n250), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n358), .A2(new_n388), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n357), .A2(new_n438), .B1(new_n388), .B2(new_n360), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT69), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n437), .A2(KEYINPUT69), .A3(new_n439), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n431), .A2(new_n432), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n431), .A2(G179), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n431), .A2(G200), .ZN(new_n447));
  OAI211_X1 g0247(.A(G190), .B(new_n423), .C1(new_n430), .C2(new_n285), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n442), .A4(new_n443), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n415), .A2(new_n422), .A3(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n315), .A2(new_n375), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n360), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n205), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n263), .A2(new_n456), .A3(new_n213), .A4(new_n249), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n425), .B1(new_n340), .B2(new_n342), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n463));
  INV_X1    g0263(.A(G107), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n462), .A2(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G97), .A3(new_n464), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n206), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n433), .A2(new_n388), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n460), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n459), .B1(new_n472), .B2(new_n251), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT4), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n320), .A2(new_n322), .A3(G244), .A4(new_n321), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(G1698), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n224), .B2(new_n277), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n479), .A2(new_n275), .B1(G33), .B2(G283), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n477), .A2(KEYINPUT81), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT81), .B1(new_n477), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n280), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G257), .A3(new_n285), .ZN(new_n490));
  OR2_X1    g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n486), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n285), .A3(G274), .A4(new_n485), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n483), .A2(G190), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n477), .A2(new_n480), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT81), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n477), .A2(KEYINPUT81), .A3(new_n480), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n285), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n494), .B(KEYINPUT82), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n474), .B(new_n496), .C1(new_n503), .C2(new_n332), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT82), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n494), .B(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n483), .A2(new_n312), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n499), .A2(new_n500), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n494), .B1(new_n508), .B2(new_n280), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n473), .C1(new_n509), .C2(G169), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n322), .A2(new_n321), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT83), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n222), .A2(G1698), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n320), .A4(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n320), .A2(new_n322), .A3(new_n514), .A4(new_n321), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT83), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G116), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n258), .A2(new_n519), .ZN(new_n520));
  AND4_X1   g0320(.A1(G244), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(G1698), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n285), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n280), .A2(new_n293), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n485), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n205), .A2(G45), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n285), .A2(G250), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(G169), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n528), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n476), .A2(new_n277), .B1(new_n258), .B2(new_n519), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n515), .B2(new_n517), .ZN(new_n532));
  OAI211_X1 g0332(.A(G179), .B(new_n530), .C1(new_n532), .C2(new_n285), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n435), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n263), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n221), .A2(G20), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n320), .A2(new_n322), .A3(new_n537), .A4(new_n321), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT68), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G107), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G87), .A2(G97), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n397), .A2(new_n206), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n387), .A2(KEYINPUT19), .A3(new_n454), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n538), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n536), .B1(new_n548), .B2(new_n250), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n457), .A2(new_n435), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT84), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n536), .B(new_n550), .C1(new_n548), .C2(new_n250), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT84), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n534), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT21), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n249), .A2(new_n213), .B1(G20), .B2(new_n519), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G283), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n560), .B(new_n206), .C1(G33), .C2(new_n454), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT20), .B1(new_n559), .B2(new_n561), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n360), .A2(new_n519), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n457), .B2(new_n519), .ZN(new_n566));
  OAI21_X1  g0366(.A(G169), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G257), .A2(G1698), .ZN(new_n568));
  INV_X1    g0368(.A(G264), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(G1698), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n570), .A2(new_n321), .A3(new_n320), .A4(new_n322), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n339), .A2(G303), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n285), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n489), .A2(new_n285), .ZN(new_n574));
  INV_X1    g0374(.A(G270), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n493), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n558), .B1(new_n567), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n573), .B2(new_n576), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n526), .B1(new_n491), .B2(new_n486), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n280), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(G270), .B1(new_n524), .B2(new_n580), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n569), .A2(G1698), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(G257), .B2(G1698), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n572), .B1(new_n323), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n280), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n586), .A3(G190), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n564), .A2(new_n566), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n579), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n573), .A2(new_n576), .A3(new_n312), .ZN(new_n590));
  INV_X1    g0390(.A(new_n457), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G116), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(new_n565), .C1(new_n562), .C2(new_n563), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n582), .A2(new_n586), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n595), .A2(KEYINPUT21), .A3(G169), .A4(new_n593), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n578), .A2(new_n589), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(G200), .B1(new_n523), .B2(new_n528), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n548), .A2(new_n250), .ZN(new_n599));
  INV_X1    g0399(.A(new_n536), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n591), .A2(G87), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G190), .B(new_n530), .C1(new_n532), .C2(new_n285), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n557), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n360), .A2(KEYINPUT25), .A3(new_n464), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT25), .B1(new_n360), .B2(new_n464), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n606), .A2(new_n607), .B1(new_n464), .B2(new_n457), .ZN(new_n608));
  AND2_X1   g0408(.A1(KEYINPUT22), .A2(G87), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n320), .A2(new_n322), .A3(new_n321), .A4(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n520), .A2(KEYINPUT23), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n541), .A2(G107), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT23), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n610), .A2(new_n611), .B1(new_n614), .B2(G20), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT22), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n339), .B2(new_n223), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G20), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT24), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n275), .A2(G87), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(new_n616), .B1(G20), .B2(new_n618), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT24), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n610), .A2(new_n611), .ZN(new_n625));
  INV_X1    g0425(.A(new_n425), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n206), .B1(new_n626), .B2(KEYINPUT23), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n608), .B1(new_n629), .B2(new_n250), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n574), .A2(new_n569), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n224), .A2(G1698), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n320), .A2(new_n322), .A3(new_n632), .A4(new_n321), .ZN(new_n633));
  NAND2_X1  g0433(.A1(G33), .A2(G294), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(G257), .A2(G1698), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n320), .A2(new_n322), .A3(new_n321), .A4(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(KEYINPUT85), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(KEYINPUT85), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n631), .B1(new_n640), .B2(new_n280), .ZN(new_n641));
  AOI21_X1  g0441(.A(G200), .B1(new_n641), .B2(new_n493), .ZN(new_n642));
  INV_X1    g0442(.A(new_n631), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n633), .A2(new_n634), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n512), .A2(new_n645), .A3(new_n320), .A4(new_n636), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n637), .A2(KEYINPUT85), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n643), .B(new_n493), .C1(new_n648), .C2(new_n285), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G190), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n630), .B1(new_n642), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT86), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n432), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n640), .A2(new_n280), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(new_n312), .A3(new_n643), .A4(new_n493), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n251), .B1(new_n621), .B2(new_n628), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n653), .B(new_n655), .C1(new_n656), .C2(new_n608), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n651), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n652), .B1(new_n651), .B2(new_n657), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n511), .B(new_n605), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n453), .A2(new_n660), .ZN(G372));
  AND2_X1   g0461(.A1(new_n371), .A2(new_n373), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n336), .A2(KEYINPUT17), .A3(new_n362), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT17), .B1(new_n336), .B2(new_n362), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n446), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n415), .A2(new_n667), .B1(new_n392), .B2(new_n421), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n662), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n310), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n314), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n557), .A2(new_n604), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n673), .B2(new_n510), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n649), .A2(new_n332), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(G190), .B2(new_n649), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n518), .A2(new_n522), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n528), .B1(new_n678), .B2(new_n280), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n679), .B2(G190), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n676), .A2(new_n630), .B1(new_n680), .B2(new_n598), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n578), .A2(new_n596), .A3(new_n594), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n657), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n681), .A2(new_n683), .A3(new_n510), .A4(new_n504), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n534), .A2(new_n552), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n432), .B1(new_n501), .B2(new_n494), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n686), .A2(new_n507), .A3(new_n473), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(new_n604), .A4(new_n685), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n674), .A2(new_n684), .A3(new_n685), .A4(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n672), .B1(new_n691), .B2(new_n453), .ZN(G369));
  NOR2_X1   g0492(.A1(new_n658), .A2(new_n659), .ZN(new_n693));
  INV_X1    g0493(.A(new_n630), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G213), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n693), .B1(new_n694), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n657), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n578), .A2(new_n596), .A3(new_n594), .ZN(new_n704));
  INV_X1    g0504(.A(new_n700), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n588), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n597), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n706), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT87), .Z(new_n711));
  NOR2_X1   g0511(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n682), .A2(new_n700), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n693), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n702), .B2(new_n705), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n717), .ZN(G399));
  NOR2_X1   g0518(.A1(new_n210), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n544), .A2(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n215), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n685), .A2(new_n604), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT26), .B1(new_n725), .B2(new_n510), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n549), .A2(new_n555), .A3(new_n551), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n555), .B1(new_n549), .B2(new_n551), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n729), .A2(new_n534), .B1(new_n680), .B2(new_n598), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n688), .A3(new_n687), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n684), .A2(new_n726), .A3(new_n731), .A4(new_n685), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n732), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT29), .B1(new_n690), .B2(new_n705), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n679), .A2(G179), .A3(new_n577), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n483), .A2(new_n506), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n649), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n679), .A2(new_n641), .A3(new_n590), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n483), .A2(new_n495), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n643), .B1(new_n648), .B2(new_n285), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n582), .A2(new_n586), .A3(G179), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n509), .A2(KEYINPUT30), .A3(new_n679), .A4(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n739), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n700), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n751), .B(new_n752), .C1(new_n660), .C2(new_n700), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n736), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n724), .B1(new_n756), .B2(G1), .ZN(G364));
  AND2_X1   g0557(.A1(new_n206), .A2(G13), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n205), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n719), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n711), .B(new_n762), .C1(G330), .C2(new_n709), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n209), .A2(new_n275), .ZN(new_n764));
  INV_X1    g0564(.A(G355), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n765), .B1(G116), .B2(new_n209), .ZN(new_n766));
  INV_X1    g0566(.A(new_n323), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n210), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n484), .B2(new_n216), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n244), .A2(new_n484), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n213), .B1(G20), .B2(new_n432), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n761), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n206), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n454), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n206), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n297), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G107), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n206), .A2(new_n312), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n786), .B1(new_n252), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n787), .A2(G190), .A3(new_n332), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n782), .B(new_n789), .C1(G58), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n783), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT88), .B(KEYINPUT32), .Z(new_n796));
  NAND3_X1  g0596(.A1(new_n795), .A2(G159), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(new_n795), .B2(G159), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(G87), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n787), .A2(new_n297), .A3(G200), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n275), .B1(new_n802), .B2(new_n221), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n787), .A2(new_n793), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n803), .B1(G77), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n792), .A2(new_n797), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  INV_X1    g0608(.A(G329), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n784), .A2(new_n808), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT89), .Z(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT33), .B(G317), .Z(new_n813));
  OAI221_X1 g0613(.A(new_n339), .B1(new_n804), .B2(new_n812), .C1(new_n802), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G322), .ZN(new_n815));
  INV_X1    g0615(.A(G326), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n790), .A2(new_n815), .B1(new_n788), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n781), .A2(new_n818), .B1(new_n799), .B2(new_n819), .ZN(new_n820));
  OR3_X1    g0620(.A1(new_n814), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n807), .B1(new_n811), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n779), .B1(new_n822), .B2(new_n776), .ZN(new_n823));
  INV_X1    g0623(.A(new_n775), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n709), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n763), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n442), .A2(new_n443), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n700), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n449), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n446), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT93), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n444), .A2(new_n445), .A3(new_n705), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n449), .A2(new_n829), .B1(new_n444), .B2(new_n445), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n444), .A2(new_n445), .A3(new_n705), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT93), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n691), .B2(new_n700), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n832), .B1(new_n831), .B2(new_n833), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT93), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n690), .A2(new_n842), .A3(new_n705), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n761), .B1(new_n844), .B2(new_n754), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n754), .B2(new_n844), .ZN(new_n846));
  INV_X1    g0646(.A(new_n776), .ZN(new_n847));
  INV_X1    g0647(.A(new_n802), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G150), .B1(new_n805), .B2(G159), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n791), .A2(G143), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n788), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n323), .B1(new_n795), .B2(G132), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n781), .A2(new_n344), .B1(new_n799), .B2(new_n252), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(G68), .B2(new_n785), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n804), .A2(new_n519), .B1(new_n794), .B2(new_n812), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n275), .B(new_n860), .C1(G283), .C2(new_n848), .ZN(new_n861));
  INV_X1    g0661(.A(new_n782), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n790), .A2(new_n818), .B1(new_n788), .B2(new_n819), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(G107), .B2(new_n800), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n785), .A2(G87), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n861), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n847), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n847), .A2(new_n774), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT90), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT91), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n762), .B(new_n867), .C1(new_n388), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT92), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n774), .B2(new_n842), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n846), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  NAND2_X1  g0676(.A1(new_n467), .A2(new_n469), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n214), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  OR3_X1    g0681(.A1(new_n215), .A2(new_n388), .A3(new_n345), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n252), .A2(G68), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n205), .B(G13), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n698), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n662), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n554), .B1(new_n529), .B2(new_n533), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n649), .A2(G179), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n630), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n704), .B1(new_n890), .B2(new_n653), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n651), .A2(new_n604), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n888), .B1(new_n893), .B2(new_n511), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n688), .B1(new_n730), .B2(new_n687), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n896));
  NOR4_X1   g0696(.A1(new_n510), .A2(new_n896), .A3(new_n888), .A4(KEYINPUT26), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n700), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n836), .B1(new_n899), .B2(new_n842), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n415), .A2(new_n422), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n393), .A2(new_n705), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n422), .B(new_n415), .C1(new_n393), .C2(new_n705), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT94), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(KEYINPUT94), .B(new_n350), .C1(new_n353), .C2(new_n354), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n337), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n355), .A2(new_n250), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(KEYINPUT95), .A3(new_n361), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT95), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT16), .B1(new_n908), .B2(new_n909), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n913), .B1(new_n918), .B2(new_n911), .ZN(new_n919));
  INV_X1    g0719(.A(new_n361), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n916), .A2(new_n921), .A3(new_n886), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n916), .A2(new_n921), .A3(new_n369), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n363), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  XNOR2_X1  g0725(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n366), .A2(new_n886), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n363), .A2(new_n370), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n922), .B1(new_n665), .B2(new_n662), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT38), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT38), .ZN(new_n933));
  INV_X1    g0733(.A(new_n928), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n924), .B2(KEYINPUT37), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n933), .B1(new_n935), .B2(new_n930), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n887), .B1(new_n907), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n935), .A2(new_n933), .A3(new_n930), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n927), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n375), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n363), .A2(new_n370), .A3(new_n927), .ZN(new_n945));
  INV_X1    g0745(.A(new_n926), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n928), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n942), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n939), .B1(new_n940), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n932), .A2(KEYINPUT39), .A3(new_n936), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n422), .A2(new_n700), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n938), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT98), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n732), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n452), .B(new_n956), .C1(new_n899), .C2(KEYINPUT29), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT99), .ZN(new_n958));
  INV_X1    g0758(.A(new_n734), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT99), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(new_n960), .A3(new_n452), .A4(new_n956), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n671), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n955), .B(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n949), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n932), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n838), .B1(new_n903), .B2(new_n904), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n753), .A2(new_n966), .A3(KEYINPUT40), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT100), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n965), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n930), .B1(new_n925), .B2(new_n928), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n949), .B1(new_n971), .B2(KEYINPUT38), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT100), .B1(new_n972), .B2(new_n967), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n753), .A2(new_n966), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT38), .B1(new_n929), .B2(new_n931), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n976), .B2(new_n940), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT40), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n753), .A2(new_n452), .ZN(new_n981));
  OAI21_X1  g0781(.A(G330), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n980), .B2(new_n981), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n963), .A2(new_n983), .B1(new_n205), .B2(new_n758), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n963), .A2(new_n983), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n885), .B1(new_n984), .B2(new_n985), .ZN(G367));
  NAND2_X1  g0786(.A1(new_n768), .A2(new_n234), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n777), .C1(new_n209), .C2(new_n435), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n781), .A2(new_n221), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G150), .B2(new_n791), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT107), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n784), .A2(new_n388), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n275), .B1(new_n794), .B2(new_n851), .C1(new_n344), .C2(new_n799), .ZN(new_n993));
  INV_X1    g0793(.A(new_n788), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n992), .B(new_n993), .C1(G143), .C2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(G159), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n802), .A2(new_n996), .B1(new_n804), .B2(new_n252), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT108), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n991), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n323), .B1(new_n788), .B2(new_n812), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n802), .A2(new_n818), .B1(new_n804), .B2(new_n808), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G317), .C2(new_n795), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n781), .A2(new_n425), .B1(new_n790), .B2(new_n819), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n784), .A2(new_n454), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n800), .A2(G116), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT46), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1002), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n999), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT47), .Z(new_n1010));
  OAI211_X1 g0810(.A(new_n761), .B(new_n988), .C1(new_n1010), .C2(new_n847), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT109), .Z(new_n1012));
  NOR2_X1   g0812(.A1(new_n602), .A2(new_n705), .ZN(new_n1013));
  MUX2_X1   g0813(.A(new_n725), .B(new_n685), .S(new_n1013), .Z(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT101), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1012), .B1(new_n824), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT110), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT106), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n712), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n511), .B1(new_n474), .B2(new_n705), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n510), .B2(new_n705), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT102), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n717), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT105), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT44), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n712), .A2(new_n1018), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1021), .B(KEYINPUT102), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n717), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT45), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1028), .B(new_n1029), .C1(new_n1031), .C2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT105), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1032), .A2(new_n717), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1038), .A2(KEYINPUT44), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1019), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1026), .B1(new_n1038), .B2(KEYINPUT44), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT44), .B2(new_n1038), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1044), .A2(new_n1045), .B1(new_n1018), .B2(new_n712), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1019), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .A4(new_n1028), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1041), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n703), .A2(new_n715), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n693), .B2(new_n715), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(new_n711), .Z(new_n1052));
  AOI21_X1  g0852(.A(new_n755), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n719), .B(KEYINPUT41), .Z(new_n1054));
  OAI21_X1  g0854(.A(new_n759), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n510), .B1(new_n1023), .B2(new_n657), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT42), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n716), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1057), .B1(new_n1023), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1032), .A2(KEYINPUT42), .A3(new_n716), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n705), .A2(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1015), .B(KEYINPUT43), .ZN(new_n1062));
  OAI21_X1  g0862(.A(KEYINPUT104), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1056), .A2(new_n705), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT104), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1062), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1015), .A2(KEYINPUT43), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1064), .A2(new_n1065), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT103), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT103), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1061), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n713), .A2(new_n1023), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1070), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1017), .B1(new_n1055), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(G387));
  INV_X1    g0882(.A(new_n1052), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1083), .A2(new_n755), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n755), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n719), .A3(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n764), .A2(new_n721), .B1(G107), .B2(new_n209), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n769), .B1(new_n240), .B2(G45), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n721), .B(KEYINPUT111), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n484), .B1(new_n221), .B2(new_n388), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n256), .A2(G50), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT50), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1090), .B(new_n1094), .C1(new_n1093), .C2(new_n1092), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1088), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G159), .A2(new_n994), .B1(new_n800), .B2(G77), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n252), .B2(new_n790), .C1(new_n435), .C2(new_n781), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n848), .A2(new_n257), .B1(new_n795), .B2(G150), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n221), .B2(new_n804), .ZN(new_n1100));
  NOR4_X1   g0900(.A1(new_n1098), .A2(new_n323), .A3(new_n1004), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n781), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(G283), .B1(new_n800), .B2(G294), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G311), .A2(new_n848), .B1(new_n994), .B2(G322), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT112), .ZN(new_n1105));
  INV_X1    g0905(.A(G317), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n790), .A2(new_n1106), .B1(new_n804), .B2(new_n819), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT113), .Z(new_n1110));
  OAI21_X1  g0910(.A(new_n1103), .B1(new_n1110), .B2(KEYINPUT48), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(KEYINPUT48), .B2(new_n1110), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1112), .A2(KEYINPUT49), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n323), .B1(new_n794), .B2(new_n816), .C1(new_n519), .C2(new_n784), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1112), .B2(KEYINPUT49), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1101), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n761), .B1(new_n778), .B2(new_n1096), .C1(new_n1116), .C2(new_n847), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n703), .B2(new_n775), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1052), .B2(new_n760), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1087), .A2(new_n1119), .ZN(G393));
  NAND2_X1  g0920(.A1(new_n768), .A2(new_n247), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n777), .C1(new_n454), .C2(new_n209), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n802), .A2(new_n252), .B1(new_n804), .B2(new_n256), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1102), .A2(G77), .B1(new_n800), .B2(G68), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n767), .A3(new_n865), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(G143), .C2(new_n795), .ZN(new_n1126));
  INV_X1    g0926(.A(G150), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n790), .A2(new_n996), .B1(new_n788), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n790), .A2(new_n812), .B1(new_n788), .B2(new_n1106), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT52), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n786), .B1(new_n808), .B2(new_n799), .C1(new_n519), .C2(new_n781), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n339), .B1(new_n802), .B2(new_n819), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n804), .A2(new_n818), .B1(new_n794), .B2(new_n815), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1126), .A2(new_n1130), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n761), .B(new_n1122), .C1(new_n1137), .C2(new_n847), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1023), .B2(new_n775), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1049), .B2(new_n760), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1084), .A2(new_n1049), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n719), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1084), .A2(new_n1049), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(G390));
  OAI22_X1  g0944(.A1(new_n804), .A2(new_n454), .B1(new_n794), .B2(new_n818), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n275), .B(new_n1145), .C1(new_n626), .C2(new_n848), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n221), .B2(new_n784), .C1(new_n223), .C2(new_n799), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G77), .A2(new_n1102), .B1(new_n791), .B2(G116), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n808), .B2(new_n788), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G128), .A2(new_n994), .B1(new_n785), .B2(G50), .ZN(new_n1150));
  INV_X1    g0950(.A(G132), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n790), .C1(new_n996), .C2(new_n781), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n848), .A2(G137), .B1(new_n795), .B2(G125), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n799), .A2(KEYINPUT53), .A3(new_n1127), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT53), .B1(new_n799), .B2(new_n1127), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n339), .B1(new_n805), .B2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1147), .A2(new_n1149), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT117), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n847), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1161), .B2(new_n1160), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1163), .B(new_n761), .C1(new_n257), .C2(new_n870), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n950), .A2(new_n951), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n773), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n753), .A2(new_n905), .A3(G330), .A4(new_n842), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(KEYINPUT115), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n732), .A2(new_n842), .A3(new_n705), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n833), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n952), .B1(new_n1171), .B2(new_n905), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n965), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1168), .A2(KEYINPUT115), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n952), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n843), .A2(new_n833), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n905), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n950), .A2(new_n951), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1169), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1176), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n932), .A2(KEYINPUT39), .A3(new_n936), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT39), .B1(new_n932), .B2(new_n964), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1172), .A2(new_n965), .B1(new_n1168), .B2(KEYINPUT115), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1169), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1166), .B1(new_n1188), .B2(new_n760), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n730), .A2(new_n510), .A3(new_n504), .A4(new_n597), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n693), .A2(new_n1190), .A3(new_n700), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n751), .A2(new_n752), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G330), .B(new_n842), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n906), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1171), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1194), .A2(new_n1167), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n900), .B1(new_n1194), .B2(new_n1167), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n753), .A2(new_n452), .A3(G330), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT116), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT116), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n753), .A2(new_n452), .A3(new_n1201), .A4(G330), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n960), .B1(new_n735), .B2(new_n452), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n957), .A2(KEYINPUT99), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n672), .B(new_n1203), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1198), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n719), .B1(new_n1188), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n962), .B(new_n1203), .C1(new_n1197), .C2(new_n1196), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1180), .B2(new_n1187), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1189), .B1(new_n1208), .B2(new_n1210), .ZN(G378));
  INV_X1    g1011(.A(KEYINPUT119), .ZN(new_n1212));
  INV_X1    g1012(.A(G330), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n977), .B2(new_n978), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n974), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT118), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n974), .A2(new_n1214), .A3(KEYINPUT118), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n311), .A2(new_n886), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n315), .B(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1220), .B(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AND4_X1   g1023(.A1(new_n1212), .A2(new_n1217), .A3(new_n1218), .A4(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n974), .A2(new_n1214), .A3(new_n1222), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT119), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n1218), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n955), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT121), .B1(new_n1210), .B2(new_n1206), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1175), .A2(new_n1179), .A3(new_n1169), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1186), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1207), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT121), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1206), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1230), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1227), .A2(new_n1212), .A3(new_n1218), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n954), .B(KEYINPUT98), .Z(new_n1239));
  AND3_X1   g1039(.A1(new_n1217), .A2(new_n1218), .A3(new_n1223), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1238), .B(new_n1239), .C1(new_n1240), .C2(new_n1226), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1229), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT57), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1229), .A2(new_n1237), .A3(new_n1241), .A4(KEYINPUT57), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n719), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT120), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1229), .A2(new_n760), .A3(new_n1241), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n761), .B1(new_n869), .B2(G50), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n802), .A2(new_n1151), .B1(new_n804), .B2(new_n851), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G150), .A2(new_n1102), .B1(new_n994), .B2(G125), .ZN(new_n1251));
  INV_X1    g1051(.A(G128), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n790), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1250), .B(new_n1253), .C1(new_n800), .C2(new_n1157), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT59), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n785), .A2(G159), .ZN(new_n1258));
  AOI211_X1 g1058(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n848), .A2(G97), .B1(new_n795), .B2(G283), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n435), .B2(new_n804), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n989), .B(new_n1262), .C1(G77), .C2(new_n800), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n790), .A2(new_n464), .B1(new_n784), .B2(new_n344), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G116), .B2(new_n994), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1263), .A2(new_n284), .A3(new_n323), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT58), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G50), .B1(new_n258), .B2(new_n284), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n767), .B2(G41), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1260), .A2(new_n1268), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1249), .B1(new_n1272), .B2(new_n776), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1222), .B2(new_n774), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1247), .B1(new_n1248), .B2(new_n1274), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1248), .A2(new_n1247), .A3(new_n1274), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1246), .B1(new_n1275), .B2(new_n1276), .ZN(G375));
  INV_X1    g1077(.A(new_n1198), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n906), .A2(new_n773), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n790), .A2(new_n851), .B1(new_n799), .B2(new_n996), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n848), .A2(new_n1157), .B1(new_n795), .B2(G128), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1127), .B2(new_n804), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n781), .A2(new_n252), .B1(new_n788), .B2(new_n1151), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n767), .B1(new_n344), .B2(new_n784), .ZN(new_n1284));
  OR4_X1    g1084(.A1(new_n1280), .A2(new_n1282), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n788), .A2(new_n818), .B1(new_n799), .B2(new_n454), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(G283), .B2(new_n791), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n275), .B1(new_n848), .B2(G116), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n626), .A2(new_n805), .B1(new_n795), .B2(G303), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n992), .B1(new_n535), .B2(new_n1102), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n847), .B1(new_n1285), .B2(new_n1291), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n762), .B(new_n1292), .C1(new_n221), .C2(new_n871), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1278), .A2(new_n760), .B1(new_n1279), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1198), .A2(new_n1206), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1207), .A2(new_n1054), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(G381));
  NOR3_X1   g1099(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1300), .B(KEYINPUT122), .Z(new_n1301));
  NOR3_X1   g1101(.A1(new_n1301), .A2(G390), .A3(G381), .ZN(new_n1302));
  INV_X1    g1102(.A(G378), .ZN(new_n1303));
  INV_X1    g1103(.A(G375), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1302), .A2(new_n1081), .A3(new_n1303), .A4(new_n1304), .ZN(G407));
  NAND2_X1  g1105(.A1(new_n699), .A2(G213), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1303), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(G407), .A2(G213), .A3(new_n1308), .ZN(G409));
  INV_X1    g1109(.A(KEYINPUT125), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1081), .A2(G390), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1081), .A2(G390), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT123), .B1(new_n1081), .B2(G390), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G393), .B(G396), .ZN(new_n1315));
  OAI22_X1  g1115(.A1(new_n1312), .A2(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1081), .A2(G390), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(G393), .B(new_n826), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1317), .A2(KEYINPUT123), .A3(new_n1311), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT124), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1316), .A2(new_n1319), .A3(KEYINPUT124), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1246), .B(G378), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1248), .B(new_n1274), .C1(new_n1242), .C2(new_n1054), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1303), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1209), .A2(KEYINPUT60), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1296), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n720), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1331), .B1(new_n1330), .B2(new_n1329), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1294), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n875), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(G384), .A3(new_n1294), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1328), .A2(new_n1306), .A3(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1307), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1341), .A2(KEYINPUT62), .A3(new_n1337), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1328), .A2(new_n1306), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1336), .A2(G2897), .A3(new_n1307), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1336), .B1(G2897), .B2(new_n1307), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT61), .B1(new_n1344), .B2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1324), .B1(new_n1343), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1344), .A2(new_n1347), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT61), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1341), .A2(KEYINPUT63), .A3(new_n1337), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1350), .A2(new_n1351), .A3(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1320), .ZN(new_n1354));
  AOI211_X1 g1154(.A(new_n1307), .B(new_n1336), .C1(new_n1325), .C2(new_n1327), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1354), .B1(new_n1355), .B2(KEYINPUT63), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1353), .A2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1310), .B1(new_n1349), .B2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT63), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1320), .B1(new_n1338), .B2(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1360), .A2(new_n1352), .A3(new_n1348), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1347), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1351), .B1(new_n1362), .B2(new_n1341), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1363), .B1(new_n1340), .B2(new_n1342), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1361), .B(KEYINPUT125), .C1(new_n1364), .C2(new_n1324), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1358), .A2(new_n1365), .ZN(G405));
  NOR2_X1   g1166(.A1(new_n1304), .A2(G378), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(KEYINPUT126), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT126), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1325), .A2(new_n1369), .ZN(new_n1370));
  OAI221_X1 g1170(.A(new_n1368), .B1(KEYINPUT127), .B2(new_n1337), .C1(new_n1367), .C2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1337), .A2(KEYINPUT127), .ZN(new_n1372));
  XNOR2_X1  g1172(.A(new_n1320), .B(new_n1372), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1371), .B(new_n1373), .ZN(G402));
endmodule


