//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT73), .ZN(new_n209));
  AND2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT73), .A3(new_n202), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n208), .A2(new_n212), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n210), .A2(new_n211), .ZN(new_n218));
  AND2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n218), .A2(new_n221), .A3(KEYINPUT73), .A4(new_n203), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G127gat), .B(G134gat), .Z(new_n226));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(G113gat), .B(G120gat), .Z(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n222), .A3(KEYINPUT3), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n225), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n228), .A2(new_n232), .A3(KEYINPUT69), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT69), .B1(new_n228), .B2(new_n232), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n217), .A2(new_n222), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n232), .A3(new_n228), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n245), .A2(new_n238), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n237), .A2(new_n243), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(KEYINPUT4), .B(new_n223), .C1(new_n239), .C2(new_n240), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n238), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n248), .A2(new_n235), .A3(new_n249), .A4(new_n236), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n233), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n245), .ZN(new_n252));
  INV_X1    g051(.A(new_n236), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n244), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT0), .ZN(new_n258));
  XNOR2_X1  g057(.A(G57gat), .B(G85gat), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT6), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n255), .A3(new_n260), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n256), .A2(KEYINPUT6), .A3(new_n261), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT22), .ZN(new_n272));
  INV_X1    g071(.A(G211gat), .ZN(new_n273));
  INV_X1    g072(.A(G218gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n271), .A3(new_n275), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT26), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n285), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT27), .B(G183gat), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT28), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n296), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n294), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n302), .B(new_n303), .C1(G169gat), .C2(G176gat), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT23), .B1(new_n286), .B2(KEYINPUT65), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307));
  INV_X1    g106(.A(G183gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n296), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT67), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n311), .A3(new_n284), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n310), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n307), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n313), .A3(new_n307), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n306), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n293), .A2(new_n304), .A3(new_n305), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n285), .A2(KEYINPUT24), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n309), .A2(KEYINPUT64), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n284), .A2(new_n310), .ZN(new_n321));
  OR3_X1    g120(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT25), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n301), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n283), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n316), .ZN(new_n328));
  OAI211_X1 g127(.A(KEYINPUT25), .B(new_n318), .C1(new_n328), .C2(new_n314), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  INV_X1    g129(.A(new_n323), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n293), .A2(new_n304), .A3(new_n305), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n282), .B1(new_n334), .B2(new_n301), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n281), .B1(new_n327), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n298), .B(new_n299), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n329), .A2(new_n333), .B1(new_n337), .B2(new_n294), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n282), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n339));
  INV_X1    g138(.A(new_n281), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n283), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n270), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n342), .A3(new_n270), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n345), .B2(KEYINPUT30), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT72), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(KEYINPUT72), .A3(new_n347), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n267), .B(new_n346), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT81), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n279), .B2(new_n280), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n242), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n354));
  AND2_X1   g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT3), .B1(new_n217), .B2(new_n222), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n281), .B1(new_n356), .B2(KEYINPUT29), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n354), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n357), .A2(new_n358), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n354), .B2(new_n357), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n362));
  OAI22_X1  g161(.A1(new_n359), .A2(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n361), .A2(new_n362), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G22gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT31), .B(G50gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  NOR3_X1   g168(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT76), .B(G22gat), .Z(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(new_n363), .B2(new_n364), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n369), .A2(KEYINPUT77), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n365), .A2(new_n371), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n365), .A2(new_n371), .A3(new_n374), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n370), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT70), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(G15gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G43gat), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n239), .A2(new_n240), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n325), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n334), .A2(new_n241), .A3(new_n301), .ZN(new_n386));
  INV_X1    g185(.A(G227gat), .ZN(new_n387));
  INV_X1    g186(.A(G233gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n383), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(KEYINPUT32), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n390), .B(KEYINPUT32), .C1(new_n383), .C2(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT34), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n385), .A2(new_n386), .ZN(new_n398));
  INV_X1    g197(.A(new_n389), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT34), .B(new_n389), .C1(new_n385), .C2(new_n386), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n394), .A3(new_n395), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(KEYINPUT35), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n352), .A2(new_n379), .A3(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n351), .A2(KEYINPUT81), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n351), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT71), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n402), .A2(new_n394), .A3(new_n395), .ZN(new_n413));
  INV_X1    g212(.A(new_n400), .ZN(new_n414));
  INV_X1    g213(.A(new_n401), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n394), .A2(new_n395), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n396), .A2(KEYINPUT71), .A3(new_n402), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n411), .A2(new_n417), .A3(new_n418), .A4(new_n379), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT35), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT36), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n406), .A2(KEYINPUT36), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n427));
  OR3_X1    g226(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n363), .A2(new_n364), .A3(new_n372), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n373), .B2(new_n374), .ZN(new_n430));
  INV_X1    g229(.A(new_n378), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT78), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n427), .A2(new_n434), .A3(new_n351), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n336), .A2(new_n342), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n270), .B1(new_n436), .B2(KEYINPUT37), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT79), .B(KEYINPUT38), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n336), .A2(new_n342), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(new_n266), .A3(new_n265), .A4(new_n344), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n443), .B(new_n438), .C1(new_n437), .C2(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n436), .A2(KEYINPUT37), .ZN(new_n445));
  INV_X1    g244(.A(new_n270), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n440), .ZN(new_n447));
  INV_X1    g246(.A(new_n438), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT80), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n442), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n436), .A2(new_n446), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n347), .B2(new_n344), .ZN(new_n452));
  INV_X1    g251(.A(new_n348), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(new_n349), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n243), .A2(new_n235), .A3(new_n246), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT39), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n253), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n260), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n251), .A2(new_n236), .A3(new_n245), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT39), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n456), .B2(new_n253), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n455), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n462), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(KEYINPUT40), .A3(new_n260), .A4(new_n458), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n465), .A3(new_n262), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n379), .B1(new_n454), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n435), .B1(new_n450), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n421), .B1(new_n426), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G113gat), .B(G141gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT82), .B(G197gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT11), .B(G169gat), .Z(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT12), .ZN(new_n475));
  NAND2_X1  g274(.A1(G229gat), .A2(G233gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(KEYINPUT13), .Z(new_n477));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n478));
  INV_X1    g277(.A(G43gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G50gat), .ZN(new_n480));
  INV_X1    g279(.A(G50gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G43gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n482), .A3(KEYINPUT15), .ZN(new_n483));
  NAND2_X1  g282(.A1(G29gat), .A2(G36gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G29gat), .ZN(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT14), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(G29gat), .B2(G36gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n485), .B1(new_n491), .B2(KEYINPUT83), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT83), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n483), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(KEYINPUT85), .A2(G29gat), .A3(G36gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n499), .A2(new_n483), .A3(new_n490), .A4(new_n488), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n479), .A2(KEYINPUT84), .A3(G50gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n504));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n478), .B1(new_n495), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n480), .A2(new_n482), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n502), .B(new_n501), .C1(new_n509), .C2(KEYINPUT84), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n484), .A2(new_n511), .ZN(new_n512));
  AND4_X1   g311(.A1(new_n490), .A2(new_n488), .A3(new_n512), .A4(new_n496), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n513), .A3(new_n483), .ZN(new_n514));
  INV_X1    g313(.A(new_n494), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n493), .B1(new_n488), .B2(new_n490), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n515), .A2(new_n516), .A3(new_n485), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n514), .B(KEYINPUT86), .C1(new_n517), .C2(new_n483), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n508), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT16), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(G1gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n523), .B(new_n524), .C1(G1gat), .C2(new_n521), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G8gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(new_n519), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n477), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n508), .A2(new_n532), .A3(new_n518), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n508), .A2(new_n518), .A3(KEYINPUT87), .A4(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n495), .A2(new_n507), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT89), .B1(new_n538), .B2(KEYINPUT17), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n540));
  NOR4_X1   g339(.A1(new_n495), .A2(new_n507), .A3(new_n540), .A4(new_n532), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n528), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n529), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n476), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n531), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n476), .A4(new_n544), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n475), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n548), .A3(new_n475), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n469), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(KEYINPUT41), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT94), .ZN(new_n557));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT95), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566));
  NAND3_X1  g365(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT96), .B1(new_n563), .B2(KEYINPUT7), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n574), .B1(new_n567), .B2(new_n565), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n561), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n565), .A2(new_n567), .ZN(new_n577));
  INV_X1    g376(.A(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n561), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n568), .A4(new_n572), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(KEYINPUT97), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n573), .A2(new_n575), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n537), .A2(new_n542), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G190gat), .B(G218gat), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n520), .A2(new_n586), .B1(KEYINPUT41), .B2(new_n555), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n590), .B1(new_n588), .B2(new_n591), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n560), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n559), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G71gat), .B(G78gat), .Z(new_n599));
  XNOR2_X1  g398(.A(G57gat), .B(G64gat), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n600), .A2(KEYINPUT90), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT9), .ZN(new_n602));
  INV_X1    g401(.A(G71gat), .ZN(new_n603));
  INV_X1    g402(.A(G78gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n600), .B2(KEYINPUT90), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n599), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G64gat), .ZN(new_n608));
  OR3_X1    g407(.A1(new_n608), .A2(KEYINPUT91), .A3(G57gat), .ZN(new_n609));
  INV_X1    g408(.A(G57gat), .ZN(new_n610));
  OR3_X1    g409(.A1(new_n610), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT91), .B1(new_n608), .B2(G57gat), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT92), .B1(new_n610), .B2(G64gat), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n609), .A2(new_n611), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n599), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n605), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n582), .A2(new_n617), .A3(new_n585), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n576), .A2(new_n581), .A3(new_n607), .A4(new_n616), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n586), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n618), .A2(new_n620), .ZN(new_n627));
  INV_X1    g426(.A(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(G231gat), .B(G233gat), .C1(new_n622), .C2(KEYINPUT21), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT21), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n617), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G127gat), .ZN(new_n645));
  INV_X1    g444(.A(G127gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n526), .B1(KEYINPUT21), .B2(new_n622), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n651), .A3(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT93), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G155gat), .ZN(new_n656));
  XOR2_X1   g455(.A(G183gat), .B(G211gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n650), .A2(new_n652), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n598), .A2(new_n639), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n553), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n267), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT98), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT98), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g472(.A(new_n346), .B1(new_n350), .B2(new_n348), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n675), .A2(G8gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(KEYINPUT42), .B2(new_n678), .ZN(G1325gat));
  AOI21_X1  g479(.A(new_n424), .B1(new_n422), .B2(KEYINPUT36), .ZN(new_n681));
  OAI21_X1  g480(.A(G15gat), .B1(new_n665), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n406), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n665), .B2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n433), .B(new_n370), .C1(new_n377), .C2(new_n378), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n665), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NOR3_X1   g490(.A1(new_n598), .A2(new_n662), .A3(new_n638), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n553), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n486), .A3(new_n671), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n408), .A2(new_n409), .B1(new_n419), .B2(KEYINPUT35), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT101), .B1(new_n468), .B2(new_n426), .ZN(new_n699));
  INV_X1    g498(.A(new_n440), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n439), .B1(new_n336), .B2(new_n342), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n700), .A2(new_n701), .A3(new_n270), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n443), .B1(new_n702), .B2(new_n438), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n267), .A2(new_n345), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n447), .A2(KEYINPUT80), .A3(new_n448), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n441), .ZN(new_n706));
  INV_X1    g505(.A(new_n466), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n432), .B1(new_n674), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n681), .A3(new_n710), .A4(new_n435), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n698), .B1(new_n699), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n697), .B1(new_n712), .B2(new_n598), .ZN(new_n713));
  INV_X1    g512(.A(new_n598), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n469), .A2(KEYINPUT44), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n638), .B(KEYINPUT100), .Z(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n552), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n662), .B(KEYINPUT99), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n722), .B2(new_n670), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n696), .A2(new_n723), .ZN(G1328gat));
  NOR3_X1   g523(.A1(new_n693), .A2(G36gat), .A3(new_n454), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT46), .ZN(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n722), .B2(new_n454), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1329gat));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n715), .A3(new_n426), .A4(new_n721), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G43gat), .ZN(new_n730));
  INV_X1    g529(.A(new_n406), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n479), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n693), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1330gat));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n432), .A3(new_n721), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n687), .A2(new_n481), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT103), .Z(new_n741));
  AOI21_X1  g540(.A(new_n739), .B1(new_n694), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n737), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n738), .B1(new_n737), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n716), .A2(new_n687), .A3(new_n721), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n745), .A2(G50gat), .B1(new_n694), .B2(new_n741), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n743), .A2(new_n744), .B1(new_n746), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI22_X1  g546(.A1(new_n687), .A2(new_n351), .B1(new_n706), .B2(new_n708), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n710), .B1(new_n748), .B2(new_n681), .ZN(new_n749));
  AND4_X1   g548(.A1(new_n710), .A2(new_n709), .A3(new_n681), .A4(new_n435), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n421), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n662), .ZN(new_n752));
  NOR4_X1   g551(.A1(new_n717), .A2(new_n714), .A3(new_n552), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n670), .B(KEYINPUT105), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(new_n610), .ZN(G1332gat));
  INV_X1    g556(.A(new_n754), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n454), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1333gat));
  NOR3_X1   g563(.A1(new_n754), .A2(G71gat), .A3(new_n406), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n758), .A2(new_n426), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(G71gat), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n754), .A2(new_n688), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n604), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n552), .A2(new_n662), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n638), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT108), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n716), .A2(new_n671), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n570), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n775), .B2(new_n774), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n699), .A2(new_n711), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n598), .B1(new_n778), .B2(new_n421), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT51), .B1(new_n779), .B2(new_n771), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  INV_X1    g580(.A(new_n771), .ZN(new_n782));
  NOR4_X1   g581(.A1(new_n712), .A2(new_n781), .A3(new_n598), .A4(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT110), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n751), .A2(new_n714), .A3(new_n771), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n781), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n779), .A2(KEYINPUT51), .A3(new_n771), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n790), .A2(new_n570), .A3(new_n638), .A4(new_n671), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n777), .A2(new_n791), .ZN(G1336gat));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n713), .A2(new_n715), .A3(new_n674), .A4(new_n773), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n718), .B1(new_n780), .B2(new_n783), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n674), .A2(new_n571), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n797), .B(new_n800), .ZN(G1337gat));
  XOR2_X1   g600(.A(KEYINPUT112), .B(G99gat), .Z(new_n802));
  NOR2_X1   g601(.A1(new_n639), .A2(new_n406), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n790), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n716), .A2(new_n773), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n426), .A2(new_n802), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT113), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  INV_X1    g608(.A(new_n803), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n784), .B2(new_n789), .ZN(new_n811));
  OAI221_X1 g610(.A(new_n809), .B1(new_n805), .B2(new_n806), .C1(new_n811), .C2(new_n802), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(G1338gat));
  OR2_X1    g612(.A1(new_n379), .A2(G106gat), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n798), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G106gat), .B1(new_n805), .B2(new_n379), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G106gat), .B1(new_n805), .B2(new_n688), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n817), .ZN(G1339gat));
  NOR2_X1   g620(.A1(new_n552), .A2(new_n663), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n628), .B1(new_n621), .B2(new_n623), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n633), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n621), .A2(new_n623), .A3(new_n628), .ZN(new_n827));
  AND4_X1   g626(.A1(new_n826), .A2(new_n626), .A3(KEYINPUT54), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n824), .B1(new_n624), .B2(new_n625), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n829), .B2(new_n827), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n825), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n626), .A2(KEYINPUT54), .A3(new_n827), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n829), .A2(new_n826), .A3(new_n827), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n825), .A2(KEYINPUT55), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n635), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n545), .A2(new_n546), .ZN(new_n840));
  AND4_X1   g639(.A1(new_n548), .A2(new_n840), .A3(new_n530), .A4(new_n475), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n833), .B(new_n839), .C1(new_n841), .C2(new_n549), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n476), .B1(new_n543), .B2(new_n544), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n527), .A2(new_n529), .A3(new_n477), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n474), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT115), .B(new_n474), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n551), .A2(new_n847), .A3(new_n638), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n714), .B1(new_n842), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n551), .A2(new_n847), .A3(new_n848), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n838), .B1(new_n828), .B2(new_n830), .ZN(new_n852));
  INV_X1    g651(.A(new_n825), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n835), .B2(new_n836), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n852), .B(new_n636), .C1(new_n854), .C2(KEYINPUT55), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n851), .A2(new_n855), .A3(new_n598), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n720), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT116), .B1(new_n850), .B2(new_n856), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n822), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n417), .A2(new_n418), .A3(new_n379), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n861), .A2(new_n674), .A3(new_n862), .A4(new_n755), .ZN(new_n863));
  AOI21_X1  g662(.A(G113gat), .B1(new_n863), .B2(new_n552), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n842), .A2(new_n849), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n598), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n851), .A2(new_n855), .A3(new_n598), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n720), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n860), .ZN(new_n870));
  INV_X1    g669(.A(new_n822), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n872), .B2(new_n688), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n874), .B(new_n687), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n670), .A2(new_n674), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n876), .A2(new_n406), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n552), .A2(G113gat), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n864), .B1(new_n879), .B2(new_n880), .ZN(G1340gat));
  AOI21_X1  g680(.A(G120gat), .B1(new_n863), .B2(new_n638), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n718), .A2(G120gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n879), .B2(new_n883), .ZN(G1341gat));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n646), .A3(new_n662), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n879), .A2(new_n720), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n646), .ZN(G1342gat));
  INV_X1    g686(.A(G134gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n863), .A2(new_n888), .A3(new_n714), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT56), .Z(new_n890));
  NAND2_X1  g689(.A1(new_n879), .A2(new_n714), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G134gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1343gat));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n426), .ZN(new_n894));
  XNOR2_X1  g693(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n872), .B2(new_n432), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n688), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n831), .A2(new_n900), .A3(new_n832), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n901), .B(new_n839), .C1(new_n841), .C2(new_n549), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n831), .B2(new_n832), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n849), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n598), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n662), .B1(new_n905), .B2(new_n867), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n899), .B1(new_n906), .B2(new_n822), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n894), .B1(new_n897), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G141gat), .B1(new_n909), .B2(new_n719), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n861), .A2(new_n755), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n681), .A2(new_n432), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n674), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n552), .A2(new_n204), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT58), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n910), .B(new_n919), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1344gat));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n379), .B1(new_n870), .B2(new_n871), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n822), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT122), .B1(new_n552), .B2(new_n663), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n687), .B1(new_n906), .B2(new_n927), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n923), .A2(new_n896), .B1(new_n928), .B2(new_n898), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n894), .A2(new_n638), .ZN(new_n930));
  OAI21_X1  g729(.A(G148gat), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g730(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n932));
  OAI211_X1 g731(.A(new_n638), .B(new_n894), .C1(new_n897), .C2(new_n908), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n205), .A2(KEYINPUT59), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n931), .A2(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n755), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n639), .A2(G148gat), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n872), .A2(new_n936), .A3(new_n914), .A4(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT120), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n922), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n933), .A2(new_n934), .ZN(new_n942));
  INV_X1    g741(.A(new_n932), .ZN(new_n943));
  AOI211_X1 g742(.A(new_n379), .B(new_n895), .C1(new_n870), .C2(new_n871), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n856), .B1(new_n904), .B2(new_n598), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n926), .B(new_n925), .C1(new_n945), .C2(new_n662), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT57), .B1(new_n946), .B2(new_n687), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n638), .B(new_n894), .C1(new_n944), .C2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n943), .B1(new_n948), .B2(G148gat), .ZN(new_n949));
  OAI211_X1 g748(.A(KEYINPUT123), .B(new_n939), .C1(new_n942), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n941), .A2(new_n950), .ZN(G1345gat));
  OAI21_X1  g750(.A(G155gat), .B1(new_n909), .B2(new_n869), .ZN(new_n952));
  INV_X1    g751(.A(new_n915), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n213), .A3(new_n662), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1346gat));
  OAI21_X1  g754(.A(G162gat), .B1(new_n909), .B2(new_n598), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n214), .A3(new_n714), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1347gat));
  NOR2_X1   g757(.A1(new_n861), .A2(new_n671), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n862), .A2(new_n454), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(G169gat), .B1(new_n962), .B2(new_n552), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n755), .A2(new_n731), .A3(new_n674), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n874), .B1(new_n861), .B2(new_n687), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n872), .A2(KEYINPUT117), .A3(new_n688), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n719), .A2(new_n289), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(G1348gat));
  INV_X1    g768(.A(new_n964), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n717), .A2(new_n290), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n970), .B(new_n971), .C1(new_n873), .C2(new_n875), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n965), .A2(new_n966), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n970), .A4(new_n971), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n290), .B1(new_n961), .B2(new_n639), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT125), .A4(new_n977), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1349gat));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n962), .A2(new_n295), .A3(new_n662), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n308), .B1(new_n967), .B2(new_n720), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n983), .B(KEYINPUT60), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n983), .A2(KEYINPUT60), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n962), .A2(new_n295), .A3(new_n662), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n876), .A2(new_n869), .A3(new_n964), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n987), .B(new_n988), .C1(new_n989), .C2(new_n308), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n986), .A2(new_n990), .ZN(G1350gat));
  NAND3_X1  g790(.A1(new_n962), .A2(new_n296), .A3(new_n714), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n967), .A2(new_n714), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n993), .B1(new_n994), .B2(G190gat), .ZN(new_n995));
  AOI211_X1 g794(.A(KEYINPUT61), .B(new_n296), .C1(new_n967), .C2(new_n714), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G1351gat));
  NOR4_X1   g796(.A1(new_n861), .A2(new_n454), .A3(new_n671), .A4(new_n913), .ZN(new_n998));
  XOR2_X1   g797(.A(KEYINPUT127), .B(G197gat), .Z(new_n999));
  NAND3_X1  g798(.A1(new_n998), .A2(new_n552), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(new_n929), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n936), .A2(new_n426), .A3(new_n454), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1003), .A2(new_n719), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1000), .B1(new_n1004), .B2(new_n999), .ZN(G1352gat));
  INV_X1    g804(.A(G204gat), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n998), .A2(new_n1006), .A3(new_n638), .ZN(new_n1007));
  XOR2_X1   g806(.A(new_n1007), .B(KEYINPUT62), .Z(new_n1008));
  OAI21_X1  g807(.A(G204gat), .B1(new_n1003), .B2(new_n717), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(G1353gat));
  NAND3_X1  g809(.A1(new_n998), .A2(new_n273), .A3(new_n662), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1001), .A2(new_n662), .A3(new_n1002), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n1012), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1013));
  AOI21_X1  g812(.A(KEYINPUT63), .B1(new_n1012), .B2(G211gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(G1354gat));
  OAI21_X1  g814(.A(G218gat), .B1(new_n1003), .B2(new_n598), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n274), .A3(new_n714), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1016), .A2(new_n1017), .ZN(G1355gat));
endmodule


