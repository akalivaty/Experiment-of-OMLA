

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764;

  AND2_X1 U377 ( .A1(n360), .A2(n359), .ZN(n753) );
  INV_X1 U378 ( .A(n622), .ZN(n359) );
  XNOR2_X1 U379 ( .A(n411), .B(n361), .ZN(n360) );
  INV_X1 U380 ( .A(KEYINPUT48), .ZN(n361) );
  NOR2_X1 U381 ( .A1(n356), .A2(n387), .ZN(n413) );
  NOR2_X1 U382 ( .A1(n616), .A2(n605), .ZN(n606) );
  XNOR2_X1 U383 ( .A(n558), .B(KEYINPUT106), .ZN(n600) );
  XNOR2_X1 U384 ( .A(n528), .B(n527), .ZN(n553) );
  XNOR2_X1 U385 ( .A(n358), .B(n523), .ZN(n373) );
  XNOR2_X1 U386 ( .A(n522), .B(n517), .ZN(n358) );
  XOR2_X1 U387 ( .A(KEYINPUT67), .B(G131), .Z(n519) );
  XOR2_X1 U388 ( .A(G125), .B(G146), .Z(n477) );
  NAND2_X1 U389 ( .A1(n384), .A2(n357), .ZN(n356) );
  INV_X1 U390 ( .A(n388), .ZN(n357) );
  NOR2_X1 U391 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U392 ( .A1(n671), .A2(n604), .ZN(n616) );
  AND2_X1 U393 ( .A1(n739), .A2(KEYINPUT2), .ZN(n624) );
  NOR2_X1 U394 ( .A1(n763), .A2(n764), .ZN(n598) );
  XNOR2_X1 U395 ( .A(n393), .B(n392), .ZN(n694) );
  XNOR2_X2 U396 ( .A(n390), .B(n462), .ZN(n680) );
  XNOR2_X1 U397 ( .A(n430), .B(n488), .ZN(n585) );
  AND2_X1 U398 ( .A1(n407), .A2(n567), .ZN(n406) );
  NAND2_X1 U399 ( .A1(n415), .A2(n414), .ZN(n416) );
  NOR2_X1 U400 ( .A1(n694), .A2(n547), .ZN(n500) );
  NOR2_X1 U401 ( .A1(n547), .A2(n533), .ZN(n534) );
  NOR2_X2 U402 ( .A1(n679), .A2(n680), .ZN(n463) );
  XNOR2_X1 U403 ( .A(n409), .B(n504), .ZN(n752) );
  XNOR2_X1 U404 ( .A(n482), .B(n519), .ZN(n409) );
  NOR2_X1 U405 ( .A1(n416), .A2(n569), .ZN(n568) );
  XNOR2_X1 U406 ( .A(n477), .B(n434), .ZN(n515) );
  XNOR2_X1 U407 ( .A(n498), .B(n497), .ZN(n547) );
  XNOR2_X1 U408 ( .A(n752), .B(n449), .ZN(n397) );
  INV_X1 U409 ( .A(G146), .ZN(n449) );
  XNOR2_X1 U410 ( .A(n546), .B(KEYINPUT110), .ZN(n590) );
  BUF_X1 U411 ( .A(n451), .Z(n754) );
  OR2_X1 U412 ( .A1(n374), .A2(KEYINPUT87), .ZN(n380) );
  NAND2_X1 U413 ( .A1(n389), .A2(n584), .ZN(n388) );
  XNOR2_X1 U414 ( .A(n581), .B(KEYINPUT47), .ZN(n385) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n516) );
  OR2_X1 U416 ( .A1(n673), .A2(n600), .ZN(n559) );
  NOR2_X1 U417 ( .A1(n362), .A2(n371), .ZN(n402) );
  INV_X1 U418 ( .A(KEYINPUT90), .ZN(n408) );
  XOR2_X1 U419 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n513) );
  XNOR2_X1 U420 ( .A(KEYINPUT11), .B(KEYINPUT100), .ZN(n512) );
  XNOR2_X1 U421 ( .A(G113), .B(G104), .ZN(n520) );
  INV_X1 U422 ( .A(G237), .ZN(n486) );
  OR2_X1 U423 ( .A1(n695), .A2(n429), .ZN(n428) );
  XNOR2_X1 U424 ( .A(n397), .B(n470), .ZN(n645) );
  XNOR2_X1 U425 ( .A(n443), .B(n368), .ZN(n633) );
  XNOR2_X1 U426 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U427 ( .A(n595), .B(n594), .ZN(n615) );
  NAND2_X1 U428 ( .A1(n610), .A2(n591), .ZN(n595) );
  INV_X1 U429 ( .A(KEYINPUT70), .ZN(n592) );
  AND2_X1 U430 ( .A1(n601), .A2(n682), .ZN(n394) );
  XNOR2_X1 U431 ( .A(n579), .B(n377), .ZN(n376) );
  INV_X1 U432 ( .A(KEYINPUT112), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n396), .B(n395), .ZN(n609) );
  INV_X1 U434 ( .A(KEYINPUT30), .ZN(n395) );
  NAND2_X1 U435 ( .A1(n590), .A2(n695), .ZN(n396) );
  NOR2_X1 U436 ( .A1(G902), .A2(n639), .ZN(n528) );
  AND2_X1 U437 ( .A1(n398), .A2(n390), .ZN(n550) );
  AND2_X1 U438 ( .A1(n562), .A2(n399), .ZN(n398) );
  NAND2_X1 U439 ( .A1(n727), .A2(G217), .ZN(n423) );
  INV_X1 U440 ( .A(n633), .ZN(n422) );
  BUF_X1 U441 ( .A(n727), .Z(n733) );
  XNOR2_X1 U442 ( .A(n397), .B(n459), .ZN(n729) );
  INV_X1 U443 ( .A(KEYINPUT35), .ZN(n391) );
  NAND2_X1 U444 ( .A1(n539), .A2(n541), .ZN(n414) );
  AND2_X1 U445 ( .A1(n374), .A2(KEYINPUT87), .ZN(n382) );
  XNOR2_X1 U446 ( .A(G137), .B(G101), .ZN(n467) );
  XNOR2_X1 U447 ( .A(n418), .B(n417), .ZN(n473) );
  XNOR2_X1 U448 ( .A(G116), .B(G113), .ZN(n418) );
  XNOR2_X1 U449 ( .A(KEYINPUT3), .B(G119), .ZN(n417) );
  XNOR2_X1 U450 ( .A(G128), .B(G119), .ZN(n438) );
  XNOR2_X1 U451 ( .A(KEYINPUT78), .B(KEYINPUT23), .ZN(n436) );
  XOR2_X1 U452 ( .A(G110), .B(KEYINPUT24), .Z(n437) );
  XNOR2_X1 U453 ( .A(n433), .B(n432), .ZN(n505) );
  INV_X1 U454 ( .A(KEYINPUT8), .ZN(n432) );
  XNOR2_X1 U455 ( .A(G143), .B(G128), .ZN(n476) );
  XOR2_X1 U456 ( .A(G137), .B(KEYINPUT68), .Z(n450) );
  XNOR2_X1 U457 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n480) );
  AND2_X1 U458 ( .A1(n609), .A2(n696), .ZN(n591) );
  NOR2_X1 U459 ( .A1(n553), .A2(n556), .ZN(n531) );
  AND2_X1 U460 ( .A1(n603), .A2(n590), .ZN(n577) );
  XNOR2_X1 U461 ( .A(n431), .B(G953), .ZN(n451) );
  INV_X1 U462 ( .A(KEYINPUT64), .ZN(n431) );
  NAND2_X1 U463 ( .A1(n406), .A2(n405), .ZN(n570) );
  NAND2_X1 U464 ( .A1(n403), .A2(n402), .ZN(n405) );
  XNOR2_X1 U465 ( .A(G116), .B(G107), .ZN(n501) );
  XNOR2_X1 U466 ( .A(n476), .B(G134), .ZN(n504) );
  XNOR2_X1 U467 ( .A(n373), .B(n518), .ZN(n639) );
  XOR2_X1 U468 ( .A(n515), .B(n514), .Z(n518) );
  XNOR2_X1 U469 ( .A(G101), .B(KEYINPUT74), .ZN(n455) );
  INV_X1 U470 ( .A(G953), .ZN(n738) );
  INV_X1 U471 ( .A(KEYINPUT33), .ZN(n392) );
  NAND2_X1 U472 ( .A1(n425), .A2(n424), .ZN(n580) );
  AND2_X1 U473 ( .A1(n426), .A2(n428), .ZN(n425) );
  NAND2_X1 U474 ( .A1(n645), .A2(n487), .ZN(n378) );
  OR2_X1 U475 ( .A1(n633), .A2(G902), .ZN(n400) );
  XNOR2_X1 U476 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n444) );
  INV_X1 U477 ( .A(n714), .ZN(n375) );
  XNOR2_X1 U478 ( .A(n597), .B(n596), .ZN(n763) );
  INV_X1 U479 ( .A(KEYINPUT40), .ZN(n596) );
  BUF_X1 U480 ( .A(n680), .Z(n374) );
  AND2_X1 U481 ( .A1(n376), .A2(n580), .ZN(n669) );
  OR2_X1 U482 ( .A1(n620), .A2(n613), .ZN(n637) );
  XOR2_X1 U483 ( .A(n555), .B(KEYINPUT107), .Z(n673) );
  XNOR2_X1 U484 ( .A(n600), .B(n599), .ZN(n671) );
  INV_X1 U485 ( .A(KEYINPUT111), .ZN(n599) );
  INV_X1 U486 ( .A(KEYINPUT122), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n421) );
  XNOR2_X1 U488 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U489 ( .A(n404), .B(n762), .ZN(G24) );
  INV_X1 U490 ( .A(n414), .ZN(n634) );
  AND2_X1 U491 ( .A1(n568), .A2(n408), .ZN(n362) );
  AND2_X1 U492 ( .A1(n414), .A2(n372), .ZN(n363) );
  INV_X1 U493 ( .A(n683), .ZN(n399) );
  AND2_X1 U494 ( .A1(n376), .A2(n375), .ZN(n364) );
  XNOR2_X1 U495 ( .A(n511), .B(n510), .ZN(n556) );
  INV_X1 U496 ( .A(n556), .ZN(n554) );
  XOR2_X1 U497 ( .A(n446), .B(n444), .Z(n365) );
  AND2_X1 U498 ( .A1(n608), .A2(KEYINPUT83), .ZN(n366) );
  XNOR2_X1 U499 ( .A(n546), .B(KEYINPUT6), .ZN(n601) );
  NAND2_X1 U500 ( .A1(n545), .A2(KEYINPUT90), .ZN(n367) );
  AND2_X1 U501 ( .A1(n505), .A2(G221), .ZN(n368) );
  AND2_X1 U502 ( .A1(n695), .A2(n429), .ZN(n369) );
  NOR2_X1 U503 ( .A1(n607), .A2(n374), .ZN(n370) );
  XNOR2_X1 U504 ( .A(n515), .B(n435), .ZN(n751) );
  AND2_X1 U505 ( .A1(n569), .A2(KEYINPUT90), .ZN(n371) );
  OR2_X1 U506 ( .A1(KEYINPUT44), .A2(KEYINPUT91), .ZN(n372) );
  OR2_X1 U507 ( .A1(n754), .A2(G952), .ZN(n655) );
  INV_X1 U508 ( .A(n553), .ZN(n557) );
  AND2_X1 U509 ( .A1(n553), .A2(n554), .ZN(n558) );
  NOR2_X1 U510 ( .A1(n366), .A2(n614), .ZN(n389) );
  XNOR2_X2 U511 ( .A(n378), .B(n471), .ZN(n546) );
  NAND2_X1 U512 ( .A1(n381), .A2(n379), .ZN(n387) );
  OR2_X1 U513 ( .A1(n607), .A2(n380), .ZN(n379) );
  NOR2_X1 U514 ( .A1(n383), .A2(n382), .ZN(n381) );
  AND2_X1 U515 ( .A1(n607), .A2(KEYINPUT87), .ZN(n383) );
  NAND2_X1 U516 ( .A1(n385), .A2(n582), .ZN(n384) );
  NAND2_X1 U517 ( .A1(n578), .A2(n390), .ZN(n579) );
  XNOR2_X2 U518 ( .A(n461), .B(n460), .ZN(n390) );
  XNOR2_X2 U519 ( .A(n530), .B(n391), .ZN(n404) );
  NAND2_X1 U520 ( .A1(n401), .A2(n602), .ZN(n393) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT72), .ZN(n401) );
  NAND2_X1 U522 ( .A1(n535), .A2(n394), .ZN(n536) );
  INV_X1 U523 ( .A(n415), .ZN(n636) );
  XNOR2_X2 U524 ( .A(n538), .B(KEYINPUT32), .ZN(n415) );
  INV_X1 U525 ( .A(n562), .ZN(n682) );
  XNOR2_X2 U526 ( .A(n400), .B(n365), .ZN(n562) );
  XNOR2_X1 U527 ( .A(n534), .B(KEYINPUT22), .ZN(n539) );
  AND2_X1 U528 ( .A1(n401), .A2(n546), .ZN(n690) );
  NAND2_X1 U529 ( .A1(n404), .A2(n568), .ZN(n403) );
  NAND2_X1 U530 ( .A1(n404), .A2(n367), .ZN(n407) );
  XNOR2_X2 U531 ( .A(n410), .B(KEYINPUT4), .ZN(n482) );
  XNOR2_X2 U532 ( .A(KEYINPUT65), .B(KEYINPUT66), .ZN(n410) );
  NAND2_X1 U533 ( .A1(n413), .A2(n412), .ZN(n411) );
  XNOR2_X1 U534 ( .A(n598), .B(KEYINPUT46), .ZN(n412) );
  NAND2_X1 U535 ( .A1(n363), .A2(n415), .ZN(n544) );
  NAND2_X1 U536 ( .A1(n416), .A2(n542), .ZN(n543) );
  XNOR2_X1 U537 ( .A(n420), .B(n419), .ZN(G66) );
  NAND2_X1 U538 ( .A1(n421), .A2(n655), .ZN(n420) );
  NAND2_X1 U539 ( .A1(n427), .A2(n369), .ZN(n424) );
  INV_X1 U540 ( .A(n585), .ZN(n427) );
  NAND2_X1 U541 ( .A1(n585), .A2(n491), .ZN(n426) );
  NAND2_X1 U542 ( .A1(n427), .A2(n695), .ZN(n605) );
  INV_X1 U543 ( .A(n491), .ZN(n429) );
  NAND2_X1 U544 ( .A1(n652), .A2(n628), .ZN(n430) );
  BUF_X1 U545 ( .A(n585), .Z(n620) );
  XNOR2_X1 U546 ( .A(KEYINPUT10), .B(G140), .ZN(n434) );
  INV_X1 U547 ( .A(n450), .ZN(n435) );
  INV_X1 U548 ( .A(G475), .ZN(n525) );
  XNOR2_X1 U549 ( .A(KEYINPUT105), .B(G478), .ZN(n510) );
  XNOR2_X1 U550 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U551 ( .A(n593), .B(n592), .ZN(n594) );
  NAND2_X1 U552 ( .A1(n451), .A2(G234), .ZN(n433) );
  XNOR2_X1 U553 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U554 ( .A(KEYINPUT95), .B(KEYINPUT69), .Z(n439) );
  XNOR2_X1 U555 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U556 ( .A(n751), .B(n442), .ZN(n443) );
  XNOR2_X1 U557 ( .A(G902), .B(KEYINPUT15), .ZN(n628) );
  NAND2_X1 U558 ( .A1(G234), .A2(n628), .ZN(n445) );
  XNOR2_X1 U559 ( .A(KEYINPUT20), .B(n445), .ZN(n447) );
  NAND2_X1 U560 ( .A1(G217), .A2(n447), .ZN(n446) );
  NAND2_X1 U561 ( .A1(n447), .A2(G221), .ZN(n448) );
  XNOR2_X1 U562 ( .A(n448), .B(KEYINPUT21), .ZN(n683) );
  NAND2_X1 U563 ( .A1(n562), .A2(n399), .ZN(n679) );
  XOR2_X1 U564 ( .A(n450), .B(G140), .Z(n453) );
  NAND2_X1 U565 ( .A1(G227), .A2(n754), .ZN(n452) );
  XNOR2_X1 U566 ( .A(n453), .B(n452), .ZN(n458) );
  XNOR2_X1 U567 ( .A(G107), .B(G104), .ZN(n454) );
  XNOR2_X1 U568 ( .A(n454), .B(G110), .ZN(n456) );
  XNOR2_X1 U569 ( .A(n456), .B(n455), .ZN(n474) );
  INV_X1 U570 ( .A(n474), .ZN(n457) );
  XNOR2_X1 U571 ( .A(n458), .B(n457), .ZN(n459) );
  NOR2_X1 U572 ( .A1(n729), .A2(G902), .ZN(n461) );
  INV_X1 U573 ( .A(G469), .ZN(n460) );
  INV_X1 U574 ( .A(KEYINPUT1), .ZN(n462) );
  XOR2_X1 U575 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n465) );
  NAND2_X1 U576 ( .A1(n516), .A2(G210), .ZN(n464) );
  XNOR2_X1 U577 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U578 ( .A(n466), .B(KEYINPUT73), .Z(n469) );
  XNOR2_X1 U579 ( .A(n473), .B(n467), .ZN(n468) );
  XNOR2_X1 U580 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U581 ( .A(G902), .ZN(n487) );
  XOR2_X1 U582 ( .A(KEYINPUT71), .B(G472), .Z(n471) );
  XNOR2_X1 U583 ( .A(KEYINPUT16), .B(G122), .ZN(n472) );
  XNOR2_X1 U584 ( .A(n473), .B(n472), .ZN(n475) );
  XNOR2_X1 U585 ( .A(n475), .B(n474), .ZN(n745) );
  NAND2_X1 U586 ( .A1(n754), .A2(G224), .ZN(n479) );
  XNOR2_X1 U587 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U588 ( .A(n479), .B(n478), .ZN(n484) );
  XNOR2_X1 U589 ( .A(n480), .B(KEYINPUT79), .ZN(n481) );
  XNOR2_X1 U590 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U591 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U592 ( .A(n745), .B(n485), .ZN(n652) );
  NAND2_X1 U593 ( .A1(n487), .A2(n486), .ZN(n489) );
  NAND2_X1 U594 ( .A1(n489), .A2(G210), .ZN(n488) );
  NAND2_X1 U595 ( .A1(n489), .A2(G214), .ZN(n695) );
  INV_X1 U596 ( .A(KEYINPUT77), .ZN(n490) );
  XNOR2_X1 U597 ( .A(n490), .B(KEYINPUT19), .ZN(n491) );
  XNOR2_X1 U598 ( .A(G898), .B(KEYINPUT94), .ZN(n741) );
  NOR2_X1 U599 ( .A1(n738), .A2(n741), .ZN(n746) );
  NAND2_X1 U600 ( .A1(n746), .A2(G902), .ZN(n492) );
  NAND2_X1 U601 ( .A1(n738), .A2(G952), .ZN(n572) );
  NAND2_X1 U602 ( .A1(n492), .A2(n572), .ZN(n495) );
  NAND2_X1 U603 ( .A1(G237), .A2(G234), .ZN(n494) );
  INV_X1 U604 ( .A(KEYINPUT14), .ZN(n493) );
  XNOR2_X1 U605 ( .A(n494), .B(n493), .ZN(n710) );
  INV_X1 U606 ( .A(n710), .ZN(n575) );
  AND2_X1 U607 ( .A1(n495), .A2(n575), .ZN(n496) );
  NAND2_X1 U608 ( .A1(n580), .A2(n496), .ZN(n498) );
  XNOR2_X1 U609 ( .A(KEYINPUT92), .B(KEYINPUT0), .ZN(n497) );
  XNOR2_X1 U610 ( .A(KEYINPUT34), .B(KEYINPUT80), .ZN(n499) );
  XNOR2_X1 U611 ( .A(n500), .B(n499), .ZN(n529) );
  XOR2_X1 U612 ( .A(KEYINPUT104), .B(G122), .Z(n502) );
  XNOR2_X1 U613 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U614 ( .A(n504), .B(n503), .ZN(n509) );
  XOR2_X1 U615 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n507) );
  NAND2_X1 U616 ( .A1(n505), .A2(G217), .ZN(n506) );
  XNOR2_X1 U617 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U618 ( .A(n509), .B(n508), .ZN(n734) );
  NOR2_X1 U619 ( .A1(G902), .A2(n734), .ZN(n511) );
  XNOR2_X1 U620 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U621 ( .A1(G214), .A2(n516), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n519), .B(KEYINPUT101), .ZN(n523) );
  XOR2_X1 U623 ( .A(G143), .B(G122), .Z(n521) );
  XNOR2_X1 U624 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U625 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n526) );
  NOR2_X1 U626 ( .A1(n554), .A2(n557), .ZN(n611) );
  NAND2_X1 U627 ( .A1(n529), .A2(n611), .ZN(n530) );
  XNOR2_X1 U628 ( .A(n531), .B(KEYINPUT109), .ZN(n699) );
  INV_X1 U629 ( .A(n699), .ZN(n532) );
  NAND2_X1 U630 ( .A1(n532), .A2(n399), .ZN(n533) );
  INV_X1 U631 ( .A(n680), .ZN(n535) );
  XNOR2_X1 U632 ( .A(n536), .B(KEYINPUT81), .ZN(n537) );
  NAND2_X1 U633 ( .A1(n539), .A2(n537), .ZN(n538) );
  NOR2_X1 U634 ( .A1(n590), .A2(n562), .ZN(n540) );
  AND2_X1 U635 ( .A1(n540), .A2(n374), .ZN(n541) );
  INV_X1 U636 ( .A(KEYINPUT91), .ZN(n542) );
  NAND2_X1 U637 ( .A1(n544), .A2(n543), .ZN(n545) );
  INV_X1 U638 ( .A(n547), .ZN(n551) );
  NAND2_X1 U639 ( .A1(n690), .A2(n551), .ZN(n549) );
  XOR2_X1 U640 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n548) );
  XNOR2_X1 U641 ( .A(n549), .B(n548), .ZN(n674) );
  XNOR2_X1 U642 ( .A(n550), .B(KEYINPUT97), .ZN(n587) );
  NOR2_X1 U643 ( .A1(n587), .A2(n546), .ZN(n552) );
  AND2_X1 U644 ( .A1(n552), .A2(n551), .ZN(n661) );
  OR2_X1 U645 ( .A1(n674), .A2(n661), .ZN(n560) );
  NOR2_X1 U646 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U647 ( .A(n559), .B(KEYINPUT108), .Z(n702) );
  INV_X1 U648 ( .A(n702), .ZN(n608) );
  NAND2_X1 U649 ( .A1(n560), .A2(n608), .ZN(n566) );
  NAND2_X1 U650 ( .A1(n539), .A2(n601), .ZN(n561) );
  XNOR2_X1 U651 ( .A(n561), .B(KEYINPUT89), .ZN(n564) );
  AND2_X1 U652 ( .A1(n374), .A2(n562), .ZN(n563) );
  AND2_X1 U653 ( .A1(n564), .A2(n563), .ZN(n659) );
  INV_X1 U654 ( .A(n659), .ZN(n565) );
  AND2_X1 U655 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U656 ( .A(KEYINPUT44), .ZN(n569) );
  XNOR2_X2 U657 ( .A(n570), .B(KEYINPUT45), .ZN(n739) );
  NOR2_X1 U658 ( .A1(n754), .A2(G900), .ZN(n571) );
  NAND2_X1 U659 ( .A1(G902), .A2(n571), .ZN(n573) );
  NAND2_X1 U660 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U661 ( .A1(n575), .A2(n574), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n682), .A2(n399), .ZN(n576) );
  NOR2_X1 U663 ( .A1(n588), .A2(n576), .ZN(n603) );
  XNOR2_X1 U664 ( .A(n577), .B(KEYINPUT28), .ZN(n578) );
  NAND2_X1 U665 ( .A1(n669), .A2(n608), .ZN(n581) );
  INV_X1 U666 ( .A(KEYINPUT83), .ZN(n582) );
  NAND2_X1 U667 ( .A1(n669), .A2(KEYINPUT47), .ZN(n583) );
  NAND2_X1 U668 ( .A1(n583), .A2(KEYINPUT83), .ZN(n584) );
  XNOR2_X1 U669 ( .A(n620), .B(KEYINPUT38), .ZN(n696) );
  NAND2_X1 U670 ( .A1(n696), .A2(n695), .ZN(n701) );
  NOR2_X1 U671 ( .A1(n699), .A2(n701), .ZN(n586) );
  XNOR2_X1 U672 ( .A(n586), .B(KEYINPUT41), .ZN(n714) );
  XNOR2_X1 U673 ( .A(KEYINPUT42), .B(n364), .ZN(n764) );
  XNOR2_X1 U674 ( .A(n589), .B(KEYINPUT76), .ZN(n610) );
  XOR2_X1 U675 ( .A(KEYINPUT88), .B(KEYINPUT39), .Z(n593) );
  NAND2_X1 U676 ( .A1(n615), .A2(n600), .ZN(n597) );
  INV_X1 U677 ( .A(n601), .ZN(n602) );
  AND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U679 ( .A(KEYINPUT36), .B(n606), .Z(n607) );
  AND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  INV_X1 U682 ( .A(n637), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n673), .ZN(n678) );
  INV_X1 U684 ( .A(n616), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n617), .A2(n695), .ZN(n618) );
  NOR2_X1 U686 ( .A1(n535), .A2(n618), .ZN(n619) );
  XOR2_X1 U687 ( .A(n619), .B(KEYINPUT43), .Z(n621) );
  NAND2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n638) );
  NAND2_X1 U689 ( .A1(n678), .A2(n638), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n624), .A2(n753), .ZN(n625) );
  XNOR2_X2 U691 ( .A(n625), .B(KEYINPUT75), .ZN(n721) );
  INV_X1 U692 ( .A(n628), .ZN(n626) );
  AND2_X1 U693 ( .A1(n739), .A2(n626), .ZN(n627) );
  NAND2_X1 U694 ( .A1(n753), .A2(n627), .ZN(n631) );
  XOR2_X1 U695 ( .A(KEYINPUT85), .B(n628), .Z(n629) );
  INV_X1 U696 ( .A(KEYINPUT2), .ZN(n717) );
  OR2_X1 U697 ( .A1(n629), .A2(n717), .ZN(n630) );
  AND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X4 U699 ( .A1(n721), .A2(n632), .ZN(n727) );
  INV_X1 U700 ( .A(n655), .ZN(n737) );
  XOR2_X1 U701 ( .A(G110), .B(n634), .Z(G12) );
  XNOR2_X1 U702 ( .A(G119), .B(KEYINPUT127), .ZN(n635) );
  XNOR2_X1 U703 ( .A(n636), .B(n635), .ZN(G21) );
  XNOR2_X1 U704 ( .A(n637), .B(G143), .ZN(G45) );
  XNOR2_X1 U705 ( .A(n638), .B(G140), .ZN(G42) );
  NAND2_X1 U706 ( .A1(n727), .A2(G475), .ZN(n641) );
  XNOR2_X1 U707 ( .A(n639), .B(KEYINPUT59), .ZN(n640) );
  XNOR2_X1 U708 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U709 ( .A1(n642), .A2(n655), .ZN(n644) );
  INV_X1 U710 ( .A(KEYINPUT60), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n644), .B(n643), .ZN(G60) );
  NAND2_X1 U712 ( .A1(n727), .A2(G472), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n645), .B(KEYINPUT62), .ZN(n646) );
  XNOR2_X1 U714 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U715 ( .A1(n648), .A2(n655), .ZN(n650) );
  XOR2_X1 U716 ( .A(KEYINPUT93), .B(KEYINPUT63), .Z(n649) );
  XNOR2_X1 U717 ( .A(n650), .B(n649), .ZN(G57) );
  NAND2_X1 U718 ( .A1(n727), .A2(G210), .ZN(n654) );
  XOR2_X1 U719 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n651) );
  XNOR2_X1 U720 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n654), .B(n653), .ZN(n656) );
  NAND2_X1 U722 ( .A1(n656), .A2(n655), .ZN(n658) );
  XOR2_X1 U723 ( .A(KEYINPUT86), .B(KEYINPUT56), .Z(n657) );
  XNOR2_X1 U724 ( .A(n658), .B(n657), .ZN(G51) );
  XOR2_X1 U725 ( .A(G101), .B(n659), .Z(G3) );
  NAND2_X1 U726 ( .A1(n671), .A2(n661), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n660), .B(G104), .ZN(G6) );
  XOR2_X1 U728 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n663) );
  NAND2_X1 U729 ( .A1(n661), .A2(n673), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(G107), .B(n664), .ZN(G9) );
  XOR2_X1 U732 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n666) );
  NAND2_X1 U733 ( .A1(n669), .A2(n673), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U735 ( .A(G128), .B(KEYINPUT113), .Z(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(G30) );
  NAND2_X1 U737 ( .A1(n669), .A2(n671), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n670), .B(G146), .ZN(G48) );
  NAND2_X1 U739 ( .A1(n671), .A2(n674), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n672), .B(G113), .ZN(G15) );
  XOR2_X1 U741 ( .A(G116), .B(KEYINPUT115), .Z(n676) );
  NAND2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n676), .B(n675), .ZN(G18) );
  XNOR2_X1 U744 ( .A(n370), .B(G125), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U746 ( .A(G134), .B(n678), .ZN(G36) );
  XNOR2_X1 U747 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n726) );
  NAND2_X1 U748 ( .A1(n374), .A2(n679), .ZN(n681) );
  XNOR2_X1 U749 ( .A(KEYINPUT50), .B(n681), .ZN(n687) );
  XOR2_X1 U750 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n685) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U754 ( .A1(n546), .A2(n688), .ZN(n689) );
  NOR2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U756 ( .A(n691), .B(KEYINPUT51), .ZN(n692) );
  XNOR2_X1 U757 ( .A(KEYINPUT117), .B(n692), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n714), .A2(n693), .ZN(n707) );
  NOR2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U760 ( .A(n697), .B(KEYINPUT118), .ZN(n698) );
  NOR2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U762 ( .A(KEYINPUT119), .B(n700), .Z(n704) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U765 ( .A1(n694), .A2(n705), .ZN(n706) );
  NOR2_X1 U766 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U767 ( .A(n708), .B(KEYINPUT52), .ZN(n709) );
  NOR2_X1 U768 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U769 ( .A1(n711), .A2(G952), .ZN(n712) );
  XNOR2_X1 U770 ( .A(n712), .B(KEYINPUT120), .ZN(n713) );
  NAND2_X1 U771 ( .A1(n713), .A2(n738), .ZN(n716) );
  NOR2_X1 U772 ( .A1(n714), .A2(n694), .ZN(n715) );
  NOR2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n724) );
  AND2_X1 U774 ( .A1(n753), .A2(n739), .ZN(n719) );
  XOR2_X1 U775 ( .A(KEYINPUT82), .B(n717), .Z(n718) );
  NOR2_X1 U776 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U778 ( .A(KEYINPUT84), .B(n722), .Z(n723) );
  NAND2_X1 U779 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U780 ( .A(n726), .B(n725), .ZN(G75) );
  NAND2_X1 U781 ( .A1(n733), .A2(G469), .ZN(n731) );
  XOR2_X1 U782 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n728) );
  XNOR2_X1 U783 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U784 ( .A1(n737), .A2(n732), .ZN(G54) );
  NAND2_X1 U785 ( .A1(n733), .A2(G478), .ZN(n735) );
  XNOR2_X1 U786 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n737), .A2(n736), .ZN(G63) );
  NAND2_X1 U788 ( .A1(n739), .A2(n738), .ZN(n744) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n740) );
  XNOR2_X1 U790 ( .A(n740), .B(KEYINPUT61), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U792 ( .A1(n744), .A2(n743), .ZN(n750) );
  XNOR2_X1 U793 ( .A(n745), .B(KEYINPUT124), .ZN(n747) );
  NOR2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U795 ( .A(KEYINPUT123), .B(n748), .Z(n749) );
  XNOR2_X1 U796 ( .A(n750), .B(n749), .ZN(G69) );
  XNOR2_X1 U797 ( .A(n752), .B(n751), .ZN(n756) );
  XNOR2_X1 U798 ( .A(n753), .B(n756), .ZN(n755) );
  NAND2_X1 U799 ( .A1(n755), .A2(n754), .ZN(n761) );
  XNOR2_X1 U800 ( .A(KEYINPUT125), .B(n756), .ZN(n757) );
  XNOR2_X1 U801 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U802 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U803 ( .A1(n759), .A2(G953), .ZN(n760) );
  NAND2_X1 U804 ( .A1(n761), .A2(n760), .ZN(G72) );
  XNOR2_X1 U805 ( .A(G122), .B(KEYINPUT126), .ZN(n762) );
  XOR2_X1 U806 ( .A(n763), .B(G131), .Z(G33) );
  XOR2_X1 U807 ( .A(G137), .B(n764), .Z(G39) );
endmodule

