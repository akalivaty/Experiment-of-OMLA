//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT72), .ZN(new_n189));
  XOR2_X1   g003(.A(G116), .B(G119), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G113), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n198), .A3(new_n201), .A4(new_n196), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n202), .A2(new_n203), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n200), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n210), .A2(KEYINPUT64), .A3(G146), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT64), .B1(new_n210), .B2(G146), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G146), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n208), .B2(G143), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(KEYINPUT64), .A3(G146), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT65), .B1(new_n222), .B2(new_n215), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n210), .A2(G146), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n209), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n225), .A2(KEYINPUT66), .A3(KEYINPUT0), .A4(G128), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n209), .A2(new_n224), .A3(KEYINPUT0), .A4(G128), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n217), .A2(new_n223), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n197), .A2(G134), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n201), .B1(new_n196), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n195), .A2(new_n198), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(KEYINPUT67), .A3(new_n201), .A4(new_n196), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n234), .B2(new_n204), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n209), .A2(new_n224), .A3(new_n236), .A4(G128), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT68), .B(G128), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(G143), .B2(new_n208), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n237), .B1(new_n240), .B2(new_n222), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n207), .A2(new_n230), .B1(new_n235), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n192), .B1(new_n242), .B2(KEYINPUT30), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n245));
  OR2_X1    g059(.A1(KEYINPUT68), .A2(G128), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT68), .A2(G128), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n213), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n244), .B1(new_n249), .B2(new_n237), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n244), .B(new_n237), .C1(new_n240), .C2(new_n222), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n235), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n230), .A2(new_n207), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT30), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n241), .A2(KEYINPUT69), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n251), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n258), .A2(new_n235), .B1(new_n230), .B2(new_n207), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT30), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n243), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n192), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n265));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G210), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n265), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n189), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n235), .A2(new_n241), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n254), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n263), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n260), .B1(new_n259), .B2(KEYINPUT30), .ZN(new_n277));
  AND4_X1   g091(.A1(new_n260), .A2(new_n253), .A3(KEYINPUT30), .A4(new_n254), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n271), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n272), .A2(new_n281), .A3(KEYINPUT31), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n262), .B2(new_n271), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n253), .A2(new_n254), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(new_n192), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT28), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n274), .A2(new_n192), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n264), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n270), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n188), .B1(new_n285), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n286), .A2(new_n192), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n288), .A2(KEYINPUT29), .A3(new_n291), .A4(new_n296), .ZN(new_n297));
  OR3_X1    g111(.A1(new_n297), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n288), .A2(new_n289), .A3(new_n291), .A4(new_n270), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n262), .A2(new_n287), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n299), .B(new_n300), .C1(new_n301), .C2(new_n270), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT75), .B1(new_n297), .B2(new_n293), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n298), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n295), .A2(KEYINPUT32), .B1(new_n305), .B2(G472), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n307));
  OAI21_X1  g121(.A(KEYINPUT74), .B1(new_n295), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  INV_X1    g123(.A(new_n307), .ZN(new_n310));
  INV_X1    g124(.A(new_n294), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n282), .B2(new_n284), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n309), .B(new_n310), .C1(new_n312), .C2(new_n188), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n306), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n317), .A2(KEYINPUT76), .A3(G125), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n317), .A2(KEYINPUT76), .A3(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n317), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n328), .B2(KEYINPUT76), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT77), .A3(KEYINPUT16), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n317), .A3(G125), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n323), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n208), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n323), .A2(new_n330), .A3(G146), .A4(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  INV_X1    g150(.A(G119), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(G128), .ZN(new_n338));
  INV_X1    g152(.A(G128), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G119), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n238), .B2(G119), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n338), .B1(new_n341), .B2(new_n336), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G110), .ZN(new_n343));
  INV_X1    g157(.A(new_n341), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n335), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n345), .ZN(new_n347));
  INV_X1    g161(.A(G110), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n348), .B(new_n338), .C1(new_n341), .C2(new_n336), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n319), .A2(new_n208), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n334), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT78), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n334), .A2(new_n350), .A3(new_n354), .A4(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G137), .ZN(new_n357));
  INV_X1    g171(.A(G953), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n358), .A2(G221), .A3(G234), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n357), .B(new_n359), .Z(new_n360));
  AND3_X1   g174(.A1(new_n346), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n346), .B2(new_n356), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .A4(new_n303), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n346), .A2(new_n356), .ZN(new_n367));
  INV_X1    g181(.A(new_n360), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n346), .A2(new_n356), .A3(new_n360), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n303), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n364), .A2(new_n365), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(G234), .B2(new_n303), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n371), .A2(new_n376), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n315), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n315), .A3(new_n378), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n314), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT95), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n385), .B2(G107), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G104), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(G107), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n386), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n388), .A2(G104), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n385), .A2(G107), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n225), .B1(G128), .B2(new_n245), .ZN(new_n397));
  INV_X1    g211(.A(new_n237), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n396), .B2(new_n241), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n207), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT12), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT82), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n386), .A2(new_n389), .A3(new_n391), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G101), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(G101), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n230), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n207), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n258), .A2(KEYINPUT10), .A3(new_n396), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n409), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G140), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n358), .A2(G227), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n403), .A2(new_n418), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(KEYINPUT81), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n418), .A2(new_n422), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n409), .A2(new_n415), .A3(new_n417), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n207), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n430), .A3(G469), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n432));
  NAND2_X1  g246(.A1(G469), .A2(G902), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n424), .A2(new_n425), .B1(new_n427), .B2(new_n429), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT83), .B(G469), .C1(new_n435), .C2(G902), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n422), .B1(new_n429), .B2(new_n418), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n403), .A2(new_n422), .A3(new_n418), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n437), .B(new_n303), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n266), .A2(G143), .A3(G214), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(G143), .B1(new_n266), .B2(G214), .ZN(new_n444));
  OAI21_X1  g258(.A(G131), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n201), .A3(new_n442), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OR3_X1    g262(.A1(new_n328), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n321), .B1(KEYINPUT90), .B2(new_n319), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT19), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n334), .B(new_n448), .C1(new_n452), .C2(G146), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n443), .A2(new_n444), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT18), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n201), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n351), .B1(new_n329), .B2(new_n208), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n456), .B(new_n457), .C1(new_n455), .C2(new_n445), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G113), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(G104), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n445), .A2(new_n447), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT92), .ZN(new_n465));
  INV_X1    g279(.A(new_n445), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n333), .A3(new_n334), .A4(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n461), .B(KEYINPUT91), .Z(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n458), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(G475), .B1(new_n462), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT20), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n303), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n473), .B2(new_n303), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(KEYINPUT93), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n473), .A2(new_n478), .A3(new_n474), .A4(new_n303), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n470), .A2(new_n458), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n461), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n472), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n303), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n477), .A2(new_n479), .B1(G475), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n238), .A2(G143), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT13), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n194), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n339), .B2(G143), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n487), .B(new_n488), .Z(new_n489));
  INV_X1    g303(.A(G116), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(G122), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(G122), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(new_n388), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n488), .B(G134), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n388), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n493), .A2(new_n499), .A3(KEYINPUT14), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n493), .B2(KEYINPUT14), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n492), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n500), .B(new_n502), .C1(KEYINPUT14), .C2(new_n493), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n497), .B(new_n498), .C1(new_n388), .C2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT9), .B(G234), .Z(new_n506));
  AND3_X1   g320(.A1(new_n506), .A2(G217), .A3(new_n358), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n505), .A2(new_n507), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n303), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G478), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n510), .B(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G221), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n506), .B2(new_n303), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n441), .A2(new_n484), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  MUX2_X1   g332(.A(new_n241), .B(new_n230), .S(G125), .Z(new_n519));
  NAND2_X1  g333(.A1(new_n358), .A2(G224), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n337), .A3(G116), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT85), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n525), .B(G113), .C1(new_n522), .C2(new_n190), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n190), .A2(new_n191), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n396), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n192), .A2(new_n414), .A3(new_n412), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT86), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g346(.A(G110), .B(G122), .Z(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(KEYINPUT86), .A3(new_n529), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n530), .A2(new_n533), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n521), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n541), .A2(new_n303), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n533), .A2(KEYINPUT8), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT87), .ZN(new_n545));
  OAI22_X1  g359(.A1(new_n528), .A2(new_n545), .B1(KEYINPUT8), .B2(new_n533), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n396), .B1(new_n526), .B2(new_n527), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n528), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n544), .B1(new_n549), .B2(new_n538), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n519), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G210), .B1(G237), .B2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT88), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n542), .A2(new_n543), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n556), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n541), .A2(new_n303), .A3(new_n553), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n558), .B1(new_n559), .B2(KEYINPUT89), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n541), .A2(new_n303), .A3(new_n553), .A4(new_n554), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G952), .ZN(new_n564));
  AOI211_X1 g378(.A(G953), .B(new_n564), .C1(G234), .C2(G237), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n303), .B(new_n358), .C1(G234), .C2(G237), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT21), .B(G898), .Z(new_n569));
  OAI21_X1  g383(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G214), .B1(G237), .B2(G902), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT84), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n563), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n384), .B1(new_n518), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n563), .A2(new_n575), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n441), .A2(new_n517), .ZN(new_n579));
  INV_X1    g393(.A(new_n484), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n513), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT95), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n383), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n585));
  INV_X1    g399(.A(new_n295), .ZN(new_n586));
  OAI21_X1  g400(.A(G472), .B1(new_n312), .B2(G902), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n377), .A2(new_n315), .A3(new_n378), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n379), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n441), .A2(new_n517), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n585), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n586), .A2(new_n587), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n382), .A2(new_n592), .A3(new_n579), .A4(KEYINPUT96), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n559), .A2(new_n555), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n561), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n575), .ZN(new_n596));
  NAND2_X1  g410(.A1(G478), .A2(G902), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n505), .B(new_n507), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n511), .A3(new_n303), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(KEYINPUT33), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n597), .B(new_n599), .C1(new_n600), .C2(new_n511), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n596), .A2(new_n601), .A3(new_n484), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n591), .A2(new_n593), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT34), .B(G104), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  NAND2_X1  g419(.A1(new_n483), .A2(G475), .ZN(new_n606));
  INV_X1    g420(.A(new_n475), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n513), .B(new_n606), .C1(new_n607), .C2(new_n476), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n596), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n591), .A2(new_n593), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  NOR2_X1   g426(.A1(new_n368), .A2(KEYINPUT36), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n367), .B(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n614), .B(new_n303), .C1(new_n375), .C2(G234), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n377), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n592), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n582), .A2(new_n577), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT37), .B(G110), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT97), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n618), .B(new_n620), .ZN(G12));
  AOI21_X1  g435(.A(new_n572), .B1(new_n594), .B2(new_n561), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n590), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n566), .B1(new_n568), .B2(G900), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n608), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n624), .A2(new_n314), .A3(new_n616), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT98), .B(G128), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G30));
  XNOR2_X1  g444(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n563), .B(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n616), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n272), .A2(new_n281), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n270), .B1(new_n296), .B2(new_n264), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n303), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n308), .A2(new_n637), .A3(new_n638), .A4(new_n313), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n484), .A2(new_n514), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n633), .A2(new_n573), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n625), .B(KEYINPUT39), .Z(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n579), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT40), .Z(new_n647));
  NAND3_X1  g461(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G143), .ZN(G45));
  NOR3_X1   g463(.A1(new_n601), .A2(new_n484), .A3(new_n626), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n624), .A2(new_n314), .A3(new_n616), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G146), .ZN(G48));
  OAI21_X1  g466(.A(new_n303), .B1(new_n438), .B2(new_n439), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(KEYINPUT101), .A3(G469), .ZN(new_n654));
  NAND2_X1  g468(.A1(KEYINPUT101), .A2(G469), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n303), .B(new_n655), .C1(new_n438), .C2(new_n439), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n654), .A2(new_n517), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n314), .A2(new_n602), .A3(new_n382), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT41), .B(G113), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G15));
  NAND4_X1  g474(.A1(new_n314), .A2(new_n609), .A3(new_n382), .A4(new_n657), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G116), .ZN(G18));
  AND3_X1   g476(.A1(new_n657), .A2(new_n570), .A3(new_n622), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n314), .A2(new_n663), .A3(new_n581), .A4(new_n616), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G119), .ZN(G21));
  NAND2_X1  g479(.A1(new_n377), .A2(new_n378), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n288), .A2(new_n291), .A3(new_n296), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n293), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n285), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n187), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT102), .B(G472), .Z(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n312), .B2(G902), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n663), .A2(new_n667), .A3(new_n640), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G122), .ZN(G24));
  NAND3_X1  g490(.A1(new_n671), .A2(new_n673), .A3(new_n616), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT103), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n671), .A2(new_n673), .A3(new_n679), .A4(new_n616), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n657), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n623), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(new_n650), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G125), .ZN(G27));
  OR2_X1    g499(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n666), .B1(new_n686), .B2(new_n306), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n557), .A2(new_n573), .A3(new_n560), .A4(new_n562), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n433), .B(KEYINPUT104), .Z(new_n690));
  NAND3_X1  g504(.A1(new_n431), .A2(new_n440), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n517), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n687), .A2(new_n650), .A3(new_n689), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n688), .A2(new_n692), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n601), .A2(new_n484), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n625), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n383), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n201), .ZN(G33));
  NAND4_X1  g516(.A1(new_n383), .A2(KEYINPUT105), .A3(new_n627), .A4(new_n696), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n314), .A2(new_n382), .A3(new_n696), .A4(new_n627), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G134), .ZN(G36));
  OAI21_X1  g522(.A(G469), .B1(new_n435), .B2(KEYINPUT45), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT106), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n435), .A2(KEYINPUT45), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n690), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT107), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n712), .A2(KEYINPUT46), .A3(new_n690), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n713), .A2(new_n718), .A3(new_n714), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n717), .A3(new_n440), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n517), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT108), .B1(new_n721), .B2(new_n644), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n580), .A2(new_n601), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT43), .ZN(new_n724));
  INV_X1    g538(.A(new_n592), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n616), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n688), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n720), .A2(new_n729), .A3(new_n517), .A4(new_n645), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n726), .A2(new_n727), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n722), .A2(new_n728), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G137), .ZN(G39));
  INV_X1    g547(.A(new_n382), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n314), .A2(new_n698), .A3(new_n688), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n720), .A2(KEYINPUT47), .A3(new_n517), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT47), .B1(new_n720), .B2(new_n517), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G140), .ZN(G42));
  NAND2_X1  g553(.A1(new_n654), .A2(new_n656), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT49), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n580), .A3(new_n601), .ZN(new_n742));
  INV_X1    g556(.A(new_n639), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n666), .A2(new_n572), .A3(new_n516), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n742), .A2(new_n632), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n667), .A2(new_n724), .A3(new_n565), .A4(new_n674), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n683), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n681), .A2(new_n650), .A3(new_n696), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n698), .B1(new_n678), .B2(new_n680), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n751), .B2(new_n696), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n704), .A2(new_n705), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n704), .A2(new_n705), .ZN(new_n754));
  OAI22_X1  g568(.A1(new_n749), .A2(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n756));
  INV_X1    g570(.A(new_n697), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n514), .A2(KEYINPUT110), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n513), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n760), .A3(new_n484), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n576), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n591), .A2(new_n593), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n606), .B1(new_n607), .B2(new_n476), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n626), .B(new_n764), .C1(new_n758), .C2(new_n760), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n590), .A2(new_n688), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n314), .A3(new_n616), .A4(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n583), .A2(new_n763), .A3(new_n618), .A4(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n755), .A2(new_n756), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n751), .A2(new_n750), .A3(new_n696), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n770), .A2(new_n771), .B1(new_n703), .B2(new_n706), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n583), .A2(new_n763), .A3(new_n618), .A4(new_n767), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT115), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n701), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n658), .A2(new_n664), .A3(new_n661), .A4(new_n675), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n624), .A2(new_n314), .A3(new_n616), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n780), .A2(new_n627), .B1(new_n751), .B2(new_n683), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n573), .A2(new_n580), .A3(new_n595), .A4(new_n513), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n692), .A2(new_n616), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n639), .A3(new_n625), .A4(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(KEYINPUT52), .A3(new_n651), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n684), .A2(new_n628), .A3(new_n651), .A4(new_n784), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n779), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n786), .A2(new_n787), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n786), .A2(new_n787), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT114), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n755), .A2(new_n768), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n658), .A2(new_n675), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(KEYINPUT109), .A3(new_n661), .A4(new_n664), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n777), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n701), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n785), .A2(new_n800), .A3(new_n788), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n793), .A2(new_n794), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n779), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n790), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n794), .A2(new_n799), .A3(KEYINPUT112), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n785), .A2(new_n788), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT112), .B1(new_n794), .B2(new_n799), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n779), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n802), .A2(new_n779), .ZN(new_n814));
  OAI211_X1 g628(.A(KEYINPUT113), .B(new_n779), .C1(new_n809), .C2(new_n810), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n806), .B1(new_n816), .B2(KEYINPUT54), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n736), .A2(new_n737), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n740), .B(KEYINPUT116), .Z(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n516), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n746), .A2(new_n689), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n818), .A2(KEYINPUT118), .A3(new_n820), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n573), .B(new_n682), .C1(KEYINPUT117), .C2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n746), .A2(new_n828), .A3(new_n632), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n682), .A2(new_n688), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n382), .A2(new_n743), .A3(new_n565), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n484), .A3(new_n601), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n724), .A2(new_n565), .A3(new_n833), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n681), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n821), .A2(new_n824), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT51), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n564), .B(G953), .C1(new_n834), .C2(new_n697), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n837), .A2(new_n687), .ZN(new_n843));
  NOR2_X1   g657(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n843), .B(new_n844), .Z(new_n845));
  AND2_X1   g659(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n747), .A2(new_n817), .A3(new_n839), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(G952), .A2(G953), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n745), .B1(new_n849), .B2(new_n850), .ZN(G75));
  AND2_X1   g665(.A1(new_n790), .A2(new_n803), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n303), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT56), .B1(new_n853), .B2(G210), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n537), .A2(new_n540), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(new_n521), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT55), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n854), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n358), .A2(G952), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G51));
  NAND2_X1  g676(.A1(new_n805), .A2(KEYINPUT121), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n790), .A2(new_n803), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n790), .A2(new_n803), .A3(new_n866), .A4(new_n804), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n690), .B(KEYINPUT120), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT57), .Z(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT122), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n438), .A2(new_n439), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n874), .A3(new_n870), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n853), .A2(new_n711), .A3(new_n710), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n861), .B1(new_n876), .B2(new_n877), .ZN(G54));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n853), .A2(KEYINPUT58), .A3(G475), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n462), .A2(new_n472), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n861), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n880), .A2(new_n882), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n880), .A2(new_n879), .A3(new_n882), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G60));
  INV_X1    g702(.A(new_n600), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n597), .B(KEYINPUT59), .Z(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n817), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n868), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n891), .A2(new_n884), .A3(new_n893), .ZN(G63));
  XNOR2_X1  g708(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n375), .A2(new_n303), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n852), .A2(new_n898), .B1(new_n362), .B2(new_n361), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n864), .A2(new_n614), .A3(new_n897), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n899), .B(new_n884), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(G66));
  NAND2_X1  g720(.A1(new_n569), .A2(G224), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(G953), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n796), .A2(new_n798), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n583), .A2(new_n763), .A3(new_n618), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n908), .B1(new_n912), .B2(G953), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT126), .ZN(new_n914));
  INV_X1    g728(.A(G898), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n855), .B1(new_n915), .B2(G953), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n914), .B(new_n916), .ZN(G69));
  OAI22_X1  g731(.A1(new_n277), .A2(new_n278), .B1(KEYINPUT30), .B2(new_n242), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n452), .ZN(new_n919));
  NAND2_X1  g733(.A1(G900), .A2(G953), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n732), .A2(new_n738), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n781), .A2(new_n651), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n923), .A2(new_n776), .A3(new_n707), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n722), .A2(new_n687), .A3(new_n730), .A4(new_n782), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(KEYINPUT127), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(KEYINPUT127), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n921), .B(new_n924), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n919), .B(new_n920), .C1(new_n928), .C2(G953), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n648), .A2(new_n923), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n646), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n757), .A2(new_n761), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n383), .A2(new_n933), .A3(new_n689), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n935), .A3(new_n921), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n936), .A2(new_n358), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n929), .B1(new_n937), .B2(new_n919), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n358), .B1(G227), .B2(G900), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G72));
  NAND4_X1  g754(.A1(new_n932), .A2(new_n921), .A3(new_n912), .A4(new_n935), .ZN(new_n941));
  NAND2_X1  g755(.A1(G472), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT63), .Z(new_n943));
  AOI21_X1  g757(.A(new_n293), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n301), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n861), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n943), .B1(new_n928), .B2(new_n911), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(new_n293), .A3(new_n301), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n634), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n270), .B2(new_n301), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n816), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n949), .B1(new_n943), .B2(new_n952), .ZN(G57));
endmodule


