//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1186, new_n1187, new_n1188, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n203), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n202), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n207), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NAND2_X1  g0022(.A1(new_n204), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  OR3_X1    g0028(.A1(new_n207), .A2(KEYINPUT65), .A3(G13), .ZN(new_n229));
  OAI21_X1  g0029(.A(KEYINPUT65), .B1(new_n207), .B2(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT0), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n222), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n211), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n214), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI211_X1 g0057(.A(G226), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  OAI211_X1 g0058(.A(G232), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n254), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n252), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G238), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n267), .B1(new_n266), .B2(new_n270), .ZN(new_n273));
  OAI21_X1  g0073(.A(G169), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT14), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT14), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n276), .B(G169), .C1(new_n272), .C2(new_n273), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n272), .A2(KEYINPUT70), .A3(new_n273), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  AOI211_X1 g0080(.A(new_n280), .B(new_n267), .C1(new_n266), .C2(new_n270), .ZN(new_n281));
  OAI21_X1  g0081(.A(G179), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n266), .A2(new_n270), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(new_n280), .A3(new_n271), .ZN(new_n287));
  INV_X1    g0087(.A(new_n281), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(KEYINPUT72), .A3(G179), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n278), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n203), .A2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n226), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n292), .B1(new_n293), .B2(new_n216), .C1(new_n295), .C2(new_n214), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n225), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT11), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT11), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n292), .A2(G1), .A3(new_n302), .ZN(new_n303));
  XOR2_X1   g0103(.A(new_n303), .B(KEYINPUT12), .Z(new_n304));
  NAND3_X1  g0104(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT68), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n251), .B2(G20), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n226), .A2(KEYINPUT68), .A3(G1), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n306), .A2(new_n298), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G68), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n300), .A2(new_n301), .A3(new_n304), .A4(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n291), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n254), .B1(new_n269), .B2(G244), .ZN(new_n316));
  OR2_X1    g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(G232), .A3(new_n255), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(G1698), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n320), .B1(new_n210), .B2(new_n319), .C1(new_n321), .C2(new_n209), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT69), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n316), .B1(new_n323), .B2(new_n264), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT8), .B(G58), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n295), .B1(new_n226), .B2(new_n216), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n293), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n298), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n306), .A2(new_n216), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n310), .A2(G77), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n326), .B(new_n335), .C1(G179), .C2(new_n324), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n312), .B1(new_n289), .B2(G190), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n286), .B2(new_n271), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT71), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G190), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n287), .B2(new_n288), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT71), .ZN(new_n344));
  NOR4_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(new_n339), .A4(new_n312), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n315), .B(new_n336), .C1(new_n341), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n319), .A2(G222), .A3(new_n255), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT67), .ZN(new_n348));
  INV_X1    g0148(.A(G223), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n321), .A2(new_n349), .B1(new_n216), .B2(new_n319), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n265), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n254), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n269), .A2(G226), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n201), .B2(new_n204), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n358), .B1(new_n359), .B2(new_n295), .C1(new_n328), .C2(new_n293), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n298), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n310), .A2(G50), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(G50), .C2(new_n305), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n357), .B(new_n363), .C1(G169), .C2(new_n355), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n355), .A2(G190), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT9), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n354), .A2(G200), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n363), .A2(new_n367), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n365), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n215), .A2(G1698), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n374), .B1(G223), .B2(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n264), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n352), .B1(new_n268), .B2(new_n219), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n338), .ZN(new_n380));
  INV_X1    g0180(.A(new_n378), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n377), .A2(KEYINPUT73), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n383), .B(new_n264), .C1(new_n375), .C2(new_n376), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n380), .B1(new_n385), .B2(G190), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n256), .A2(new_n257), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n387), .B2(new_n226), .ZN(new_n388));
  AND4_X1   g0188(.A1(KEYINPUT7), .A2(new_n317), .A3(new_n226), .A4(new_n318), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n294), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n204), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n391), .A4(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n298), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n328), .A2(new_n306), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n310), .A2(new_n327), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n386), .A2(new_n399), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT17), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n385), .A2(G179), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n379), .A2(new_n325), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n404), .A2(KEYINPUT18), .A3(new_n405), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n324), .A2(G200), .ZN(new_n412));
  INV_X1    g0212(.A(new_n335), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(new_n342), .C2(new_n324), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n373), .A2(new_n403), .A3(new_n411), .A4(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n346), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n251), .A2(G45), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT76), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G41), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT76), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n251), .A4(G45), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n420), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(new_n264), .ZN(new_n427));
  OAI211_X1 g0227(.A(G257), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n319), .A2(KEYINPUT83), .A3(G257), .A4(G1698), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n319), .A2(G250), .A3(new_n255), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G294), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n430), .A2(new_n431), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n427), .A2(G264), .B1(new_n434), .B2(new_n265), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n420), .A2(new_n425), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n436), .A2(G274), .A3(new_n264), .A4(new_n421), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n325), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n265), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n426), .A2(G264), .A3(new_n264), .ZN(new_n440));
  AND4_X1   g0240(.A1(G179), .A2(new_n439), .A3(new_n440), .A4(new_n437), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT84), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n440), .A3(new_n437), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G169), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT84), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n444), .B(new_n445), .C1(new_n356), .C2(new_n443), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n226), .A2(G107), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT23), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n226), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n451), .A2(KEYINPUT22), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(KEYINPUT22), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n449), .B(new_n450), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT81), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n451), .B(KEYINPUT22), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(KEYINPUT81), .A3(new_n449), .A4(new_n450), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(KEYINPUT24), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT24), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n454), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n298), .A3(new_n461), .ZN(new_n462));
  OR2_X1    g0262(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n306), .A2(new_n210), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(KEYINPUT82), .B(KEYINPUT25), .C1(new_n305), .C2(G107), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n251), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n305), .A2(new_n467), .A3(new_n225), .A4(new_n297), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G107), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n462), .A2(new_n465), .A3(new_n466), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n447), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT85), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n447), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT21), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT78), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n321), .B2(new_n211), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n319), .A2(KEYINPUT78), .A3(G264), .A4(G1698), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n387), .A2(G303), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n319), .A2(G257), .A3(new_n255), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(new_n265), .B1(new_n427), .B2(G270), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n484), .A2(new_n437), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n468), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT79), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  INV_X1    g0290(.A(G97), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n490), .B(new_n226), .C1(G33), .C2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n298), .C1(new_n226), .C2(G116), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT20), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n251), .A2(new_n486), .A3(G13), .A4(G20), .ZN(new_n496));
  XOR2_X1   g0296(.A(new_n496), .B(KEYINPUT80), .Z(new_n497));
  NAND3_X1  g0297(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G169), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n477), .B1(new_n485), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n484), .A2(new_n437), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(KEYINPUT21), .A3(G169), .A4(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n485), .A2(G179), .A3(new_n498), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n476), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n338), .B1(new_n435), .B2(new_n437), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n443), .A2(new_n342), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n471), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G1698), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n511), .B(G244), .C1(new_n257), .C2(new_n256), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n217), .B1(new_n317), .B2(new_n318), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(KEYINPUT4), .ZN(new_n514));
  OAI21_X1  g0314(.A(G250), .B1(new_n256), .B2(new_n257), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n255), .B1(new_n515), .B2(KEYINPUT4), .ZN(new_n516));
  INV_X1    g0316(.A(new_n490), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT75), .B1(new_n518), .B2(new_n264), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n426), .A2(new_n253), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n427), .A2(G257), .B1(new_n520), .B2(new_n264), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n515), .A2(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G1698), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n510), .B1(new_n387), .B2(new_n217), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n523), .A2(new_n490), .A3(new_n512), .A4(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT75), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n526), .A3(new_n265), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n519), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G200), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n426), .A2(G257), .A3(new_n264), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n437), .B(new_n530), .C1(new_n518), .C2(new_n264), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n531), .A2(new_n342), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n305), .A2(G97), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n468), .A2(new_n491), .ZN(new_n535));
  OAI21_X1  g0335(.A(G107), .B1(new_n388), .B2(new_n389), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n210), .A2(KEYINPUT74), .ZN(new_n537));
  OR2_X1    g0337(.A1(KEYINPUT6), .A2(G97), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT74), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G107), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n537), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n537), .A2(new_n540), .B1(new_n538), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g0343(.A(G20), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n294), .A2(G77), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n536), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n535), .B1(new_n546), .B2(new_n298), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n529), .A2(new_n532), .A3(new_n534), .A4(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n226), .B(G68), .C1(new_n256), .C2(new_n257), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  INV_X1    g0350(.A(G87), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n491), .A3(new_n210), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n260), .A2(new_n226), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n550), .A2(new_n226), .A3(G33), .A4(G97), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(KEYINPUT77), .B(new_n549), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n298), .A3(new_n559), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n468), .A2(new_n330), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n330), .A2(new_n306), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n217), .A2(G1698), .ZN(new_n564));
  OAI221_X1 g0364(.A(new_n564), .B1(G238), .B2(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G116), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n264), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G250), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n419), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n251), .A2(new_n253), .A3(G45), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n264), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n325), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n317), .A2(new_n318), .B1(new_n209), .B2(new_n255), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n564), .B1(G33), .B2(G116), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n356), .B(new_n571), .C1(new_n575), .C2(new_n264), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n563), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n338), .B1(new_n567), .B2(new_n572), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n342), .B(new_n571), .C1(new_n575), .C2(new_n264), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n469), .A2(G87), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(new_n562), .A3(new_n560), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n519), .A2(new_n521), .A3(new_n527), .A4(new_n356), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n547), .A2(new_n534), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n531), .A2(new_n325), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n548), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n509), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n485), .A2(new_n338), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n501), .A2(new_n342), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n592), .A2(new_n498), .A3(new_n593), .ZN(new_n594));
  NOR4_X1   g0394(.A1(new_n417), .A2(new_n506), .A3(new_n591), .A4(new_n594), .ZN(G372));
  NOR2_X1   g0395(.A1(new_n341), .A2(new_n345), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n336), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n403), .B1(new_n597), .B2(new_n314), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n411), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n371), .A2(new_n372), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n365), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n444), .B1(new_n356), .B2(new_n443), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n504), .B1(new_n471), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n591), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT87), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n534), .A2(new_n547), .B1(new_n531), .B2(new_n325), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(new_n578), .A3(new_n583), .A4(new_n586), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT26), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n589), .B2(new_n584), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT86), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n612), .B(new_n608), .C1(new_n589), .C2(new_n584), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n578), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n605), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n607), .A2(new_n608), .ZN(new_n617));
  INV_X1    g0417(.A(new_n613), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n607), .B2(new_n608), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(KEYINPUT87), .A3(new_n578), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n604), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n601), .B1(new_n417), .B2(new_n622), .ZN(G369));
  NAND3_X1  g0423(.A1(new_n251), .A2(new_n226), .A3(G13), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G213), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g0427(.A(new_n627), .B(KEYINPUT88), .Z(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G343), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n504), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n471), .A2(new_n631), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(new_n509), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n476), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n472), .A2(new_n632), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT90), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n642), .B(new_n639), .C1(new_n476), .C2(new_n637), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n634), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n471), .A2(new_n602), .A3(new_n632), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n641), .A2(new_n643), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n631), .A2(new_n498), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n504), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n594), .A2(new_n504), .A3(new_n648), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n651), .B2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n646), .A2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n231), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G41), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n552), .A2(G116), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n658), .A2(new_n251), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n224), .B2(new_n658), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT28), .Z(new_n662));
  NOR3_X1   g0462(.A1(new_n509), .A2(new_n590), .A3(new_n594), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(new_n476), .A3(new_n505), .A4(new_n632), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n571), .B1(new_n575), .B2(new_n264), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n531), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(new_n441), .A3(new_n484), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT30), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n666), .A2(KEYINPUT30), .A3(new_n441), .A4(new_n484), .ZN(new_n670));
  AOI21_X1  g0470(.A(G179), .B1(new_n484), .B2(new_n437), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n443), .A3(new_n665), .A4(new_n528), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n631), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT31), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n548), .A2(new_n589), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n471), .A2(new_n507), .A3(new_n508), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n506), .A2(new_n583), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n615), .B1(new_n617), .B2(new_n610), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT29), .A3(new_n632), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n616), .A2(new_n621), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n591), .A2(new_n603), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n631), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n677), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n662), .B1(new_n690), .B2(G1), .ZN(G364));
  OR2_X1    g0491(.A1(new_n653), .A2(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n302), .A2(G20), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n251), .B1(new_n693), .B2(G45), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n658), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n692), .A2(new_n654), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(G13), .A2(G33), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G20), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n652), .B(new_n701), .C1(new_n651), .C2(new_n649), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n225), .B1(G20), .B2(new_n325), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n246), .A2(G45), .ZN(new_n707));
  INV_X1    g0507(.A(G45), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n223), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n319), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G355), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n231), .B1(new_n711), .B2(new_n387), .ZN(new_n712));
  OAI221_X1 g0512(.A(new_n706), .B1(new_n486), .B2(new_n231), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G179), .A2(G200), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(G20), .A3(new_n342), .ZN(new_n715));
  INV_X1    g0515(.A(G159), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT32), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n226), .A2(G179), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(G190), .A3(G200), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n551), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n226), .B1(new_n714), .B2(G190), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n491), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n721), .A2(new_n723), .A3(new_n387), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n342), .A3(G200), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n718), .B(new_n724), .C1(new_n210), .C2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n226), .A2(new_n356), .A3(G190), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n338), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT92), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(G20), .A2(G179), .A3(G190), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n338), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n734), .A2(G77), .B1(G50), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n735), .A2(G200), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n202), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n727), .A2(G200), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n726), .B(new_n741), .C1(G68), .C2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G317), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT33), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(KEYINPUT33), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G294), .ZN(new_n749));
  INV_X1    g0549(.A(G303), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n748), .B1(new_n749), .B2(new_n722), .C1(new_n750), .C2(new_n720), .ZN(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n733), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n736), .A2(G326), .ZN(new_n754));
  INV_X1    g0554(.A(new_n725), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n319), .B1(new_n755), .B2(G283), .ZN(new_n756));
  INV_X1    g0556(.A(new_n715), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G329), .ZN(new_n758));
  INV_X1    g0558(.A(G322), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n756), .B(new_n758), .C1(new_n739), .C2(new_n759), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n751), .A2(new_n753), .A3(new_n754), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n703), .B1(new_n744), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n702), .A2(new_n713), .A3(new_n696), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n698), .A2(new_n763), .ZN(G396));
  OAI21_X1  g0564(.A(new_n414), .B1(new_n413), .B2(new_n632), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n336), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n336), .A2(new_n631), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT95), .B1(new_n687), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT95), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n622), .A2(new_n771), .A3(new_n631), .A4(new_n768), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n770), .A2(new_n772), .B1(new_n687), .B2(new_n769), .ZN(new_n773));
  INV_X1    g0573(.A(new_n677), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n697), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n768), .A2(new_n699), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n703), .A2(new_n699), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n216), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n387), .B1(new_n752), .B2(new_n715), .C1(new_n733), .C2(new_n486), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n720), .A2(new_n210), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n755), .A2(G87), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT94), .B(G283), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n742), .B2(new_n784), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n780), .A2(new_n723), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n736), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n786), .B1(new_n749), .B2(new_n739), .C1(new_n750), .C2(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n743), .A2(G150), .B1(G143), .B2(new_n738), .ZN(new_n789));
  INV_X1    g0589(.A(G137), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n789), .B1(new_n790), .B2(new_n787), .C1(new_n733), .C2(new_n716), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT34), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n792), .B1(new_n214), .B2(new_n720), .C1(new_n203), .C2(new_n725), .ZN(new_n793));
  INV_X1    g0593(.A(G132), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n319), .B1(new_n715), .B2(new_n794), .C1(new_n202), .C2(new_n722), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n788), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n703), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n777), .A2(new_n696), .A3(new_n779), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n776), .A2(new_n798), .ZN(G384));
  OAI211_X1 g0599(.A(new_n683), .B(new_n416), .C1(KEYINPUT29), .C2(new_n687), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n601), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT102), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT38), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n404), .A2(new_n628), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n804), .A2(new_n402), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT37), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n805), .A2(KEYINPUT101), .A3(new_n806), .A4(new_n407), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n407), .A2(new_n804), .A3(new_n806), .A4(new_n402), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT101), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n407), .A2(new_n402), .A3(new_n804), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(KEYINPUT37), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n807), .A2(KEYINPUT100), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n804), .B1(new_n411), .B2(new_n403), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n807), .A2(new_n810), .B1(new_n812), .B2(KEYINPUT100), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n803), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n812), .A2(new_n808), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n815), .A2(KEYINPUT38), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n632), .A2(new_n313), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n314), .B2(new_n596), .ZN(new_n823));
  INV_X1    g0623(.A(new_n822), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n341), .B2(new_n345), .C1(new_n291), .C2(new_n313), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n676), .A2(new_n826), .A3(new_n769), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n821), .A2(new_n827), .A3(KEYINPUT40), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT40), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n676), .A2(new_n826), .A3(new_n769), .ZN(new_n830));
  INV_X1    g0630(.A(new_n819), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n803), .B1(new_n831), .B2(new_n814), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n820), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n829), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n828), .A2(G330), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n774), .A2(new_n416), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n828), .A2(new_n676), .A3(new_n834), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n417), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n802), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n767), .B(KEYINPUT97), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n770), .B2(new_n772), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n820), .A2(new_n832), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n826), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n411), .A2(new_n628), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT39), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n821), .B2(new_n847), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n314), .A2(new_n632), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n846), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n840), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n251), .B2(new_n693), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n542), .A2(new_n543), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n486), .B1(new_n856), .B2(KEYINPUT35), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n857), .B(new_n227), .C1(KEYINPUT35), .C2(new_n856), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT36), .ZN(new_n859));
  OR3_X1    g0659(.A1(new_n201), .A2(KEYINPUT96), .A3(new_n203), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n224), .A2(G77), .A3(new_n392), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT96), .B1(new_n201), .B2(new_n203), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(G1), .A3(new_n302), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n855), .A2(new_n859), .A3(new_n864), .ZN(G367));
  NAND2_X1  g0665(.A1(new_n734), .A2(new_n201), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n725), .A2(new_n216), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n720), .A2(new_n202), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n867), .B(new_n868), .C1(G150), .C2(new_n738), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n722), .A2(new_n203), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n736), .A2(G143), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n790), .B2(new_n715), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n870), .B(new_n872), .C1(G159), .C2(new_n743), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n866), .A2(new_n319), .A3(new_n869), .A4(new_n873), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n387), .B1(new_n715), .B2(new_n745), .C1(new_n739), .C2(new_n750), .ZN(new_n875));
  INV_X1    g0675(.A(new_n722), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(G107), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n720), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(G116), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT46), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n755), .A2(G97), .B1(G311), .B2(new_n736), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n743), .A2(G294), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n877), .A2(new_n880), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n733), .A2(new_n784), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n874), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT47), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n703), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n657), .A2(new_n319), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n706), .B1(new_n231), .B2(new_n330), .C1(new_n242), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n696), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT110), .ZN(new_n892));
  INV_X1    g0692(.A(new_n701), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n560), .A2(new_n562), .A3(new_n582), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n631), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n585), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n615), .A2(new_n894), .A3(new_n631), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n887), .B(new_n892), .C1(new_n893), .C2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT106), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT42), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n447), .A2(new_n471), .A3(new_n474), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n474), .B1(new_n447), .B2(new_n471), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n679), .A2(new_n635), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n640), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n642), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n638), .A2(KEYINPUT90), .A3(new_n640), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n633), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n631), .A2(new_n587), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n548), .A2(new_n589), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT104), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n606), .A2(new_n631), .A3(new_n586), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n901), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n589), .B1(new_n912), .B2(new_n476), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT105), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT105), .B(new_n589), .C1(new_n912), .C2(new_n476), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n632), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n900), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n909), .A2(new_n901), .A3(new_n914), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n634), .B(new_n914), .C1(new_n641), .C2(new_n643), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(KEYINPUT106), .A3(new_n920), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n898), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(KEYINPUT43), .B2(new_n898), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n922), .A2(new_n929), .A3(new_n923), .A4(new_n926), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT107), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n655), .A2(new_n914), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT108), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n931), .B(new_n938), .C1(new_n934), .C2(new_n935), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n644), .A2(new_n645), .A3(new_n914), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT45), .ZN(new_n944));
  INV_X1    g0744(.A(new_n914), .ZN(new_n945));
  INV_X1    g0745(.A(new_n645), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n909), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT44), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT44), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n646), .A2(new_n949), .A3(new_n945), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n655), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n948), .A2(new_n950), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT45), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n943), .B(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n655), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT109), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n654), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n647), .A2(new_n633), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n644), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n644), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n653), .A2(G330), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n689), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n952), .A2(new_n957), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n690), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n658), .B(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n695), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n899), .B1(new_n942), .B2(new_n969), .ZN(G387));
  OAI22_X1  g0770(.A1(new_n733), .A2(new_n203), .B1(new_n330), .B2(new_n722), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n725), .A2(new_n491), .B1(new_n359), .B2(new_n715), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n720), .A2(new_n216), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n972), .A2(new_n973), .A3(new_n387), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT111), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n971), .B(new_n975), .C1(G50), .C2(new_n738), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n716), .B2(new_n787), .C1(new_n328), .C2(new_n742), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n743), .A2(G311), .B1(G317), .B2(new_n738), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n759), .B2(new_n787), .C1(new_n733), .C2(new_n750), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT48), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n749), .B2(new_n720), .C1(new_n722), .C2(new_n784), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT49), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n755), .A2(G116), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n757), .A2(G326), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n983), .A2(new_n387), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n982), .A2(KEYINPUT49), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n977), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n703), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n239), .A2(new_n708), .A3(new_n319), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n328), .A2(KEYINPUT50), .A3(G50), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT50), .B1(new_n328), .B2(G50), .ZN(new_n992));
  NAND2_X1  g0792(.A1(G68), .A2(G77), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n708), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n659), .B1(new_n994), .B2(new_n387), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n231), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n996), .B(new_n706), .C1(new_n210), .C2(new_n231), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n696), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n647), .B2(new_n701), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n961), .A2(new_n964), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n695), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n658), .B1(new_n1000), .B2(new_n690), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n965), .ZN(G393));
  NAND2_X1  g0803(.A1(new_n952), .A2(new_n957), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n965), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(new_n658), .A3(new_n966), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n952), .A2(new_n957), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n945), .A2(new_n701), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n231), .A2(new_n491), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1010), .B(new_n705), .C1(new_n249), .C2(new_n888), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n738), .A2(G159), .B1(new_n736), .B2(G150), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n757), .A2(G143), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1014), .A2(new_n319), .A3(new_n782), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n733), .A2(new_n328), .B1(new_n216), .B2(new_n722), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(G68), .C2(new_n878), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n201), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n742), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT113), .Z(new_n1021));
  NOR2_X1   g0821(.A1(new_n742), .A2(new_n750), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n387), .B1(new_n759), .B2(new_n715), .C1(new_n733), .C2(new_n749), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G107), .B2(new_n755), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n738), .A2(G311), .B1(new_n736), .B2(G317), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT52), .Z(new_n1026));
  AOI22_X1  g0826(.A1(new_n878), .A2(new_n783), .B1(new_n876), .B2(G116), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1021), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n697), .B(new_n1011), .C1(new_n1029), .C2(new_n703), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1008), .A2(new_n695), .B1(new_n1009), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1007), .A2(new_n1031), .ZN(G390));
  NAND4_X1  g0832(.A1(new_n676), .A2(new_n826), .A3(G330), .A4(new_n769), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT114), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n851), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n631), .B1(new_n680), .B2(new_n681), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n841), .B1(new_n1038), .B2(new_n769), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n826), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n821), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n851), .B1(new_n843), .B2(new_n826), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1036), .B(new_n1041), .C1(new_n1042), .C2(new_n849), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1041), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT98), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n841), .B(new_n1045), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n614), .A2(new_n605), .A3(new_n615), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT87), .B1(new_n620), .B2(new_n578), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n686), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n632), .A3(new_n769), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n771), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n687), .A2(KEYINPUT95), .A3(new_n769), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1046), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1037), .B1(new_n1053), .B2(new_n1040), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n849), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1044), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1033), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1043), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n800), .A2(new_n601), .A3(new_n836), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n676), .A2(G330), .A3(new_n769), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n1040), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n1033), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n843), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1034), .A2(new_n1035), .A3(new_n1061), .A4(new_n1039), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1059), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1041), .B1(new_n1042), .B2(new_n849), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n1033), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1065), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n1043), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1066), .A2(new_n658), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1055), .A2(new_n699), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n778), .A2(new_n328), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n734), .A2(G97), .B1(G107), .B2(new_n743), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT117), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT117), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n725), .A2(new_n203), .B1(new_n749), .B2(new_n715), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n387), .B1(new_n739), .B2(new_n486), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G283), .C2(new_n736), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n721), .B(new_n1080), .C1(G77), .C2(new_n876), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n722), .A2(new_n716), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n387), .B1(new_n755), .B2(new_n201), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT54), .B(G143), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n734), .B2(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n742), .A2(new_n790), .B1(new_n739), .B2(new_n794), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1083), .B2(KEYINPUT115), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n720), .A2(new_n359), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1090));
  XNOR2_X1  g0890(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n736), .A2(G128), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1086), .A2(new_n1088), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1082), .B(new_n1093), .C1(G125), .C2(new_n757), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n703), .B1(new_n1081), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1072), .A2(new_n696), .A3(new_n1073), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1058), .B2(new_n695), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1071), .A2(new_n1098), .ZN(G378));
  AOI21_X1  g0899(.A(new_n1059), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n658), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(KEYINPUT57), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n694), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT121), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT120), .B1(new_n853), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT119), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n600), .A2(new_n364), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT118), .Z(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1110), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n373), .A2(new_n1112), .ZN(new_n1113));
  AND4_X1   g0913(.A1(new_n363), .A2(new_n1111), .A3(new_n628), .A4(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1111), .A2(new_n1113), .B1(new_n363), .B2(new_n628), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n835), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n828), .A2(new_n1116), .A3(G330), .A4(new_n834), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(KEYINPUT120), .A3(new_n1119), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1106), .A2(new_n1120), .B1(new_n1122), .B2(new_n853), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1104), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n700), .ZN(new_n1126));
  INV_X1    g0926(.A(G124), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n262), .B1(new_n715), .B2(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n742), .A2(new_n794), .B1(new_n722), .B2(new_n359), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1085), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n733), .A2(new_n790), .B1(new_n720), .B2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1129), .B(new_n1131), .C1(G125), .C2(new_n736), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n739), .ZN(new_n1134));
  AOI211_X1 g0934(.A(G41), .B(new_n1128), .C1(new_n1134), .C2(KEYINPUT59), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(KEYINPUT59), .B2(new_n1134), .C1(new_n716), .C2(new_n725), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n733), .A2(new_n330), .B1(new_n203), .B2(new_n722), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n319), .B(new_n1137), .C1(G283), .C2(new_n757), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n263), .B1(new_n725), .B2(new_n202), .C1(new_n742), .C2(new_n491), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n973), .B(new_n1139), .C1(G107), .C2(new_n738), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(new_n486), .C2(new_n787), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT58), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n214), .B1(new_n256), .B2(G41), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n703), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n778), .A2(new_n1019), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1126), .A2(new_n697), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1120), .B(new_n853), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1069), .B1(new_n1068), .B2(new_n1043), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n1059), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n658), .A2(KEYINPUT57), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1124), .A2(new_n1154), .ZN(G375));
  OAI221_X1 g0955(.A(new_n387), .B1(new_n715), .B2(new_n750), .C1(new_n720), .C2(new_n491), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n734), .B2(G107), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n743), .A2(G116), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n738), .A2(G283), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n787), .A2(new_n749), .B1(new_n330), .B2(new_n722), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(new_n867), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n734), .A2(G150), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n736), .A2(G132), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n319), .B1(new_n1133), .B2(new_n715), .C1(new_n1130), .C2(new_n742), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G137), .B2(new_n738), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n755), .A2(G58), .B1(new_n876), .B2(G50), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n720), .A2(new_n716), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n703), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n696), .B(new_n1171), .C1(new_n826), .C2(new_n700), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n203), .B2(new_n778), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n695), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT122), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1063), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1069), .A2(new_n968), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(G381));
  NOR2_X1   g0980(.A1(G375), .A2(G378), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(G381), .A2(G384), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G393), .A2(G396), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(G387), .A2(G390), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(G407));
  NAND2_X1  g0985(.A1(new_n630), .A2(G213), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT123), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1181), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(G407), .A2(G213), .A3(new_n1188), .ZN(G409));
  INV_X1    g0989(.A(KEYINPUT62), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1058), .A2(new_n695), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1096), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1151), .A2(new_n1101), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1070), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1124), .B2(new_n1154), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1123), .B(new_n968), .C1(new_n1151), .C2(new_n1059), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1149), .B1(new_n1150), .B2(new_n695), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1196), .A2(new_n1098), .A3(new_n1071), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1187), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT60), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1178), .B1(new_n1065), .B2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1063), .A2(new_n1059), .A3(new_n1064), .A4(KEYINPUT60), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n1203), .A3(new_n658), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT124), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1202), .A2(new_n1203), .A3(KEYINPUT124), .A4(new_n658), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1177), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(G384), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1206), .A2(new_n1177), .A3(G384), .A4(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1195), .A2(new_n1200), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1190), .B1(new_n1213), .B2(KEYINPUT127), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT61), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT125), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1210), .A2(new_n1216), .A3(new_n1211), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1187), .A2(G2897), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1217), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1150), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1153), .B1(new_n1100), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1149), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1123), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1102), .B1(new_n1151), .B2(new_n1059), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n694), .ZN(new_n1229));
  OAI21_X1  g1029(.A(G378), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1222), .A2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1210), .A2(new_n1216), .A3(new_n1211), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1219), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1221), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1222), .A2(new_n1230), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT127), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1237), .A3(KEYINPUT62), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1214), .A2(new_n1215), .A3(new_n1234), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT126), .ZN(new_n1240));
  INV_X1    g1040(.A(G390), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(G387), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(G393), .B(G396), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G390), .B(new_n899), .C1(new_n942), .C2(new_n969), .ZN(new_n1244));
  AND4_X1   g1044(.A1(new_n1240), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(KEYINPUT126), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1246), .A2(new_n1243), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1239), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1213), .A2(KEYINPUT63), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1248), .A2(KEYINPUT61), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1230), .A2(new_n1222), .B1(new_n1232), .B2(new_n1219), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1253), .B2(new_n1221), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1250), .B(new_n1251), .C1(new_n1254), .C2(new_n1213), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1249), .A2(new_n1255), .ZN(G405));
  OR2_X1    g1056(.A1(new_n1181), .A2(new_n1195), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1248), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1181), .A2(new_n1195), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1212), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1258), .A2(new_n1260), .A3(new_n1235), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(G402));
endmodule


