//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n626, new_n628, new_n629, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n453), .A2(G567), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT68), .B(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(new_n464), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND3_X1  g055(.A1(new_n474), .A2(G2105), .A3(new_n464), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(G136), .B2(new_n477), .ZN(G162));
  AND2_X1   g063(.A1(new_n464), .A2(new_n465), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n475), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n477), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n482), .A2(G126), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n494), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G651), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G88), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n504), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT70), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n514));
  OAI211_X1 g089(.A(G543), .B(new_n507), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n500), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n512), .A2(new_n517), .A3(new_n500), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n509), .A2(G62), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(KEYINPUT72), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n509), .A2(new_n523), .A3(G62), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n504), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n518), .A2(new_n520), .B1(new_n527), .B2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NOR2_X1   g105(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n503), .B2(new_n505), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(G89), .A3(new_n509), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n537), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n509), .A2(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n515), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n532), .A2(KEYINPUT74), .A3(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n540), .B1(new_n544), .B2(G51), .ZN(G168));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OR2_X1    g121(.A1(KEYINPUT5), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(KEYINPUT5), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(G77), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n506), .A2(G90), .A3(new_n507), .A4(new_n509), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n544), .B2(G52), .ZN(G171));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n542), .B2(new_n543), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n532), .A2(G81), .A3(new_n509), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n547), .B2(new_n548), .ZN(new_n559));
  AND2_X1   g134(.A1(G68), .A2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n532), .A2(new_n509), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(G91), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n516), .A2(G53), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI211_X1 g150(.A(KEYINPUT75), .B(KEYINPUT9), .C1(new_n515), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n504), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n572), .A2(new_n577), .A3(new_n579), .ZN(G299));
  AND4_X1   g155(.A1(KEYINPUT74), .A2(new_n506), .A3(G543), .A4(new_n507), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT74), .B1(new_n532), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(G52), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n553), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G301));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  INV_X1    g161(.A(G51), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n542), .B2(new_n543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n588), .B2(new_n540), .ZN(new_n589));
  OAI21_X1  g164(.A(G51), .B1(new_n581), .B2(new_n582), .ZN(new_n590));
  INV_X1    g165(.A(new_n540), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT77), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(G286));
  NAND3_X1  g168(.A1(new_n570), .A2(G87), .A3(new_n571), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n509), .A2(G74), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n516), .A2(G49), .B1(new_n595), .B2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G288));
  AOI22_X1  g172(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n504), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n532), .A2(G48), .A3(G543), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n570), .A2(G86), .A3(new_n571), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G305));
  AND2_X1   g179(.A1(new_n544), .A2(G47), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n504), .ZN(new_n607));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n569), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n605), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n570), .A2(G92), .A3(new_n571), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n613), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n570), .A2(G92), .A3(new_n571), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n510), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n544), .A2(G54), .B1(G651), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n614), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n611), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n611), .B1(new_n621), .B2(G868), .ZN(G321));
  MUX2_X1   g198(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g199(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n621), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n621), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g206(.A(G323), .B(new_n631), .ZN(G282));
  NOR2_X1   g207(.A1(new_n490), .A2(new_n470), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n477), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n482), .A2(G123), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n639), .A2(new_n475), .A3(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n475), .B2(G111), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n637), .B(new_n638), .C1(new_n640), .C2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n636), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT83), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G14), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(G401));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT84), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(new_n684), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT20), .Z(new_n688));
  AOI211_X1 g263(.A(new_n686), .B(new_n688), .C1(new_n681), .C2(new_n685), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G29), .A2(G35), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G162), .B2(G29), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT29), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G2090), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n701), .A2(G33), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT25), .Z(new_n704));
  INV_X1    g279(.A(G139), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI221_X1 g281(.A(new_n704), .B1(new_n476), .B2(new_n705), .C1(new_n706), .C2(new_n475), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n702), .B1(new_n707), .B2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G2072), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT91), .Z(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NOR2_X1   g287(.A1(G168), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n712), .B2(G21), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT92), .B(G1966), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G16), .A2(G19), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n563), .B2(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G1341), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n714), .B2(new_n715), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n700), .A2(new_n711), .A3(new_n716), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n701), .A2(G32), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n477), .A2(G141), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n482), .A2(G129), .ZN(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT26), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n471), .A2(G105), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n723), .A2(new_n724), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n722), .B1(new_n731), .B2(new_n701), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT27), .ZN(new_n733));
  INV_X1    g308(.A(G1996), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n621), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G4), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT89), .B(G1348), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n712), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G1956), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n737), .A2(new_n738), .ZN(new_n746));
  NOR4_X1   g321(.A1(new_n735), .A2(new_n739), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n748), .B2(KEYINPUT24), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(KEYINPUT24), .B2(new_n748), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n479), .B2(new_n701), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G11), .ZN(new_n755));
  INV_X1    g330(.A(G28), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n758), .A2(KEYINPUT94), .B1(KEYINPUT30), .B2(new_n756), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n755), .B1(new_n759), .B2(new_n760), .C1(new_n708), .C2(new_n709), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n753), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n701), .B2(new_n645), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n701), .A2(G27), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT95), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n701), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(G2078), .ZN(new_n767));
  NOR2_X1   g342(.A1(G171), .A2(new_n712), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G5), .B2(new_n712), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n766), .A2(G2078), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n767), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n701), .A2(G26), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n477), .A2(G140), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n482), .A2(G128), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n475), .A2(G116), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n777), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2067), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G1341), .B2(new_n718), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n763), .A2(new_n774), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n721), .A2(new_n747), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT97), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT88), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n712), .A2(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n712), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT87), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n712), .A2(G6), .ZN(new_n798));
  INV_X1    g373(.A(G305), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n712), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT32), .B(G1981), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n712), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(G288), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n712), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n796), .A2(new_n797), .A3(new_n802), .A4(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n701), .A2(G25), .ZN(new_n810));
  OAI21_X1  g385(.A(KEYINPUT85), .B1(G95), .B2(G2105), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR3_X1   g387(.A1(KEYINPUT85), .A2(G95), .A3(G2105), .ZN(new_n813));
  OAI221_X1 g388(.A(G2104), .B1(G107), .B2(new_n475), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G131), .ZN(new_n815));
  INV_X1    g390(.A(G119), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n814), .B1(new_n476), .B2(new_n815), .C1(new_n816), .C2(new_n481), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT86), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n810), .B1(new_n818), .B2(new_n701), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n712), .A2(G24), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n605), .A2(new_n609), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(new_n712), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1986), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n822), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n808), .B2(KEYINPUT34), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n789), .B(new_n790), .C1(new_n809), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n788), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n809), .A2(new_n829), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n790), .B1(new_n832), .B2(new_n789), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n809), .A2(new_n829), .A3(new_n789), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(G311));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n789), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n836), .A2(KEYINPUT36), .A3(new_n834), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n837), .A2(new_n830), .A3(new_n788), .ZN(G150));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n616), .A3(new_n620), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n626), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT99), .B1(new_n556), .B2(new_n562), .ZN(new_n841));
  OAI21_X1  g416(.A(G43), .B1(new_n581), .B2(new_n582), .ZN(new_n842));
  INV_X1    g417(.A(new_n562), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(G55), .B1(new_n581), .B2(new_n582), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n847));
  AND2_X1   g422(.A1(G80), .A2(G543), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n509), .B2(G67), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n849), .B2(new_n504), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n547), .B2(new_n548), .ZN(new_n852));
  OAI211_X1 g427(.A(KEYINPUT98), .B(G651), .C1(new_n852), .C2(new_n848), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n511), .A2(G93), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n846), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n841), .A2(new_n845), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n850), .A2(new_n853), .B1(new_n511), .B2(G93), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n563), .A2(new_n844), .A3(new_n846), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n840), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  AOI21_X1  g439(.A(G860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n856), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  XOR2_X1   g445(.A(new_n817), .B(KEYINPUT103), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n634), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n730), .B(new_n707), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G164), .B(new_n782), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n482), .A2(G130), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n877), .A2(new_n475), .A3(G118), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n475), .B2(G118), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n876), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(G142), .B2(new_n477), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n875), .B(new_n882), .Z(new_n883));
  OR2_X1    g458(.A1(new_n874), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n874), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n645), .B(G160), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G162), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT106), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(KEYINPUT105), .B(G37), .Z(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n888), .A3(new_n885), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n892), .A2(KEYINPUT104), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(KEYINPUT104), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n890), .B(new_n891), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g471(.A(new_n628), .B(KEYINPUT107), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n860), .ZN(new_n898));
  INV_X1    g473(.A(G299), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n621), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n839), .A2(G299), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT41), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n900), .A2(KEYINPUT41), .A3(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n860), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n897), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n839), .B(new_n899), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(new_n804), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n825), .A2(G288), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n525), .B(new_n526), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n512), .A2(new_n517), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT71), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n519), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n918), .A3(G305), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G305), .B1(new_n915), .B2(new_n918), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(G303), .A2(new_n799), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(new_n912), .A3(new_n919), .A4(new_n913), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n911), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n911), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n856), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(G868), .B2(new_n930), .ZN(G295));
  OAI21_X1  g506(.A(new_n929), .B1(G868), .B2(new_n930), .ZN(G331));
  INV_X1    g507(.A(KEYINPUT112), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n590), .A2(new_n591), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT108), .B1(new_n935), .B2(G171), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n937));
  NAND3_X1  g512(.A1(G301), .A2(G168), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n589), .A2(new_n592), .A3(G171), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n905), .ZN(new_n942));
  AOI22_X1  g517(.A1(G286), .A2(G171), .B1(new_n936), .B2(new_n938), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n860), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n907), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT110), .B1(new_n943), .B2(new_n860), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n905), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n943), .B2(new_n860), .ZN(new_n950));
  AND4_X1   g525(.A1(new_n949), .A2(new_n860), .A3(new_n940), .A4(new_n939), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n946), .B(new_n948), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n903), .A2(new_n902), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n925), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n934), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI211_X1 g531(.A(new_n945), .B(new_n925), .C1(new_n953), .C2(new_n952), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT43), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n960), .B(KEYINPUT43), .C1(new_n956), .C2(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n942), .A2(new_n944), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n953), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n908), .B2(new_n952), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n925), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n954), .A2(new_n955), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n891), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n961), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT43), .A4(new_n891), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n967), .B1(new_n956), .B2(new_n957), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n933), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g551(.A(KEYINPUT112), .B(new_n974), .C1(new_n969), .C2(new_n970), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n494), .B2(new_n498), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT113), .B(G40), .Z(new_n984));
  NAND4_X1  g559(.A1(new_n473), .A2(new_n478), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n478), .A2(new_n469), .A3(new_n472), .A4(new_n984), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT114), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n982), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  AND2_X1   g564(.A1(G290), .A2(G1986), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n734), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(new_n730), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT115), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n782), .B(G2067), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n731), .A2(new_n734), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n988), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n817), .B(new_n821), .Z(new_n998));
  NAND2_X1  g573(.A1(new_n988), .A2(new_n998), .ZN(new_n999));
  AND4_X1   g574(.A1(new_n991), .A2(new_n994), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n498), .ZN(new_n1001));
  INV_X1    g576(.A(new_n492), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT4), .B1(new_n476), .B2(new_n491), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n987), .A2(new_n985), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n982), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G2078), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1008), .B2(G2078), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1007), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1014), .B(new_n979), .C1(new_n494), .C2(new_n498), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n770), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1012), .A2(new_n1013), .A3(G301), .A4(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT125), .Z(new_n1020));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1006), .A2(new_n982), .ZN(new_n1022));
  NAND3_X1  g597(.A1(G160), .A2(G40), .A3(new_n1011), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1013), .B(new_n1018), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1021), .B1(new_n1024), .B2(G171), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n1007), .B2(new_n1005), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n804), .A2(G1976), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1028), .A2(KEYINPUT117), .A3(KEYINPUT52), .A4(new_n1029), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  NAND3_X1  g610(.A1(G288), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G305), .A2(G1981), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT118), .B(G86), .Z(new_n1041));
  OAI21_X1  g616(.A(new_n601), .B1(new_n569), .B2(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1042), .A2(KEYINPUT119), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n599), .B1(new_n1042), .B2(KEYINPUT119), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1038), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1028), .A3(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1037), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT116), .B(G1971), .Z(new_n1051));
  NAND2_X1  g626(.A1(new_n1008), .A2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n980), .A2(KEYINPUT50), .B1(new_n987), .B2(new_n985), .ZN(new_n1053));
  INV_X1    g628(.A(G2090), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1016), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(G8), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1050), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1016), .B1(new_n1015), .B2(KEYINPUT121), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1053), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1062), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1017), .B1(new_n1053), .B2(new_n1064), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1015), .A2(KEYINPUT121), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(KEYINPUT122), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1054), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1027), .B1(new_n1070), .B2(new_n1052), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1059), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1061), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1012), .A2(new_n1013), .A3(new_n1018), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G171), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(G171), .B2(new_n1024), .ZN(new_n1077));
  INV_X1    g652(.A(G1966), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1008), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1053), .A2(new_n752), .A3(new_n1016), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(G168), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  AOI21_X1  g657(.A(G168), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT51), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1085), .A3(G8), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1077), .A2(new_n1021), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1026), .A2(new_n1074), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  XOR2_X1   g664(.A(G299), .B(KEYINPUT57), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n744), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT123), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1094), .A3(new_n744), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1009), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1090), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1090), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1098), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1100), .B(new_n1101), .C1(new_n1093), .C2(new_n1095), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1089), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1096), .A2(new_n1090), .A3(new_n1098), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1090), .B(KEYINPUT124), .Z(new_n1106));
  OAI211_X1 g681(.A(new_n1104), .B(KEYINPUT61), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1008), .A2(G1996), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT58), .B(G1341), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1007), .B2(new_n1005), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n563), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g688(.A(G2067), .B(new_n980), .C1(new_n985), .C2(new_n987), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n738), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n621), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1113), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n621), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n1116), .A3(new_n839), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1103), .A2(new_n1107), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1121), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1104), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1088), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1060), .A2(new_n1037), .A3(new_n1049), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1027), .B(G286), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1056), .A2(G8), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1073), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1130), .A2(KEYINPUT63), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1130), .B(new_n1131), .C1(new_n1071), .C2(new_n1059), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1136), .B2(KEYINPUT63), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1138), .A2(KEYINPUT62), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1076), .B1(new_n1138), .B2(KEYINPUT62), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n1074), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1049), .A2(new_n1035), .A3(new_n804), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(G1981), .B2(G305), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1060), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1143), .A2(new_n1028), .B1(new_n1050), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1137), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1000), .B1(new_n1129), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n988), .B1(new_n730), .B2(new_n995), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT126), .Z(new_n1149));
  XNOR2_X1  g724(.A(new_n992), .B(KEYINPUT46), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT47), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n994), .A2(new_n997), .A3(new_n999), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n988), .A2(new_n989), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT48), .Z(new_n1155));
  OAI21_X1  g730(.A(new_n1152), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n994), .A2(new_n818), .A3(new_n821), .A4(new_n997), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(G2067), .B2(new_n782), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n988), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1147), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g735(.A1(new_n460), .A2(G227), .ZN(new_n1162));
  OAI21_X1  g736(.A(new_n1162), .B1(new_n664), .B2(new_n665), .ZN(new_n1163));
  XOR2_X1   g737(.A(new_n1163), .B(KEYINPUT127), .Z(new_n1164));
  NAND4_X1  g738(.A1(new_n1164), .A2(new_n895), .A3(new_n695), .A4(new_n969), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


