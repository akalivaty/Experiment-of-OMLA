

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n529, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776;

  INV_X1 U372 ( .A(KEYINPUT22), .ZN(n350) );
  NOR2_X1 U373 ( .A1(n712), .A2(n604), .ZN(n592) );
  OR2_X1 U374 ( .A1(n551), .A2(n560), .ZN(n728) );
  XNOR2_X1 U375 ( .A(n526), .B(n351), .ZN(n531) );
  XNOR2_X1 U376 ( .A(n527), .B(n352), .ZN(n351) );
  INV_X1 U377 ( .A(n529), .ZN(n352) );
  XNOR2_X1 U378 ( .A(G116), .B(G113), .ZN(n508) );
  XNOR2_X1 U379 ( .A(G128), .B(KEYINPUT24), .ZN(n493) );
  XNOR2_X1 U380 ( .A(G104), .B(G101), .ZN(n482) );
  AND2_X2 U381 ( .A1(n372), .A2(n410), .ZN(n409) );
  NAND2_X4 U382 ( .A1(G214), .A2(n474), .ZN(n725) );
  OR2_X2 U383 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X2 U384 ( .A1(n613), .A2(n432), .ZN(n431) );
  NOR2_X2 U385 ( .A1(n625), .A2(n632), .ZN(n620) );
  XNOR2_X2 U386 ( .A(n489), .B(KEYINPUT10), .ZN(n526) );
  NAND2_X1 U387 ( .A1(n574), .A2(n775), .ZN(n575) );
  NAND2_X1 U388 ( .A1(n458), .A2(n710), .ZN(n574) );
  INV_X2 U389 ( .A(n468), .ZN(n489) );
  INV_X1 U390 ( .A(n386), .ZN(n565) );
  NAND2_X1 U391 ( .A1(n386), .A2(n562), .ZN(n554) );
  XNOR2_X2 U392 ( .A(n553), .B(n350), .ZN(n386) );
  XNOR2_X2 U393 ( .A(n660), .B(KEYINPUT59), .ZN(n661) );
  NAND2_X4 U394 ( .A1(n560), .A2(n551), .ZN(n368) );
  XOR2_X2 U395 ( .A(KEYINPUT15), .B(G902), .Z(n640) );
  XNOR2_X1 U396 ( .A(KEYINPUT5), .B(G137), .ZN(n434) );
  XNOR2_X1 U397 ( .A(KEYINPUT76), .B(G107), .ZN(n485) );
  XNOR2_X1 U398 ( .A(n405), .B(KEYINPUT33), .ZN(n418) );
  XNOR2_X1 U399 ( .A(n550), .B(n549), .ZN(n555) );
  NAND2_X1 U400 ( .A1(n413), .A2(n411), .ZN(n550) );
  XNOR2_X1 U401 ( .A(n450), .B(n358), .ZN(n357) );
  NOR2_X1 U402 ( .A1(n723), .A2(n609), .ZN(n612) );
  INV_X1 U403 ( .A(n418), .ZN(n412) );
  XNOR2_X1 U404 ( .A(n404), .B(KEYINPUT98), .ZN(n720) );
  AND2_X1 U405 ( .A1(n712), .A2(n713), .ZN(n708) );
  XNOR2_X1 U406 ( .A(n532), .B(n531), .ZN(n660) );
  INV_X1 U407 ( .A(KEYINPUT97), .ZN(n358) );
  INV_X1 U408 ( .A(n698), .ZN(n445) );
  INV_X1 U409 ( .A(n357), .ZN(n675) );
  NAND2_X1 U410 ( .A1(n361), .A2(n389), .ZN(n449) );
  XNOR2_X1 U411 ( .A(n606), .B(KEYINPUT40), .ZN(n776) );
  AND2_X1 U412 ( .A1(n437), .A2(n369), .ZN(n415) );
  AND2_X1 U413 ( .A1(n638), .A2(n685), .ZN(n606) );
  XNOR2_X1 U414 ( .A(n427), .B(KEYINPUT39), .ZN(n638) );
  NAND2_X1 U415 ( .A1(n514), .A2(n403), .ZN(n405) );
  AND2_X1 U416 ( .A1(n571), .A2(n562), .ZN(n385) );
  NOR2_X1 U417 ( .A1(n605), .A2(n604), .ZN(n622) );
  OR2_X1 U418 ( .A1(G902), .A2(n745), .ZN(n544) );
  AND2_X1 U419 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U420 ( .A(n443), .B(n484), .ZN(n442) );
  XNOR2_X1 U421 ( .A(n526), .B(n491), .ZN(n762) );
  XNOR2_X1 U422 ( .A(n356), .B(n353), .ZN(n443) );
  XNOR2_X1 U423 ( .A(n516), .B(G134), .ZN(n455) );
  XNOR2_X1 U424 ( .A(n490), .B(n485), .ZN(n353) );
  XNOR2_X1 U425 ( .A(n435), .B(n434), .ZN(n433) );
  XNOR2_X1 U426 ( .A(n548), .B(KEYINPUT35), .ZN(n549) );
  XOR2_X1 U427 ( .A(n547), .B(KEYINPUT34), .Z(n369) );
  XNOR2_X2 U428 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n465) );
  XNOR2_X1 U429 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n435) );
  XNOR2_X2 U430 ( .A(G119), .B(G110), .ZN(n492) );
  XOR2_X2 U431 ( .A(G113), .B(G104), .Z(n527) );
  XOR2_X2 U432 ( .A(G146), .B(G125), .Z(n468) );
  INV_X2 U433 ( .A(KEYINPUT66), .ZN(n480) );
  NAND2_X1 U434 ( .A1(n668), .A2(n488), .ZN(n384) );
  XNOR2_X2 U435 ( .A(n442), .B(n512), .ZN(n668) );
  XNOR2_X2 U436 ( .A(n402), .B(n401), .ZN(n514) );
  XNOR2_X1 U437 ( .A(n455), .B(n354), .ZN(n764) );
  XNOR2_X1 U438 ( .A(n354), .B(n472), .ZN(n419) );
  XNOR2_X2 U439 ( .A(n538), .B(KEYINPUT4), .ZN(n354) );
  XNOR2_X1 U440 ( .A(n377), .B(KEYINPUT92), .ZN(n355) );
  XNOR2_X1 U441 ( .A(n377), .B(KEYINPUT92), .ZN(n437) );
  BUF_X1 U442 ( .A(n486), .Z(n356) );
  INV_X1 U443 ( .A(KEYINPUT72), .ZN(n401) );
  XOR2_X1 U444 ( .A(n635), .B(KEYINPUT38), .Z(n726) );
  AND2_X2 U445 ( .A1(n430), .A2(n364), .ZN(n359) );
  XNOR2_X1 U446 ( .A(n575), .B(KEYINPUT85), .ZN(n580) );
  INV_X1 U447 ( .A(n776), .ZN(n421) );
  XNOR2_X1 U448 ( .A(G143), .B(G122), .ZN(n515) );
  XOR2_X1 U449 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n518) );
  OR2_X1 U450 ( .A1(G237), .A2(G902), .ZN(n474) );
  AND2_X1 U451 ( .A1(n359), .A2(KEYINPUT2), .ZN(n426) );
  OR2_X2 U452 ( .A1(n749), .A2(G902), .ZN(n388) );
  NAND2_X1 U453 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U454 ( .A(n512), .B(n513), .ZN(n653) );
  XNOR2_X1 U455 ( .A(n436), .B(n433), .ZN(n511) );
  INV_X2 U456 ( .A(G140), .ZN(n483) );
  NAND2_X1 U457 ( .A1(n623), .A2(n428), .ZN(n427) );
  AND2_X1 U458 ( .A1(n622), .A2(n726), .ZN(n428) );
  NOR2_X1 U459 ( .A1(G953), .A2(G237), .ZN(n521) );
  NAND2_X1 U460 ( .A1(n514), .A2(n716), .ZN(n404) );
  INV_X1 U461 ( .A(G902), .ZN(n380) );
  XNOR2_X1 U462 ( .A(n508), .B(KEYINPUT73), .ZN(n436) );
  XNOR2_X1 U463 ( .A(n420), .B(KEYINPUT46), .ZN(n613) );
  NAND2_X1 U464 ( .A1(n422), .A2(n421), .ZN(n420) );
  INV_X1 U465 ( .A(KEYINPUT99), .ZN(n529) );
  XNOR2_X1 U466 ( .A(G140), .B(KEYINPUT12), .ZN(n517) );
  INV_X1 U467 ( .A(KEYINPUT82), .ZN(n440) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n477) );
  NAND2_X1 U469 ( .A1(n412), .A2(n369), .ZN(n411) );
  INV_X1 U470 ( .A(KEYINPUT31), .ZN(n394) );
  INV_X1 U471 ( .A(KEYINPUT16), .ZN(n441) );
  AND2_X1 U472 ( .A1(n359), .A2(n371), .ZN(n446) );
  XNOR2_X1 U473 ( .A(n454), .B(n453), .ZN(n723) );
  XNOR2_X1 U474 ( .A(n607), .B(n608), .ZN(n453) );
  NOR2_X1 U475 ( .A1(n729), .A2(n728), .ZN(n454) );
  XNOR2_X1 U476 ( .A(n373), .B(n475), .ZN(n597) );
  XNOR2_X1 U477 ( .A(n603), .B(n429), .ZN(n623) );
  INV_X1 U478 ( .A(KEYINPUT30), .ZN(n429) );
  XNOR2_X1 U479 ( .A(n716), .B(KEYINPUT6), .ZN(n616) );
  XNOR2_X1 U480 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U481 ( .A(n649), .B(n648), .ZN(n752) );
  INV_X1 U482 ( .A(n449), .ZN(n690) );
  NOR2_X1 U483 ( .A1(n716), .A2(n554), .ZN(n458) );
  XOR2_X1 U484 ( .A(KEYINPUT87), .B(KEYINPUT0), .Z(n360) );
  AND2_X1 U485 ( .A1(n393), .A2(n392), .ZN(n361) );
  AND2_X1 U486 ( .A1(n602), .A2(n601), .ZN(n362) );
  XOR2_X1 U487 ( .A(n504), .B(KEYINPUT25), .Z(n363) );
  AND2_X1 U488 ( .A1(n639), .A2(n696), .ZN(n364) );
  OR2_X1 U489 ( .A1(n479), .A2(n360), .ZN(n365) );
  NOR2_X1 U490 ( .A1(n412), .A2(n733), .ZN(n366) );
  NOR2_X1 U491 ( .A1(n723), .A2(n412), .ZN(n367) );
  NAND2_X1 U492 ( .A1(n640), .A2(KEYINPUT2), .ZN(n370) );
  AND2_X1 U493 ( .A1(KEYINPUT2), .A2(n448), .ZN(n371) );
  INV_X1 U494 ( .A(KEYINPUT74), .ZN(n448) );
  NAND2_X1 U495 ( .A1(n597), .A2(n360), .ZN(n372) );
  NAND2_X1 U496 ( .A1(n614), .A2(n725), .ZN(n373) );
  XNOR2_X1 U497 ( .A(n557), .B(KEYINPUT1), .ZN(n374) );
  XNOR2_X1 U498 ( .A(n557), .B(KEYINPUT1), .ZN(n631) );
  NAND2_X2 U499 ( .A1(n382), .A2(n378), .ZN(n557) );
  BUF_X1 U500 ( .A(n597), .Z(n375) );
  NAND2_X1 U501 ( .A1(n391), .A2(n390), .ZN(n389) );
  NAND2_X2 U502 ( .A1(n409), .A2(n408), .ZN(n377) );
  BUF_X1 U503 ( .A(n614), .Z(n635) );
  BUF_X1 U504 ( .A(n666), .Z(n748) );
  XNOR2_X1 U505 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X2 U506 ( .A1(n609), .A2(n375), .ZN(n686) );
  OR2_X1 U507 ( .A1(n597), .A2(n365), .ZN(n408) );
  INV_X1 U508 ( .A(n700), .ZN(n376) );
  NOR2_X1 U509 ( .A1(n377), .A2(n728), .ZN(n552) );
  NOR2_X1 U510 ( .A1(n377), .A2(n394), .ZN(n390) );
  NAND2_X1 U511 ( .A1(n377), .A2(n394), .ZN(n392) );
  OR2_X1 U512 ( .A1(n668), .A2(n379), .ZN(n378) );
  INV_X1 U513 ( .A(n488), .ZN(n381) );
  NAND2_X1 U514 ( .A1(n488), .A2(G902), .ZN(n383) );
  NAND2_X1 U515 ( .A1(n386), .A2(n385), .ZN(n573) );
  XNOR2_X2 U516 ( .A(n387), .B(n407), .ZN(n644) );
  XNOR2_X2 U517 ( .A(n452), .B(n451), .ZN(n387) );
  XNOR2_X1 U518 ( .A(n387), .B(KEYINPUT125), .ZN(n758) );
  NAND2_X1 U519 ( .A1(n644), .A2(n501), .ZN(n406) );
  INV_X2 U520 ( .A(KEYINPUT91), .ZN(n397) );
  INV_X2 U521 ( .A(G119), .ZN(n400) );
  INV_X1 U522 ( .A(n616), .ZN(n403) );
  NAND2_X1 U523 ( .A1(n631), .A2(n708), .ZN(n402) );
  XNOR2_X2 U524 ( .A(n388), .B(n363), .ZN(n712) );
  INV_X1 U525 ( .A(n720), .ZN(n391) );
  NAND2_X1 U526 ( .A1(n720), .A2(n394), .ZN(n393) );
  NAND2_X1 U527 ( .A1(n395), .A2(n561), .ZN(n566) );
  NAND2_X1 U528 ( .A1(n357), .A2(n449), .ZN(n395) );
  XNOR2_X2 U529 ( .A(n396), .B(G472), .ZN(n716) );
  NAND2_X1 U530 ( .A1(n653), .A2(n380), .ZN(n396) );
  XNOR2_X2 U531 ( .A(n397), .B(G110), .ZN(n486) );
  XNOR2_X2 U532 ( .A(n509), .B(n398), .ZN(n452) );
  XNOR2_X2 U533 ( .A(n486), .B(n441), .ZN(n398) );
  XNOR2_X2 U534 ( .A(n399), .B(n460), .ZN(n509) );
  XNOR2_X2 U535 ( .A(n400), .B(G101), .ZN(n399) );
  NOR2_X1 U536 ( .A1(n355), .A2(n369), .ZN(n417) );
  XNOR2_X2 U537 ( .A(n406), .B(n457), .ZN(n614) );
  XNOR2_X1 U538 ( .A(n419), .B(n473), .ZN(n407) );
  NAND2_X1 U539 ( .A1(n479), .A2(n360), .ZN(n410) );
  AND2_X2 U540 ( .A1(n414), .A2(n416), .ZN(n413) );
  NOR2_X1 U541 ( .A1(n415), .A2(n368), .ZN(n414) );
  NAND2_X1 U542 ( .A1(n418), .A2(n417), .ZN(n416) );
  INV_X1 U543 ( .A(n773), .ZN(n422) );
  XNOR2_X1 U544 ( .A(n587), .B(n440), .ZN(n439) );
  NAND2_X1 U545 ( .A1(n423), .A2(KEYINPUT74), .ZN(n425) );
  NAND2_X1 U546 ( .A1(n445), .A2(n426), .ZN(n423) );
  XNOR2_X2 U547 ( .A(n424), .B(n641), .ZN(n666) );
  NAND2_X1 U548 ( .A1(n447), .A2(n697), .ZN(n424) );
  NAND2_X1 U549 ( .A1(n425), .A2(n444), .ZN(n697) );
  XNOR2_X1 U550 ( .A(n431), .B(n630), .ZN(n430) );
  NAND2_X1 U551 ( .A1(n362), .A2(n628), .ZN(n432) );
  OR2_X1 U552 ( .A1(n355), .A2(n558), .ZN(n450) );
  NAND2_X1 U553 ( .A1(n438), .A2(n370), .ZN(n447) );
  NAND2_X1 U554 ( .A1(n439), .A2(n359), .ZN(n438) );
  XNOR2_X2 U555 ( .A(n764), .B(G146), .ZN(n512) );
  NAND2_X1 U556 ( .A1(n445), .A2(n446), .ZN(n444) );
  XNOR2_X2 U557 ( .A(n536), .B(n527), .ZN(n451) );
  XNOR2_X2 U558 ( .A(n459), .B(G122), .ZN(n536) );
  BUF_X1 U559 ( .A(n555), .Z(n578) );
  AND2_X1 U560 ( .A1(n374), .A2(n616), .ZN(n571) );
  AND2_X1 U561 ( .A1(n521), .A2(G210), .ZN(n456) );
  AND2_X1 U562 ( .A1(G210), .A2(n474), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n516), .B(n515), .ZN(n520) );
  XNOR2_X1 U564 ( .A(n509), .B(n456), .ZN(n510) );
  XNOR2_X1 U565 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U566 ( .A(n629), .B(KEYINPUT67), .ZN(n630) );
  INV_X1 U567 ( .A(n490), .ZN(n491) );
  INV_X1 U568 ( .A(n640), .ZN(n501) );
  XNOR2_X2 U569 ( .A(G116), .B(G107), .ZN(n459) );
  XNOR2_X2 U570 ( .A(KEYINPUT70), .B(KEYINPUT3), .ZN(n460) );
  INV_X1 U571 ( .A(KEYINPUT17), .ZN(n461) );
  NAND2_X1 U572 ( .A1(n461), .A2(KEYINPUT18), .ZN(n464) );
  INV_X1 U573 ( .A(KEYINPUT18), .ZN(n462) );
  NAND2_X1 U574 ( .A1(n462), .A2(KEYINPUT17), .ZN(n463) );
  NAND2_X1 U575 ( .A1(n464), .A2(n463), .ZN(n466) );
  XNOR2_X1 U576 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U577 ( .A1(n467), .A2(n489), .ZN(n471) );
  INV_X1 U578 ( .A(n467), .ZN(n469) );
  NAND2_X1 U579 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U580 ( .A1(n471), .A2(n470), .ZN(n473) );
  INV_X2 U581 ( .A(G953), .ZN(n769) );
  NAND2_X1 U582 ( .A1(G224), .A2(n769), .ZN(n472) );
  XNOR2_X2 U583 ( .A(G143), .B(G128), .ZN(n538) );
  INV_X1 U584 ( .A(KEYINPUT19), .ZN(n475) );
  NOR2_X1 U585 ( .A1(G898), .A2(n769), .ZN(n759) );
  NAND2_X1 U586 ( .A1(n759), .A2(G902), .ZN(n476) );
  NAND2_X1 U587 ( .A1(G952), .A2(n769), .ZN(n589) );
  NAND2_X1 U588 ( .A1(n476), .A2(n589), .ZN(n478) );
  XNOR2_X1 U589 ( .A(n477), .B(KEYINPUT14), .ZN(n706) );
  NAND2_X1 U590 ( .A1(n478), .A2(n706), .ZN(n479) );
  XNOR2_X2 U591 ( .A(n480), .B(G131), .ZN(n516) );
  AND2_X1 U592 ( .A1(n769), .A2(G227), .ZN(n481) );
  XNOR2_X1 U593 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U594 ( .A(n483), .B(G137), .ZN(n490) );
  INV_X1 U595 ( .A(KEYINPUT69), .ZN(n487) );
  XNOR2_X1 U596 ( .A(n487), .B(G469), .ZN(n488) );
  XOR2_X1 U597 ( .A(n492), .B(KEYINPUT75), .Z(n496) );
  XOR2_X1 U598 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n494) );
  XNOR2_X1 U599 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U600 ( .A(n496), .B(n495), .ZN(n499) );
  NAND2_X1 U601 ( .A1(G234), .A2(n769), .ZN(n497) );
  XOR2_X1 U602 ( .A(KEYINPUT8), .B(n497), .Z(n537) );
  NAND2_X1 U603 ( .A1(G221), .A2(n537), .ZN(n498) );
  XNOR2_X1 U604 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U605 ( .A(n762), .B(n500), .ZN(n749) );
  NAND2_X1 U606 ( .A1(n501), .A2(G234), .ZN(n503) );
  XNOR2_X1 U607 ( .A(KEYINPUT20), .B(KEYINPUT94), .ZN(n502) );
  XNOR2_X1 U608 ( .A(n503), .B(n502), .ZN(n505) );
  NAND2_X1 U609 ( .A1(G217), .A2(n505), .ZN(n504) );
  NAND2_X1 U610 ( .A1(n505), .A2(G221), .ZN(n507) );
  INV_X1 U611 ( .A(KEYINPUT21), .ZN(n506) );
  XNOR2_X1 U612 ( .A(n507), .B(n506), .ZN(n713) );
  XNOR2_X1 U613 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U614 ( .A(n520), .B(n519), .ZN(n525) );
  XOR2_X1 U615 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n523) );
  NAND2_X1 U616 ( .A1(G214), .A2(n521), .ZN(n522) );
  XNOR2_X1 U617 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U618 ( .A(n525), .B(n524), .ZN(n532) );
  NAND2_X1 U619 ( .A1(n660), .A2(n380), .ZN(n534) );
  XOR2_X1 U620 ( .A(KEYINPUT13), .B(G475), .Z(n533) );
  XNOR2_X1 U621 ( .A(n534), .B(n533), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n535) );
  XNOR2_X1 U623 ( .A(G478), .B(n535), .ZN(n545) );
  XNOR2_X1 U624 ( .A(G134), .B(KEYINPUT7), .ZN(n542) );
  NAND2_X1 U625 ( .A1(G217), .A2(n537), .ZN(n540) );
  XNOR2_X1 U626 ( .A(n538), .B(KEYINPUT9), .ZN(n539) );
  XNOR2_X1 U627 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U628 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U629 ( .A(n536), .B(n543), .ZN(n745) );
  XNOR2_X1 U630 ( .A(n545), .B(n544), .ZN(n551) );
  INV_X1 U631 ( .A(n551), .ZN(n559) );
  NAND2_X1 U632 ( .A1(n560), .A2(n559), .ZN(n618) );
  INV_X1 U633 ( .A(n618), .ZN(n685) );
  NAND2_X1 U634 ( .A1(n690), .A2(n685), .ZN(n546) );
  XNOR2_X1 U635 ( .A(n546), .B(G113), .ZN(G15) );
  INV_X1 U636 ( .A(KEYINPUT80), .ZN(n547) );
  INV_X1 U637 ( .A(KEYINPUT79), .ZN(n548) );
  XOR2_X1 U638 ( .A(n578), .B(G122), .Z(G24) );
  NAND2_X1 U639 ( .A1(n552), .A2(n713), .ZN(n553) );
  INV_X1 U640 ( .A(n374), .ZN(n710) );
  XNOR2_X1 U641 ( .A(n574), .B(G110), .ZN(G12) );
  NAND2_X1 U642 ( .A1(n555), .A2(KEYINPUT44), .ZN(n556) );
  XNOR2_X1 U643 ( .A(n556), .B(KEYINPUT84), .ZN(n569) );
  NAND2_X1 U644 ( .A1(n708), .A2(n557), .ZN(n605) );
  OR2_X1 U645 ( .A1(n605), .A2(n716), .ZN(n558) );
  OR2_X1 U646 ( .A1(n560), .A2(n559), .ZN(n637) );
  AND2_X1 U647 ( .A1(n618), .A2(n637), .ZN(n730) );
  INV_X1 U648 ( .A(n730), .ZN(n561) );
  INV_X1 U649 ( .A(n712), .ZN(n562) );
  NOR2_X1 U650 ( .A1(n374), .A2(n562), .ZN(n563) );
  NAND2_X1 U651 ( .A1(n616), .A2(n563), .ZN(n564) );
  OR2_X1 U652 ( .A1(n565), .A2(n564), .ZN(n672) );
  NAND2_X1 U653 ( .A1(n566), .A2(n672), .ZN(n567) );
  XNOR2_X1 U654 ( .A(n567), .B(KEYINPUT105), .ZN(n568) );
  NAND2_X1 U655 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U656 ( .A(n570), .B(KEYINPUT83), .ZN(n585) );
  XOR2_X1 U657 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n572) );
  XNOR2_X1 U658 ( .A(n573), .B(n572), .ZN(n775) );
  INV_X1 U659 ( .A(n580), .ZN(n577) );
  INV_X1 U660 ( .A(KEYINPUT44), .ZN(n576) );
  NAND2_X1 U661 ( .A1(n577), .A2(n576), .ZN(n583) );
  INV_X1 U662 ( .A(n578), .ZN(n579) );
  NAND2_X1 U663 ( .A1(n579), .A2(n576), .ZN(n581) );
  NAND2_X1 U664 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U665 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U666 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X2 U667 ( .A(n586), .B(KEYINPUT45), .ZN(n753) );
  NAND2_X1 U668 ( .A1(n753), .A2(n640), .ZN(n587) );
  NOR2_X1 U669 ( .A1(n730), .A2(KEYINPUT71), .ZN(n598) );
  NOR2_X1 U670 ( .A1(G900), .A2(n769), .ZN(n588) );
  NAND2_X1 U671 ( .A1(n588), .A2(G902), .ZN(n590) );
  NAND2_X1 U672 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n591), .A2(n706), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n713), .A2(n592), .ZN(n593) );
  XNOR2_X1 U675 ( .A(KEYINPUT68), .B(n593), .ZN(n615) );
  INV_X1 U676 ( .A(n716), .ZN(n594) );
  NOR2_X1 U677 ( .A1(n615), .A2(n594), .ZN(n595) );
  XNOR2_X1 U678 ( .A(KEYINPUT28), .B(n595), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n596), .A2(n557), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n598), .A2(n686), .ZN(n599) );
  XOR2_X1 U681 ( .A(n599), .B(KEYINPUT47), .Z(n602) );
  AND2_X1 U682 ( .A1(n730), .A2(KEYINPUT71), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n600), .A2(n686), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n716), .A2(n725), .ZN(n603) );
  INV_X1 U685 ( .A(KEYINPUT108), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n726), .A2(n725), .ZN(n729) );
  XNOR2_X1 U687 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n607) );
  XOR2_X1 U688 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n610) );
  XNOR2_X1 U689 ( .A(KEYINPUT110), .B(n610), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n612), .B(n611), .ZN(n773) );
  INV_X1 U691 ( .A(n635), .ZN(n625) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n619), .A2(n725), .ZN(n632) );
  XOR2_X1 U694 ( .A(KEYINPUT36), .B(n620), .Z(n621) );
  NOR2_X1 U695 ( .A1(n621), .A2(n710), .ZN(n693) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n626), .B(KEYINPUT107), .ZN(n627) );
  NOR2_X1 U699 ( .A1(n627), .A2(n368), .ZN(n684) );
  NOR2_X1 U700 ( .A1(n693), .A2(n684), .ZN(n628) );
  INV_X1 U701 ( .A(KEYINPUT48), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n632), .A2(n374), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n633), .B(KEYINPUT43), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U705 ( .A(KEYINPUT106), .B(n636), .ZN(n774) );
  INV_X1 U706 ( .A(n774), .ZN(n639) );
  INV_X1 U707 ( .A(n637), .ZN(n689) );
  NAND2_X1 U708 ( .A1(n638), .A2(n689), .ZN(n696) );
  INV_X1 U709 ( .A(n753), .ZN(n698) );
  INV_X1 U710 ( .A(KEYINPUT2), .ZN(n699) );
  INV_X1 U711 ( .A(KEYINPUT64), .ZN(n641) );
  NAND2_X1 U712 ( .A1(n666), .A2(G210), .ZN(n646) );
  XNOR2_X1 U713 ( .A(KEYINPUT86), .B(KEYINPUT54), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n642), .B(KEYINPUT55), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(n650) );
  INV_X1 U716 ( .A(G952), .ZN(n647) );
  NAND2_X1 U717 ( .A1(n647), .A2(G953), .ZN(n649) );
  INV_X1 U718 ( .A(KEYINPUT90), .ZN(n648) );
  NOR2_X2 U719 ( .A1(n650), .A2(n752), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U721 ( .A1(n666), .A2(G472), .ZN(n655) );
  XOR2_X1 U722 ( .A(KEYINPUT88), .B(KEYINPUT62), .Z(n652) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U724 ( .A1(n656), .A2(n752), .ZN(n659) );
  XNOR2_X1 U725 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n657), .B(KEYINPUT89), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(G57) );
  NAND2_X1 U728 ( .A1(n666), .A2(G475), .ZN(n662) );
  XNOR2_X1 U729 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X2 U730 ( .A1(n663), .A2(n752), .ZN(n665) );
  XNOR2_X1 U731 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n665), .B(n664), .ZN(G60) );
  NAND2_X1 U733 ( .A1(n748), .A2(G469), .ZN(n670) );
  XOR2_X1 U734 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U737 ( .A1(n671), .A2(n752), .ZN(G54) );
  XOR2_X1 U738 ( .A(n672), .B(G101), .Z(n673) );
  XNOR2_X1 U739 ( .A(n673), .B(KEYINPUT113), .ZN(G3) );
  NAND2_X1 U740 ( .A1(n675), .A2(n685), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n674), .B(G104), .ZN(G6) );
  XNOR2_X1 U742 ( .A(G107), .B(KEYINPUT27), .ZN(n679) );
  XOR2_X1 U743 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n677) );
  NAND2_X1 U744 ( .A1(n675), .A2(n689), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n679), .B(n678), .ZN(G9) );
  XOR2_X1 U747 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n681) );
  NAND2_X1 U748 ( .A1(n686), .A2(n689), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(n683) );
  XOR2_X1 U750 ( .A(G128), .B(KEYINPUT115), .Z(n682) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(G30) );
  XOR2_X1 U752 ( .A(G143), .B(n684), .Z(G45) );
  XOR2_X1 U753 ( .A(G146), .B(KEYINPUT117), .Z(n688) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n688), .B(n687), .ZN(G48) );
  NAND2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n691), .B(KEYINPUT118), .ZN(n692) );
  XNOR2_X1 U758 ( .A(G116), .B(n692), .ZN(G18) );
  XNOR2_X1 U759 ( .A(n693), .B(G125), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n694), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U761 ( .A(G134), .B(KEYINPUT119), .Z(n695) );
  XNOR2_X1 U762 ( .A(n696), .B(n695), .ZN(G36) );
  INV_X1 U763 ( .A(n697), .ZN(n705) );
  BUF_X1 U764 ( .A(n698), .Z(n700) );
  NAND2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n703) );
  NOR2_X1 U766 ( .A1(KEYINPUT2), .A2(n359), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n701), .B(KEYINPUT81), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n742) );
  NAND2_X1 U770 ( .A1(G952), .A2(n706), .ZN(n737) );
  XNOR2_X1 U771 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n707), .B(KEYINPUT51), .ZN(n722) );
  INV_X1 U773 ( .A(n708), .ZN(n709) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U775 ( .A(n711), .B(KEYINPUT50), .ZN(n718) );
  NOR2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U777 ( .A(KEYINPUT49), .B(n714), .Z(n715) );
  NOR2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U779 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U781 ( .A(n722), .B(n721), .Z(n724) );
  NOR2_X1 U782 ( .A1(n724), .A2(n723), .ZN(n734) );
  NOR2_X1 U783 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U784 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U785 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U787 ( .A1(n734), .A2(n366), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n735), .B(KEYINPUT52), .ZN(n736) );
  NOR2_X1 U789 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U790 ( .A(n738), .B(KEYINPUT122), .ZN(n739) );
  NOR2_X1 U791 ( .A1(n739), .A2(n367), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT123), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U794 ( .A1(n769), .A2(n743), .ZN(n744) );
  XOR2_X1 U795 ( .A(KEYINPUT53), .B(n744), .Z(G75) );
  NAND2_X1 U796 ( .A1(n748), .A2(G478), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U798 ( .A1(n752), .A2(n747), .ZN(G63) );
  NAND2_X1 U799 ( .A1(n748), .A2(G217), .ZN(n750) );
  XNOR2_X1 U800 ( .A(n749), .B(n750), .ZN(n751) );
  NOR2_X1 U801 ( .A1(n752), .A2(n751), .ZN(G66) );
  NAND2_X1 U802 ( .A1(n376), .A2(n769), .ZN(n757) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n754) );
  XNOR2_X1 U804 ( .A(KEYINPUT61), .B(n754), .ZN(n755) );
  NAND2_X1 U805 ( .A1(n755), .A2(G898), .ZN(n756) );
  NAND2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n761) );
  NOR2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U808 ( .A(n761), .B(n760), .ZN(G69) );
  XNOR2_X1 U809 ( .A(n762), .B(KEYINPUT126), .ZN(n763) );
  XOR2_X1 U810 ( .A(n764), .B(n763), .Z(n768) );
  XNOR2_X1 U811 ( .A(n768), .B(KEYINPUT127), .ZN(n765) );
  XNOR2_X1 U812 ( .A(G227), .B(n765), .ZN(n766) );
  NAND2_X1 U813 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U814 ( .A1(n767), .A2(G953), .ZN(n772) );
  XNOR2_X1 U815 ( .A(n359), .B(n768), .ZN(n770) );
  NAND2_X1 U816 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U817 ( .A1(n772), .A2(n771), .ZN(G72) );
  XOR2_X1 U818 ( .A(G137), .B(n773), .Z(G39) );
  XOR2_X1 U819 ( .A(G140), .B(n774), .Z(G42) );
  XNOR2_X1 U820 ( .A(n775), .B(G119), .ZN(G21) );
  XOR2_X1 U821 ( .A(G131), .B(n776), .Z(G33) );
endmodule

