

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757;

  INV_X4 U372 ( .A(G953), .ZN(n750) );
  OR2_X1 U373 ( .A1(n658), .A2(G902), .ZN(n426) );
  XNOR2_X2 U374 ( .A(n462), .B(KEYINPUT79), .ZN(n548) );
  NOR2_X2 U375 ( .A1(n521), .A2(n386), .ZN(n421) );
  XNOR2_X2 U376 ( .A(n586), .B(n585), .ZN(n724) );
  AND2_X1 U377 ( .A1(n734), .A2(n371), .ZN(n614) );
  OR2_X1 U378 ( .A1(n590), .A2(n589), .ZN(n592) );
  NOR2_X1 U379 ( .A1(n695), .A2(n692), .ZN(n512) );
  XNOR2_X1 U380 ( .A(KEYINPUT10), .B(G140), .ZN(n427) );
  AND2_X1 U381 ( .A1(n732), .A2(n750), .ZN(n733) );
  XNOR2_X1 U382 ( .A(n510), .B(n355), .ZN(n639) );
  XOR2_X1 U383 ( .A(KEYINPUT106), .B(n524), .Z(n553) );
  AND2_X1 U384 ( .A1(n518), .A2(n517), .ZN(n673) );
  AND2_X1 U385 ( .A1(n578), .A2(n523), .ZN(n524) );
  NOR2_X1 U386 ( .A1(n602), .A2(n459), .ZN(n460) );
  XNOR2_X1 U387 ( .A(n385), .B(n532), .ZN(n669) );
  AND2_X1 U388 ( .A1(n599), .A2(n597), .ZN(n584) );
  NAND2_X1 U389 ( .A1(n529), .A2(n597), .ZN(n602) );
  OR2_X1 U390 ( .A1(n551), .A2(n386), .ZN(n385) );
  XNOR2_X1 U391 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U392 ( .A1(n617), .A2(n616), .ZN(n350) );
  NAND2_X1 U393 ( .A1(n617), .A2(n616), .ZN(n619) );
  AND2_X1 U394 ( .A1(n619), .A2(n381), .ZN(n351) );
  AND2_X1 U395 ( .A1(n350), .A2(n381), .ZN(n352) );
  AND2_X1 U396 ( .A1(n619), .A2(n381), .ZN(n653) );
  BUF_X1 U397 ( .A(n548), .Z(n353) );
  XNOR2_X2 U398 ( .A(n354), .B(G472), .ZN(n521) );
  NOR2_X1 U399 ( .A1(n631), .A2(G902), .ZN(n354) );
  XNOR2_X2 U400 ( .A(n471), .B(n427), .ZN(n498) );
  XNOR2_X2 U401 ( .A(n469), .B(G134), .ZN(n483) );
  XNOR2_X2 U402 ( .A(n745), .B(n409), .ZN(n425) );
  XNOR2_X2 U403 ( .A(n483), .B(n408), .ZN(n745) );
  NAND2_X1 U404 ( .A1(n546), .A2(n369), .ZN(n368) );
  AND2_X1 U405 ( .A1(n547), .A2(n637), .ZN(n369) );
  XNOR2_X1 U406 ( .A(n378), .B(KEYINPUT48), .ZN(n377) );
  INV_X1 U407 ( .A(n629), .ZN(n402) );
  AND2_X1 U408 ( .A1(n389), .A2(n387), .ZN(n393) );
  NAND2_X1 U409 ( .A1(n388), .A2(n394), .ZN(n387) );
  NAND2_X1 U410 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U411 ( .A(n468), .B(n467), .ZN(n740) );
  XNOR2_X1 U412 ( .A(n400), .B(n359), .ZN(n560) );
  NOR2_X1 U413 ( .A1(n618), .A2(n620), .ZN(n363) );
  INV_X1 U414 ( .A(KEYINPUT46), .ZN(n379) );
  NAND2_X1 U415 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U416 ( .A(KEYINPUT44), .ZN(n396) );
  NAND2_X1 U417 ( .A1(n398), .A2(n397), .ZN(n388) );
  INV_X1 U418 ( .A(KEYINPUT89), .ZN(n397) );
  AND2_X1 U419 ( .A1(n627), .A2(n626), .ZN(n593) );
  XNOR2_X1 U420 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n464) );
  XOR2_X1 U421 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n438) );
  INV_X1 U422 ( .A(KEYINPUT2), .ZN(n371) );
  XNOR2_X1 U423 ( .A(G107), .B(KEYINPUT7), .ZN(n485) );
  XOR2_X1 U424 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n486) );
  XOR2_X1 U425 ( .A(n525), .B(KEYINPUT38), .Z(n689) );
  NAND2_X1 U426 ( .A1(n402), .A2(n401), .ZN(n376) );
  XNOR2_X1 U427 ( .A(G128), .B(G110), .ZN(n432) );
  XNOR2_X1 U428 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n429) );
  XOR2_X1 U429 ( .A(G122), .B(G104), .Z(n501) );
  XNOR2_X1 U430 ( .A(n384), .B(n383), .ZN(n466) );
  XNOR2_X1 U431 ( .A(G107), .B(G104), .ZN(n384) );
  XNOR2_X1 U432 ( .A(KEYINPUT91), .B(G110), .ZN(n383) );
  OR2_X1 U433 ( .A1(n647), .A2(n381), .ZN(n482) );
  XNOR2_X1 U434 ( .A(n569), .B(n568), .ZN(n605) );
  INV_X1 U435 ( .A(KEYINPUT0), .ZN(n568) );
  NOR2_X1 U436 ( .A1(n669), .A2(n567), .ZN(n569) );
  NAND2_X1 U437 ( .A1(n380), .A2(n701), .ZN(n594) );
  NOR2_X1 U438 ( .A1(n618), .A2(n630), .ZN(n364) );
  NOR2_X2 U439 ( .A1(n560), .A2(n680), .ZN(n510) );
  NAND2_X1 U440 ( .A1(n550), .A2(n535), .ZN(n680) );
  INV_X1 U441 ( .A(n661), .ZN(n624) );
  XOR2_X1 U442 ( .A(n509), .B(KEYINPUT40), .Z(n355) );
  NAND2_X1 U443 ( .A1(n629), .A2(KEYINPUT87), .ZN(n356) );
  NOR2_X1 U444 ( .A1(n579), .A2(n578), .ZN(n357) );
  AND2_X1 U445 ( .A1(n376), .A2(n638), .ZN(n358) );
  XNOR2_X1 U446 ( .A(KEYINPUT73), .B(KEYINPUT39), .ZN(n359) );
  XNOR2_X1 U447 ( .A(n531), .B(KEYINPUT111), .ZN(n754) );
  XOR2_X1 U448 ( .A(n572), .B(KEYINPUT65), .Z(n360) );
  INV_X1 U449 ( .A(n618), .ZN(n381) );
  XOR2_X1 U450 ( .A(n621), .B(KEYINPUT124), .Z(n361) );
  AND2_X1 U451 ( .A1(KEYINPUT89), .A2(KEYINPUT44), .ZN(n362) );
  INV_X1 U452 ( .A(KEYINPUT87), .ZN(n401) );
  AND2_X1 U453 ( .A1(n350), .A2(n363), .ZN(n622) );
  AND2_X1 U454 ( .A1(n350), .A2(n364), .ZN(n633) );
  XNOR2_X1 U455 ( .A(n365), .B(n379), .ZN(n366) );
  NAND2_X1 U456 ( .A1(n639), .A2(n757), .ZN(n365) );
  XNOR2_X1 U457 ( .A(n520), .B(n519), .ZN(n757) );
  NAND2_X1 U458 ( .A1(n367), .A2(n366), .ZN(n378) );
  NOR2_X1 U459 ( .A1(n754), .A2(n368), .ZN(n367) );
  NAND2_X1 U460 ( .A1(n593), .A2(n370), .ZN(n611) );
  XNOR2_X1 U461 ( .A(n370), .B(G122), .ZN(G24) );
  XNOR2_X2 U462 ( .A(n592), .B(n591), .ZN(n370) );
  XNOR2_X2 U463 ( .A(n613), .B(KEYINPUT45), .ZN(n734) );
  AND2_X2 U464 ( .A1(n372), .A2(n358), .ZN(n749) );
  NAND2_X1 U465 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U466 ( .A1(n377), .A2(KEYINPUT87), .ZN(n373) );
  NAND2_X1 U467 ( .A1(n375), .A2(n356), .ZN(n374) );
  INV_X1 U468 ( .A(n377), .ZN(n375) );
  NAND2_X1 U469 ( .A1(n393), .A2(n390), .ZN(n612) );
  NAND2_X1 U470 ( .A1(n380), .A2(n357), .ZN(n583) );
  XNOR2_X1 U471 ( .A(n573), .B(n360), .ZN(n380) );
  XNOR2_X1 U472 ( .A(n740), .B(n382), .ZN(n647) );
  XNOR2_X1 U473 ( .A(n477), .B(n476), .ZN(n382) );
  INV_X1 U474 ( .A(n688), .ZN(n386) );
  NAND2_X1 U475 ( .A1(n611), .A2(n362), .ZN(n389) );
  AND2_X1 U476 ( .A1(n610), .A2(n397), .ZN(n391) );
  INV_X1 U477 ( .A(n611), .ZN(n392) );
  NAND2_X1 U478 ( .A1(n610), .A2(n395), .ZN(n394) );
  INV_X1 U479 ( .A(n610), .ZN(n398) );
  XNOR2_X2 U480 ( .A(n399), .B(G143), .ZN(n469) );
  XNOR2_X2 U481 ( .A(G128), .B(KEYINPUT82), .ZN(n399) );
  NAND2_X1 U482 ( .A1(n548), .A2(n689), .ZN(n400) );
  XNOR2_X1 U483 ( .A(n403), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U484 ( .A1(n404), .A2(n624), .ZN(n403) );
  XNOR2_X1 U485 ( .A(n622), .B(n361), .ZN(n404) );
  BUF_X1 U486 ( .A(n551), .Z(n558) );
  OR2_X1 U487 ( .A1(n611), .A2(KEYINPUT44), .ZN(n405) );
  AND2_X1 U488 ( .A1(n575), .A2(n570), .ZN(n597) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n658) );
  BUF_X1 U490 ( .A(n521), .Z(n704) );
  XNOR2_X1 U491 ( .A(KEYINPUT69), .B(G131), .ZN(n502) );
  INV_X1 U492 ( .A(KEYINPUT4), .ZN(n406) );
  XNOR2_X1 U493 ( .A(n406), .B(G137), .ZN(n407) );
  XNOR2_X1 U494 ( .A(n502), .B(n407), .ZN(n408) );
  XNOR2_X1 U495 ( .A(KEYINPUT66), .B(G101), .ZN(n474) );
  XNOR2_X1 U496 ( .A(n474), .B(G146), .ZN(n409) );
  NOR2_X1 U497 ( .A1(G953), .A2(G237), .ZN(n494) );
  AND2_X1 U498 ( .A1(n494), .A2(G210), .ZN(n411) );
  XNOR2_X1 U499 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n410) );
  XNOR2_X1 U500 ( .A(n411), .B(n410), .ZN(n416) );
  XNOR2_X1 U501 ( .A(G119), .B(G116), .ZN(n413) );
  XNOR2_X1 U502 ( .A(G113), .B(KEYINPUT70), .ZN(n412) );
  XNOR2_X1 U503 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U504 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n414) );
  XNOR2_X1 U505 ( .A(n415), .B(n414), .ZN(n467) );
  XNOR2_X1 U506 ( .A(n416), .B(n467), .ZN(n417) );
  XNOR2_X1 U507 ( .A(n425), .B(n417), .ZN(n631) );
  INV_X1 U508 ( .A(G472), .ZN(n630) );
  NOR2_X1 U509 ( .A1(G902), .A2(G237), .ZN(n419) );
  INV_X1 U510 ( .A(KEYINPUT77), .ZN(n418) );
  XNOR2_X1 U511 ( .A(n419), .B(n418), .ZN(n478) );
  INV_X1 U512 ( .A(G214), .ZN(n420) );
  OR2_X1 U513 ( .A1(n478), .A2(n420), .ZN(n688) );
  XNOR2_X1 U514 ( .A(n421), .B(KEYINPUT30), .ZN(n461) );
  NAND2_X1 U515 ( .A1(n750), .A2(G227), .ZN(n422) );
  XNOR2_X1 U516 ( .A(n422), .B(G140), .ZN(n423) );
  XNOR2_X1 U517 ( .A(n466), .B(n423), .ZN(n424) );
  XNOR2_X2 U518 ( .A(n426), .B(G469), .ZN(n529) );
  XNOR2_X2 U519 ( .A(G146), .B(G125), .ZN(n471) );
  INV_X1 U520 ( .A(G119), .ZN(n428) );
  XNOR2_X1 U521 ( .A(n428), .B(G137), .ZN(n430) );
  XNOR2_X1 U522 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U523 ( .A(n498), .B(n431), .ZN(n436) );
  XNOR2_X1 U524 ( .A(n432), .B(KEYINPUT80), .ZN(n434) );
  XNOR2_X1 U525 ( .A(KEYINPUT96), .B(KEYINPUT23), .ZN(n433) );
  XNOR2_X1 U526 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U527 ( .A(n436), .B(n435), .ZN(n442) );
  NAND2_X1 U528 ( .A1(G234), .A2(n750), .ZN(n437) );
  XNOR2_X1 U529 ( .A(n438), .B(n437), .ZN(n440) );
  INV_X1 U530 ( .A(KEYINPUT68), .ZN(n439) );
  XNOR2_X1 U531 ( .A(n440), .B(n439), .ZN(n484) );
  NAND2_X1 U532 ( .A1(n484), .A2(G221), .ZN(n441) );
  XNOR2_X1 U533 ( .A(n442), .B(n441), .ZN(n654) );
  OR2_X1 U534 ( .A1(n654), .A2(G902), .ZN(n447) );
  XNOR2_X1 U535 ( .A(KEYINPUT15), .B(G902), .ZN(n618) );
  NAND2_X1 U536 ( .A1(n618), .A2(G234), .ZN(n443) );
  XNOR2_X1 U537 ( .A(n443), .B(KEYINPUT20), .ZN(n448) );
  NAND2_X1 U538 ( .A1(n448), .A2(G217), .ZN(n445) );
  XNOR2_X1 U539 ( .A(KEYINPUT97), .B(KEYINPUT25), .ZN(n444) );
  XNOR2_X1 U540 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U541 ( .A(n447), .B(n446), .ZN(n575) );
  INV_X1 U542 ( .A(n448), .ZN(n450) );
  INV_X1 U543 ( .A(G221), .ZN(n449) );
  OR2_X1 U544 ( .A1(n450), .A2(n449), .ZN(n452) );
  INV_X1 U545 ( .A(KEYINPUT21), .ZN(n451) );
  XNOR2_X1 U546 ( .A(n452), .B(n451), .ZN(n570) );
  NAND2_X1 U547 ( .A1(G234), .A2(G237), .ZN(n453) );
  XNOR2_X1 U548 ( .A(n453), .B(KEYINPUT14), .ZN(n457) );
  NAND2_X1 U549 ( .A1(G902), .A2(n457), .ZN(n454) );
  XOR2_X1 U550 ( .A(KEYINPUT92), .B(n454), .Z(n455) );
  NAND2_X1 U551 ( .A1(G953), .A2(n455), .ZN(n561) );
  XOR2_X1 U552 ( .A(KEYINPUT105), .B(n561), .Z(n456) );
  OR2_X1 U553 ( .A1(n456), .A2(G900), .ZN(n458) );
  NAND2_X1 U554 ( .A1(G952), .A2(n457), .ZN(n721) );
  OR2_X1 U555 ( .A1(n721), .A2(G953), .ZN(n563) );
  NAND2_X1 U556 ( .A1(n458), .A2(n563), .ZN(n513) );
  INV_X1 U557 ( .A(n513), .ZN(n459) );
  NAND2_X1 U558 ( .A1(n461), .A2(n460), .ZN(n462) );
  INV_X1 U559 ( .A(G122), .ZN(n463) );
  XNOR2_X1 U560 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U561 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U562 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n470) );
  XNOR2_X1 U563 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U564 ( .A(n469), .B(n472), .ZN(n477) );
  NAND2_X1 U565 ( .A1(n750), .A2(G224), .ZN(n473) );
  XNOR2_X1 U566 ( .A(n473), .B(KEYINPUT4), .ZN(n475) );
  XNOR2_X1 U567 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U568 ( .A(n478), .ZN(n479) );
  AND2_X1 U569 ( .A1(n479), .A2(G210), .ZN(n480) );
  XNOR2_X1 U570 ( .A(n480), .B(KEYINPUT83), .ZN(n481) );
  XNOR2_X1 U571 ( .A(n482), .B(n481), .ZN(n551) );
  INV_X1 U572 ( .A(n551), .ZN(n525) );
  NAND2_X1 U573 ( .A1(G217), .A2(n484), .ZN(n491) );
  XNOR2_X1 U574 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U575 ( .A(n487), .B(KEYINPUT103), .Z(n489) );
  XNOR2_X1 U576 ( .A(G116), .B(G122), .ZN(n488) );
  XNOR2_X1 U577 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U578 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U579 ( .A(n483), .B(n492), .ZN(n621) );
  INV_X1 U580 ( .A(G902), .ZN(n506) );
  NAND2_X1 U581 ( .A1(n621), .A2(n506), .ZN(n493) );
  INV_X1 U582 ( .A(G478), .ZN(n620) );
  XNOR2_X1 U583 ( .A(n493), .B(n620), .ZN(n550) );
  XOR2_X1 U584 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n496) );
  NAND2_X1 U585 ( .A1(G214), .A2(n494), .ZN(n495) );
  XNOR2_X1 U586 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U587 ( .A(KEYINPUT11), .B(n497), .ZN(n499) );
  XNOR2_X1 U588 ( .A(n499), .B(n498), .ZN(n505) );
  XNOR2_X1 U589 ( .A(G113), .B(G143), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n501), .B(n500), .ZN(n503) );
  XNOR2_X1 U591 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U592 ( .A(n505), .B(n504), .ZN(n641) );
  NAND2_X1 U593 ( .A1(n641), .A2(n506), .ZN(n508) );
  XOR2_X1 U594 ( .A(KEYINPUT13), .B(G475), .Z(n507) );
  XNOR2_X1 U595 ( .A(n508), .B(n507), .ZN(n535) );
  INV_X1 U596 ( .A(KEYINPUT109), .ZN(n509) );
  NAND2_X1 U597 ( .A1(n689), .A2(n688), .ZN(n695) );
  INV_X1 U598 ( .A(n535), .ZN(n549) );
  NAND2_X1 U599 ( .A1(n550), .A2(n549), .ZN(n692) );
  XOR2_X1 U600 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n511) );
  XNOR2_X1 U601 ( .A(n512), .B(n511), .ZN(n725) );
  NAND2_X1 U602 ( .A1(n513), .A2(n570), .ZN(n514) );
  OR2_X1 U603 ( .A1(n575), .A2(n514), .ZN(n522) );
  OR2_X1 U604 ( .A1(n521), .A2(n522), .ZN(n516) );
  INV_X1 U605 ( .A(KEYINPUT28), .ZN(n515) );
  XNOR2_X1 U606 ( .A(n516), .B(n515), .ZN(n518) );
  XNOR2_X1 U607 ( .A(n529), .B(KEYINPUT108), .ZN(n517) );
  AND2_X1 U608 ( .A1(n725), .A2(n673), .ZN(n520) );
  INV_X1 U609 ( .A(KEYINPUT42), .ZN(n519) );
  XNOR2_X1 U610 ( .A(n521), .B(KEYINPUT6), .ZN(n578) );
  INV_X1 U611 ( .A(n522), .ZN(n523) );
  INV_X1 U612 ( .A(n680), .ZN(n674) );
  AND2_X1 U613 ( .A1(n525), .A2(n688), .ZN(n526) );
  NAND2_X1 U614 ( .A1(n674), .A2(n526), .ZN(n527) );
  NOR2_X1 U615 ( .A1(n553), .A2(n527), .ZN(n528) );
  XNOR2_X1 U616 ( .A(n528), .B(KEYINPUT36), .ZN(n530) );
  XNOR2_X2 U617 ( .A(n529), .B(KEYINPUT1), .ZN(n599) );
  NAND2_X1 U618 ( .A1(n530), .A2(n599), .ZN(n531) );
  INV_X1 U619 ( .A(KEYINPUT19), .ZN(n532) );
  INV_X1 U620 ( .A(n669), .ZN(n675) );
  AND2_X1 U621 ( .A1(n675), .A2(KEYINPUT76), .ZN(n533) );
  NAND2_X1 U622 ( .A1(n673), .A2(n533), .ZN(n534) );
  INV_X1 U623 ( .A(KEYINPUT85), .ZN(n543) );
  NAND2_X1 U624 ( .A1(n534), .A2(n543), .ZN(n536) );
  OR2_X1 U625 ( .A1(n550), .A2(n535), .ZN(n682) );
  NAND2_X1 U626 ( .A1(n680), .A2(n682), .ZN(n693) );
  NAND2_X1 U627 ( .A1(n536), .A2(n693), .ZN(n537) );
  NAND2_X1 U628 ( .A1(n537), .A2(KEYINPUT47), .ZN(n547) );
  NAND2_X1 U629 ( .A1(n673), .A2(n675), .ZN(n539) );
  OR2_X1 U630 ( .A1(KEYINPUT47), .A2(n543), .ZN(n538) );
  NAND2_X1 U631 ( .A1(n539), .A2(n538), .ZN(n545) );
  XNOR2_X1 U632 ( .A(KEYINPUT76), .B(n693), .ZN(n541) );
  INV_X1 U633 ( .A(KEYINPUT47), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U635 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U637 ( .A1(n550), .A2(n549), .ZN(n589) );
  NOR2_X1 U638 ( .A1(n589), .A2(n558), .ZN(n552) );
  NAND2_X1 U639 ( .A1(n353), .A2(n552), .ZN(n637) );
  NOR2_X1 U640 ( .A1(n680), .A2(n553), .ZN(n554) );
  NAND2_X1 U641 ( .A1(n554), .A2(n688), .ZN(n555) );
  XNOR2_X1 U642 ( .A(KEYINPUT107), .B(n555), .ZN(n556) );
  INV_X1 U643 ( .A(n599), .ZN(n701) );
  NAND2_X1 U644 ( .A1(n556), .A2(n701), .ZN(n557) );
  XNOR2_X1 U645 ( .A(n557), .B(KEYINPUT43), .ZN(n559) );
  NAND2_X1 U646 ( .A1(n559), .A2(n558), .ZN(n629) );
  OR2_X1 U647 ( .A1(n560), .A2(n682), .ZN(n638) );
  XNOR2_X1 U648 ( .A(n749), .B(KEYINPUT78), .ZN(n615) );
  NOR2_X1 U649 ( .A1(G898), .A2(n561), .ZN(n562) );
  XOR2_X1 U650 ( .A(KEYINPUT93), .B(n562), .Z(n565) );
  INV_X1 U651 ( .A(n563), .ZN(n564) );
  NOR2_X1 U652 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U653 ( .A(n566), .B(KEYINPUT94), .ZN(n567) );
  INV_X1 U654 ( .A(n570), .ZN(n705) );
  OR2_X1 U655 ( .A1(n692), .A2(n705), .ZN(n571) );
  NOR2_X1 U656 ( .A1(n605), .A2(n571), .ZN(n573) );
  XNOR2_X1 U657 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n572) );
  INV_X1 U658 ( .A(KEYINPUT104), .ZN(n574) );
  XNOR2_X1 U659 ( .A(n594), .B(n574), .ZN(n577) );
  INV_X1 U660 ( .A(n575), .ZN(n706) );
  AND2_X1 U661 ( .A1(n704), .A2(n706), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n577), .A2(n576), .ZN(n627) );
  NAND2_X1 U663 ( .A1(n599), .A2(n706), .ZN(n579) );
  XNOR2_X1 U664 ( .A(KEYINPUT81), .B(KEYINPUT32), .ZN(n581) );
  INV_X1 U665 ( .A(KEYINPUT64), .ZN(n580) );
  XNOR2_X1 U666 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U667 ( .A(n583), .B(n582), .ZN(n626) );
  NAND2_X1 U668 ( .A1(n584), .A2(n578), .ZN(n586) );
  XOR2_X1 U669 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n585) );
  NOR2_X1 U670 ( .A1(n724), .A2(n605), .ZN(n588) );
  INV_X1 U671 ( .A(KEYINPUT34), .ZN(n587) );
  XNOR2_X1 U672 ( .A(n588), .B(n587), .ZN(n590) );
  INV_X1 U673 ( .A(KEYINPUT35), .ZN(n591) );
  INV_X1 U674 ( .A(n594), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n578), .A2(n706), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n625) );
  INV_X1 U677 ( .A(n597), .ZN(n700) );
  NOR2_X1 U678 ( .A1(n704), .A2(n700), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n712) );
  OR2_X1 U680 ( .A1(n605), .A2(n712), .ZN(n601) );
  XOR2_X1 U681 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n600) );
  XNOR2_X1 U682 ( .A(n601), .B(n600), .ZN(n683) );
  INV_X1 U683 ( .A(n602), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n603), .A2(n704), .ZN(n604) );
  OR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n607) );
  INV_X1 U686 ( .A(KEYINPUT99), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n607), .B(n606), .ZN(n665) );
  NAND2_X1 U688 ( .A1(n683), .A2(n665), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n608), .A2(n693), .ZN(n609) );
  AND2_X1 U690 ( .A1(n625), .A2(n609), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n612), .A2(n405), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n734), .A2(n749), .ZN(n685) );
  NAND2_X1 U694 ( .A1(n685), .A2(KEYINPUT2), .ZN(n616) );
  INV_X1 U695 ( .A(G952), .ZN(n623) );
  AND2_X1 U696 ( .A1(n623), .A2(G953), .ZN(n661) );
  XNOR2_X1 U697 ( .A(n625), .B(G101), .ZN(G3) );
  XNOR2_X1 U698 ( .A(n626), .B(G119), .ZN(G21) );
  XNOR2_X1 U699 ( .A(n627), .B(G110), .ZN(G12) );
  XOR2_X1 U700 ( .A(G140), .B(KEYINPUT115), .Z(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(G42) );
  XOR2_X1 U702 ( .A(KEYINPUT62), .B(n631), .Z(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n634), .A2(n661), .ZN(n636) );
  XOR2_X1 U705 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n635) );
  XNOR2_X1 U706 ( .A(n636), .B(n635), .ZN(G57) );
  XNOR2_X1 U707 ( .A(n637), .B(G143), .ZN(G45) );
  XNOR2_X1 U708 ( .A(n638), .B(G134), .ZN(G36) );
  XNOR2_X1 U709 ( .A(n639), .B(G131), .ZN(G33) );
  NAND2_X1 U710 ( .A1(n351), .A2(G475), .ZN(n643) );
  XOR2_X1 U711 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n640) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(n644) );
  NOR2_X2 U713 ( .A1(n644), .A2(n661), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n645), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U715 ( .A1(n653), .A2(G210), .ZN(n649) );
  XOR2_X1 U716 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X2 U719 ( .A1(n650), .A2(n661), .ZN(n652) );
  XNOR2_X1 U720 ( .A(KEYINPUT88), .B(KEYINPUT56), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(G51) );
  NAND2_X1 U722 ( .A1(n352), .A2(G217), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n656), .A2(n661), .ZN(G66) );
  NAND2_X1 U725 ( .A1(n352), .A2(G469), .ZN(n660) );
  XOR2_X1 U726 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n657) );
  XNOR2_X1 U727 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n660), .B(n659), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(G54) );
  NOR2_X1 U730 ( .A1(n680), .A2(n665), .ZN(n663) );
  XOR2_X1 U731 ( .A(KEYINPUT112), .B(n663), .Z(n664) );
  XNOR2_X1 U732 ( .A(G104), .B(n664), .ZN(G6) );
  NOR2_X1 U733 ( .A1(n682), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U736 ( .A(G107), .B(n668), .ZN(G9) );
  XOR2_X1 U737 ( .A(G128), .B(KEYINPUT29), .Z(n672) );
  NOR2_X1 U738 ( .A1(n669), .A2(n682), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n673), .A2(n670), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n672), .B(n671), .ZN(G30) );
  INV_X1 U741 ( .A(n673), .ZN(n677) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n679) );
  XNOR2_X1 U744 ( .A(G146), .B(KEYINPUT113), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n679), .B(n678), .ZN(G48) );
  NOR2_X1 U746 ( .A1(n683), .A2(n680), .ZN(n681) );
  XOR2_X1 U747 ( .A(G113), .B(n681), .Z(G15) );
  NOR2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U749 ( .A(G116), .B(n684), .Z(G18) );
  NAND2_X1 U750 ( .A1(n685), .A2(KEYINPUT84), .ZN(n687) );
  XOR2_X1 U751 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n686) );
  XNOR2_X1 U752 ( .A(n687), .B(n686), .ZN(n730) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U754 ( .A(n690), .B(KEYINPUT118), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U756 ( .A(n693), .ZN(n694) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U759 ( .A1(n724), .A2(n698), .ZN(n699) );
  XNOR2_X1 U760 ( .A(n699), .B(KEYINPUT119), .ZN(n718) );
  NAND2_X1 U761 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U762 ( .A(n702), .B(KEYINPUT116), .ZN(n703) );
  XNOR2_X1 U763 ( .A(KEYINPUT50), .B(n703), .ZN(n711) );
  INV_X1 U764 ( .A(n704), .ZN(n709) );
  NAND2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U766 ( .A(n707), .B(KEYINPUT49), .ZN(n708) );
  NOR2_X1 U767 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U768 ( .A1(n711), .A2(n710), .ZN(n713) );
  AND2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U770 ( .A(n714), .B(KEYINPUT51), .Z(n715) );
  XNOR2_X1 U771 ( .A(KEYINPUT117), .B(n715), .ZN(n716) );
  NAND2_X1 U772 ( .A1(n716), .A2(n725), .ZN(n717) );
  NAND2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n720) );
  XOR2_X1 U774 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(n722) );
  NOR2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(KEYINPUT121), .ZN(n728) );
  INV_X1 U778 ( .A(n724), .ZN(n726) );
  NAND2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U782 ( .A(n731), .B(KEYINPUT122), .ZN(n732) );
  XNOR2_X1 U783 ( .A(KEYINPUT53), .B(n733), .ZN(G75) );
  NAND2_X1 U784 ( .A1(n734), .A2(n750), .ZN(n739) );
  NAND2_X1 U785 ( .A1(G224), .A2(G953), .ZN(n735) );
  XNOR2_X1 U786 ( .A(n735), .B(KEYINPUT61), .ZN(n736) );
  XNOR2_X1 U787 ( .A(KEYINPUT126), .B(n736), .ZN(n737) );
  NAND2_X1 U788 ( .A1(n737), .A2(G898), .ZN(n738) );
  NAND2_X1 U789 ( .A1(n739), .A2(n738), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n740), .B(G101), .ZN(n742) );
  NOR2_X1 U791 ( .A1(G898), .A2(n750), .ZN(n741) );
  NOR2_X1 U792 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n745), .B(n498), .ZN(n748) );
  XOR2_X1 U795 ( .A(G227), .B(n748), .Z(n746) );
  NAND2_X1 U796 ( .A1(G900), .A2(n746), .ZN(n747) );
  NAND2_X1 U797 ( .A1(n747), .A2(G953), .ZN(n753) );
  XNOR2_X1 U798 ( .A(n749), .B(n748), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(G72) );
  XNOR2_X1 U801 ( .A(n754), .B(KEYINPUT37), .ZN(n755) );
  XNOR2_X1 U802 ( .A(n755), .B(KEYINPUT114), .ZN(n756) );
  XNOR2_X1 U803 ( .A(G125), .B(n756), .ZN(G27) );
  XNOR2_X1 U804 ( .A(n757), .B(G137), .ZN(G39) );
endmodule

