//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(KEYINPUT31), .ZN(new_n187));
  INV_X1    g001(.A(G113), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT2), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G113), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n189), .B(new_n191), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(new_n191), .ZN(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT30), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(G131), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n202), .B2(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XOR2_X1   g025(.A(KEYINPUT65), .B(G131), .Z(new_n212));
  OAI21_X1  g026(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G128), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n217), .B(new_n219), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT65), .B(G131), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n226), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT66), .A3(new_n206), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n215), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n211), .A2(G131), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n227), .ZN(new_n231));
  XNOR2_X1  g045(.A(G143), .B(G146), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT0), .B(G128), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n220), .A2(KEYINPUT64), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n201), .B1(new_n229), .B2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n227), .A2(new_n222), .A3(new_n224), .A4(new_n206), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n238), .A2(new_n201), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n200), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n243));
  INV_X1    g057(.A(G237), .ZN(new_n244));
  INV_X1    g058(.A(G953), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n244), .A2(new_n245), .A3(G210), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n243), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G101), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n200), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n229), .A2(new_n251), .A3(new_n238), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n242), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n253), .B1(new_n250), .B2(new_n252), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n187), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n256), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n258), .A2(KEYINPUT31), .A3(new_n242), .A4(new_n254), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n229), .A2(new_n251), .A3(new_n238), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n251), .B1(new_n238), .B2(new_n240), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT28), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n261), .B2(KEYINPUT28), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n252), .A2(KEYINPUT69), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n249), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT32), .ZN(new_n271));
  NOR2_X1   g085(.A1(G472), .A2(G902), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n257), .A2(new_n259), .B1(new_n268), .B2(new_n249), .ZN(new_n274));
  INV_X1    g088(.A(new_n272), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT32), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n238), .A2(new_n201), .A3(new_n240), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n222), .A2(new_n224), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n214), .B2(new_n213), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n234), .A2(new_n237), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n281), .A2(new_n228), .B1(new_n282), .B2(new_n231), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n279), .B1(new_n283), .B2(new_n201), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n261), .B1(new_n284), .B2(new_n200), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n278), .B1(new_n285), .B2(new_n250), .ZN(new_n286));
  AND4_X1   g100(.A1(new_n263), .A2(new_n265), .A3(new_n267), .A4(new_n250), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT70), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n242), .A2(new_n252), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT29), .B1(new_n289), .B2(new_n249), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n290), .B(new_n291), .C1(new_n268), .C2(new_n249), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n251), .B1(new_n229), .B2(new_n238), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT28), .B1(new_n261), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n249), .A2(new_n278), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(new_n265), .A3(new_n267), .A4(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(new_n292), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G472), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n277), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT76), .B(KEYINPUT25), .ZN(new_n303));
  INV_X1    g117(.A(G110), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT24), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G110), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n194), .A2(G128), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n223), .A2(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT71), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n194), .B2(G128), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n311), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G110), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT16), .ZN(new_n326));
  OR3_X1    g140(.A1(new_n324), .A2(KEYINPUT16), .A3(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G146), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G146), .B1(new_n326), .B2(new_n327), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n316), .B(new_n321), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n245), .A2(G221), .A3(G234), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G137), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n333), .B2(new_n335), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n324), .A2(G140), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n322), .A2(G125), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT74), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n216), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n314), .B1(new_n310), .B2(new_n315), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT72), .B(G110), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n320), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n344), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n328), .A2(KEYINPUT73), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n326), .A2(new_n327), .A3(new_n350), .A4(G146), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n331), .B(new_n338), .C1(new_n348), .C2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT71), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT71), .B1(new_n305), .B2(new_n307), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n313), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n346), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n358), .A2(new_n311), .A3(new_n319), .A4(new_n318), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n360), .A2(new_n349), .A3(new_n351), .A4(new_n344), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n338), .B1(new_n361), .B2(new_n331), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n297), .B(new_n303), .C1(new_n354), .C2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G217), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(G234), .B2(new_n297), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(KEYINPUT76), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n331), .B1(new_n348), .B2(new_n352), .ZN(new_n370));
  INV_X1    g184(.A(new_n338), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n353), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n373), .B2(new_n297), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n302), .B1(new_n366), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n297), .B1(new_n354), .B2(new_n362), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n368), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(KEYINPUT77), .A3(new_n363), .A4(new_n365), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n365), .A2(G902), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n301), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT9), .B(G234), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n384), .A2(new_n364), .A3(G953), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n192), .A2(G122), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT90), .B(G122), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(new_n192), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G107), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n390), .B(new_n386), .C1(new_n387), .C2(new_n192), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n218), .A2(G128), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n223), .A2(G143), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(new_n202), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n218), .A2(KEYINPUT13), .A3(G128), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT91), .B1(new_n399), .B2(G134), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n399), .A2(KEYINPUT91), .A3(G134), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n392), .B(new_n395), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n192), .A3(G122), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT92), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n387), .B2(new_n192), .ZN(new_n407));
  OAI21_X1  g221(.A(G107), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n393), .A2(new_n394), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G134), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n395), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n391), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n385), .B1(new_n402), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n402), .A2(new_n412), .A3(new_n385), .ZN(new_n415));
  AOI21_X1  g229(.A(G902), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G478), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT15), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n416), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n326), .A2(new_n327), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n216), .ZN(new_n421));
  NOR2_X1   g235(.A1(G237), .A2(G953), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n422), .A2(G143), .A3(G214), .ZN(new_n423));
  AOI21_X1  g237(.A(G143), .B1(new_n422), .B2(G214), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n212), .B(KEYINPUT17), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT89), .A4(new_n328), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n244), .A2(new_n245), .A3(G214), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n218), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(G143), .A3(G214), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n212), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT17), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n226), .A3(new_n429), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n421), .A2(new_n425), .A3(new_n328), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT74), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT74), .B1(new_n323), .B2(new_n325), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(G146), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n323), .A2(new_n325), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G146), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT86), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n344), .A2(new_n446), .A3(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(KEYINPUT18), .A2(G131), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n430), .A2(KEYINPUT85), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n430), .A2(KEYINPUT85), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n430), .B2(KEYINPUT85), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n435), .A2(new_n438), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  INV_X1    g269(.A(G104), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n454), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n297), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G475), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT19), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n342), .A2(new_n462), .A3(new_n343), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n442), .A2(KEYINPUT19), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n216), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n349), .A2(new_n351), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n431), .A2(new_n433), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n463), .A2(new_n469), .A3(new_n216), .A4(new_n464), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n452), .A2(new_n451), .ZN(new_n472));
  INV_X1    g286(.A(new_n450), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n344), .A2(new_n446), .A3(new_n443), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n446), .B1(new_n344), .B2(new_n443), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n457), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n477), .A2(KEYINPUT88), .B1(new_n454), .B2(new_n457), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n476), .ZN(new_n479));
  INV_X1    g293(.A(new_n457), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n461), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n485), .ZN(new_n487));
  AOI211_X1 g301(.A(KEYINPUT20), .B(new_n487), .C1(new_n478), .C2(new_n483), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n419), .B(new_n460), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n245), .A2(G952), .ZN(new_n490));
  NAND2_X1  g304(.A1(G234), .A2(G237), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n491), .A2(G902), .A3(G953), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT3), .B1(new_n456), .B2(G107), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT3), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n390), .A3(G104), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n456), .A2(G107), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(G101), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n501), .A2(G101), .ZN(new_n504));
  INV_X1    g318(.A(G101), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n497), .A2(new_n499), .A3(new_n505), .A4(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n200), .B(new_n503), .C1(new_n504), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT79), .ZN(new_n509));
  XNOR2_X1  g323(.A(G104), .B(G107), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n505), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n390), .A2(G104), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n500), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT79), .A3(G101), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT5), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n188), .B1(new_n193), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n194), .A2(G116), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n192), .A2(G119), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT5), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n517), .A2(new_n520), .B1(new_n198), .B2(new_n197), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n521), .A3(new_n506), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n508), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(G110), .B(G122), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n508), .A2(new_n524), .A3(new_n522), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(KEYINPUT6), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n234), .A2(new_n237), .A3(G125), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(G125), .B2(new_n280), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n245), .A2(G224), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT81), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n530), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT6), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n523), .A2(new_n534), .A3(new_n525), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n528), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT83), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n511), .A2(new_n514), .B1(new_n538), .B2(new_n505), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n539), .B2(new_n521), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT82), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n542), .A3(new_n521), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT79), .B1(new_n513), .B2(G101), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n509), .B(new_n505), .C1(new_n512), .C2(new_n500), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n506), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n521), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT83), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n540), .A2(new_n541), .A3(new_n543), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n524), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n530), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n529), .B(new_n552), .C1(G125), .C2(new_n280), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n527), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n536), .A2(new_n557), .A3(new_n297), .ZN(new_n558));
  OAI21_X1  g372(.A(G210), .B1(G237), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(G902), .B1(new_n551), .B2(new_n556), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n559), .A3(new_n536), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(KEYINPUT84), .A3(new_n563), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n563), .A2(KEYINPUT84), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G214), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G221), .B1(new_n384), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n546), .A2(new_n280), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n515), .A2(new_n506), .B1(new_n224), .B2(new_n222), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n231), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT12), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n546), .B2(new_n280), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n501), .A2(G101), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(KEYINPUT4), .A3(new_n506), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n282), .A2(new_n579), .A3(new_n503), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n225), .A2(KEYINPUT10), .A3(new_n506), .A4(new_n515), .ZN(new_n581));
  INV_X1    g395(.A(new_n231), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n577), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n584), .B(new_n231), .C1(new_n572), .C2(new_n573), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(G110), .B(G140), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT78), .ZN(new_n588));
  INV_X1    g402(.A(G227), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(G953), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n588), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n231), .ZN(new_n594));
  INV_X1    g408(.A(new_n591), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n583), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n592), .A2(G469), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G469), .A2(G902), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n594), .A2(new_n583), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n591), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n575), .A2(new_n595), .A3(new_n583), .A4(new_n585), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(KEYINPUT80), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G469), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n600), .A2(new_n605), .A3(new_n591), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n603), .A2(new_n604), .A3(new_n297), .A4(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n571), .B1(new_n599), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n496), .A2(new_n569), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n383), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT93), .B(G101), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G3));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n402), .B2(new_n412), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n415), .A3(new_n414), .ZN(new_n617));
  INV_X1    g431(.A(new_n415), .ZN(new_n618));
  OAI22_X1  g432(.A1(new_n618), .A2(new_n413), .B1(new_n614), .B2(new_n615), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G478), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n417), .A2(new_n297), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n297), .B1(new_n618), .B2(new_n413), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(G478), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n479), .A2(KEYINPUT88), .A3(new_n480), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n435), .A2(new_n438), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n457), .A3(new_n476), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n477), .A2(KEYINPUT88), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n485), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT20), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n484), .A2(new_n461), .A3(new_n485), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n627), .B1(new_n636), .B2(new_n460), .ZN(new_n637));
  INV_X1    g451(.A(new_n495), .ZN(new_n638));
  INV_X1    g452(.A(new_n563), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n559), .B1(new_n562), .B2(new_n536), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n567), .B(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT95), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(G475), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n458), .B2(new_n297), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n634), .B2(new_n635), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n646), .A2(new_n641), .A3(new_n647), .A4(new_n627), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n607), .A2(new_n598), .A3(new_n597), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n650), .A2(new_n382), .A3(new_n570), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n274), .A2(new_n275), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n270), .A2(new_n297), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n652), .B1(new_n653), .B2(G472), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT34), .B(G104), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  XNOR2_X1  g472(.A(new_n624), .B(new_n418), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n659), .B(new_n460), .C1(new_n486), .C2(new_n488), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n641), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n651), .A2(new_n661), .A3(new_n654), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NOR2_X1   g478(.A1(new_n338), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n370), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n379), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n375), .A2(new_n378), .A3(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n650), .A2(new_n570), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n496), .A3(new_n654), .A4(new_n569), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  AOI21_X1  g486(.A(new_n568), .B1(new_n561), .B2(new_n563), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n570), .A2(new_n650), .A3(new_n673), .A4(new_n668), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n301), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n492), .B1(new_n493), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n636), .A2(new_n659), .A3(new_n460), .A4(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XNOR2_X1  g496(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n566), .B(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n668), .ZN(new_n685));
  INV_X1    g499(.A(G472), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n258), .A2(new_n242), .A3(new_n254), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n249), .B1(new_n261), .B2(new_n293), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n686), .B1(new_n689), .B2(new_n297), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n277), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n646), .A2(new_n568), .A3(new_n419), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n684), .A2(new_n685), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n677), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n608), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT40), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n218), .ZN(G45));
  NOR3_X1   g513(.A1(new_n646), .A2(new_n627), .A3(new_n677), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n675), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  AOI21_X1  g516(.A(new_n381), .B1(new_n277), .B2(new_n300), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n603), .A2(new_n297), .A3(new_n606), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n705), .A2(new_n570), .A3(new_n607), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n703), .B(new_n706), .C1(new_n643), .C2(new_n648), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND3_X1  g523(.A1(new_n703), .A2(new_n661), .A3(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  AND4_X1   g525(.A1(new_n570), .A2(new_n705), .A3(new_n607), .A4(new_n673), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n301), .A2(new_n496), .A3(new_n668), .A4(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT97), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n194), .ZN(G21));
  OAI21_X1  g530(.A(new_n460), .B1(new_n486), .B2(new_n488), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n639), .A2(new_n640), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n717), .A2(new_n567), .A3(new_n719), .A4(new_n659), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n265), .A2(new_n294), .A3(new_n267), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n260), .B1(new_n250), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n272), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT98), .B(G472), .Z(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n274), .B2(G902), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n724), .A2(new_n382), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n721), .A2(new_n638), .A3(new_n727), .A4(new_n706), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  AND3_X1   g543(.A1(new_n724), .A2(new_n668), .A3(new_n726), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n700), .A3(new_n712), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NAND2_X1  g546(.A1(new_n592), .A2(KEYINPUT99), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT99), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n586), .A2(new_n734), .A3(new_n591), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(G469), .A3(new_n596), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n607), .A2(new_n736), .A3(new_n598), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n566), .A3(new_n567), .A4(new_n570), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n703), .A2(new_n739), .A3(new_n700), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n703), .A2(new_n739), .A3(KEYINPUT42), .A4(new_n700), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NAND3_X1  g559(.A1(new_n703), .A2(new_n739), .A3(new_n680), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  OAI21_X1  g561(.A(KEYINPUT102), .B1(new_n654), .B2(new_n685), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n625), .B1(G478), .B2(new_n620), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n749), .B(new_n460), .C1(new_n486), .C2(new_n488), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT101), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n751), .B(new_n460), .C1(new_n486), .C2(new_n488), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n646), .B(new_n749), .C1(new_n751), .C2(KEYINPUT43), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(G472), .B1(new_n274), .B2(G902), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n270), .A2(new_n272), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n685), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT102), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n748), .A2(new_n756), .A3(KEYINPUT44), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n566), .A2(new_n567), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n695), .ZN(new_n766));
  INV_X1    g580(.A(new_n607), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n592), .A2(new_n596), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n604), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n733), .A2(KEYINPUT45), .A3(new_n596), .A4(new_n735), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT100), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n772), .B1(new_n770), .B2(new_n771), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n598), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n767), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(KEYINPUT46), .B(new_n598), .C1(new_n773), .C2(new_n774), .ZN(new_n778));
  AOI211_X1 g592(.A(new_n571), .B(new_n766), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n754), .A2(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n780));
  AOI211_X1 g594(.A(KEYINPUT103), .B(KEYINPUT44), .C1(new_n780), .C2(new_n748), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT103), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n748), .A2(new_n756), .A3(new_n761), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n765), .B(new_n779), .C1(new_n781), .C2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  AOI22_X1  g601(.A1(new_n276), .A2(new_n273), .B1(new_n299), .B2(G472), .ZN(new_n788));
  AND4_X1   g602(.A1(new_n788), .A2(new_n764), .A3(new_n700), .A4(new_n381), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n790), .B(new_n571), .C1(new_n777), .C2(new_n778), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n775), .A2(new_n776), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n607), .A3(new_n778), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT47), .B1(new_n793), .B2(new_n570), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n789), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  AND2_X1   g610(.A1(new_n705), .A2(new_n607), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT49), .ZN(new_n798));
  INV_X1    g612(.A(new_n684), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n690), .B1(new_n273), .B2(new_n276), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n750), .A2(new_n381), .A3(new_n568), .A4(new_n571), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n490), .ZN(new_n803));
  INV_X1    g617(.A(new_n706), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n763), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n382), .A2(new_n805), .A3(new_n492), .A4(new_n800), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n803), .B1(new_n806), .B2(new_n637), .ZN(new_n807));
  INV_X1    g621(.A(new_n492), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n754), .B2(new_n755), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n712), .A3(new_n727), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(KEYINPUT112), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT112), .B1(new_n807), .B2(new_n810), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n805), .A3(new_n703), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT48), .Z(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n806), .A2(new_n646), .A3(new_n627), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n809), .A2(new_n805), .A3(new_n730), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n809), .A2(new_n727), .ZN(new_n819));
  OR4_X1    g633(.A1(new_n567), .A2(new_n819), .A3(new_n684), .A4(new_n804), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n820), .A2(new_n822), .ZN(new_n824));
  OAI211_X1 g638(.A(KEYINPUT51), .B(new_n818), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n791), .A2(new_n794), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n797), .A2(new_n571), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n763), .B(new_n819), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n811), .B(new_n815), .C1(new_n825), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n823), .A2(new_n824), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n818), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n375), .A2(new_n378), .A3(new_n667), .A4(new_n678), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT104), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n737), .A2(new_n570), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT105), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT104), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n838), .B(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n840), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT105), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n800), .A2(new_n720), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n841), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n301), .B(new_n674), .C1(new_n680), .C2(new_n700), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n731), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n837), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n841), .A2(new_n846), .A3(new_n847), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n731), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n707), .A2(new_n710), .A3(new_n728), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n715), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n739), .A2(new_n700), .A3(new_n730), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n489), .A2(new_n677), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n301), .A2(new_n669), .A3(new_n764), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n746), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n660), .B1(new_n646), .B2(new_n627), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n567), .A2(new_n564), .A3(new_n565), .A4(new_n638), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n651), .A3(new_n654), .A4(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n863), .B(new_n670), .C1(new_n383), .C2(new_n609), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n854), .A2(new_n856), .A3(new_n744), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n851), .A2(new_n853), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n713), .B(KEYINPUT97), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n707), .A2(new_n710), .A3(new_n728), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n870), .A3(new_n744), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n867), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n868), .A2(KEYINPUT106), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT106), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n866), .A2(new_n875), .A3(new_n867), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(KEYINPUT54), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT107), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n866), .A2(KEYINPUT107), .A3(new_n867), .ZN(new_n880));
  XOR2_X1   g694(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n881));
  OAI21_X1  g695(.A(KEYINPUT108), .B1(new_n715), .B2(new_n855), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT108), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n870), .A2(new_n871), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n744), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n854), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n879), .A2(new_n880), .A3(new_n881), .A4(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n836), .A2(new_n877), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(G952), .A2(G953), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT113), .Z(new_n891));
  OAI21_X1  g705(.A(new_n802), .B1(new_n889), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n245), .A2(G952), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT114), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n879), .A2(new_n880), .A3(new_n887), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(G210), .A3(G902), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n528), .A2(new_n535), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n533), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n902), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n895), .B1(new_n903), .B2(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n887), .A2(new_n881), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n907), .A2(new_n879), .A3(new_n908), .A4(new_n880), .ZN(new_n909));
  INV_X1    g723(.A(new_n881), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n896), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n598), .B(KEYINPUT57), .Z(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n603), .A3(new_n606), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n773), .A2(new_n774), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n896), .A2(G902), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n893), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND4_X1  g732(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT116), .ZN(new_n920));
  INV_X1    g734(.A(new_n484), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n893), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n919), .B2(new_n921), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(G60));
  XNOR2_X1  g740(.A(new_n622), .B(KEYINPUT59), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n877), .B2(new_n888), .ZN(new_n928));
  INV_X1    g742(.A(new_n620), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n894), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n620), .A2(new_n927), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n912), .B2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT117), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n896), .A2(new_n666), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n896), .A2(KEYINPUT118), .A3(new_n666), .A4(new_n935), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n373), .B1(new_n896), .B2(new_n935), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(new_n895), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n940), .A2(KEYINPUT61), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(G66));
  NOR3_X1   g761(.A1(new_n715), .A2(new_n864), .A3(new_n855), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(G953), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT119), .ZN(new_n950));
  INV_X1    g764(.A(G224), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n494), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n900), .B1(G898), .B2(new_n245), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  NAND2_X1  g769(.A1(new_n463), .A2(new_n464), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n284), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n676), .A2(G953), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n779), .A2(new_n703), .A3(new_n721), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n744), .B2(new_n746), .ZN(new_n961));
  NOR4_X1   g775(.A1(new_n788), .A2(new_n738), .A3(new_n381), .A4(new_n679), .ZN(new_n962));
  AOI211_X1 g776(.A(KEYINPUT124), .B(new_n962), .C1(new_n742), .C2(new_n743), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n795), .B(new_n959), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n850), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n781), .A2(new_n785), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n571), .B1(new_n777), .B2(new_n778), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n967), .A2(new_n695), .A3(new_n764), .A4(new_n762), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n965), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT123), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT123), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n786), .A2(new_n971), .A3(new_n965), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n964), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n958), .B1(new_n973), .B2(G953), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n957), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(KEYINPUT125), .B(new_n958), .C1(new_n973), .C2(G953), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n589), .B2(new_n676), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT122), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n694), .A2(new_n697), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(KEYINPUT62), .A3(new_n965), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n698), .B2(new_n850), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n985), .A2(new_n795), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n696), .A2(new_n763), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n703), .A3(new_n861), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n786), .A2(KEYINPUT120), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT120), .B1(new_n786), .B2(new_n988), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT121), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT121), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n986), .B(new_n993), .C1(new_n989), .C2(new_n990), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n995), .A2(new_n245), .A3(new_n957), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n978), .A2(new_n980), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n980), .B1(new_n978), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n997), .A2(new_n998), .ZN(G72));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n289), .A2(new_n249), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n687), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n874), .A2(new_n876), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n285), .A2(new_n249), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n961), .A2(new_n963), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n795), .A2(new_n959), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n971), .B1(new_n786), .B2(new_n965), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n786), .A2(new_n971), .A3(new_n965), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1010), .B(new_n948), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1007), .B1(new_n1013), .B2(new_n1001), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1006), .B1(new_n1014), .B2(new_n893), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1002), .B1(new_n973), .B2(new_n948), .ZN(new_n1016));
  OAI211_X1 g830(.A(KEYINPUT127), .B(new_n923), .C1(new_n1016), .C2(new_n1007), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1005), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT126), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n992), .A2(new_n948), .A3(new_n994), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n1001), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n285), .A2(new_n249), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1022), .ZN(new_n1024));
  AOI211_X1 g838(.A(KEYINPUT126), .B(new_n1024), .C1(new_n1020), .C2(new_n1001), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1018), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(G57));
endmodule


