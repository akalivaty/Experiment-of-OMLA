//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n592, new_n594, new_n595, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1129, new_n1130,
    new_n1131, new_n1132;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n459), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT66), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n472), .B2(G2105), .ZN(G160));
  NOR2_X1   g048(.A1(new_n460), .A2(new_n461), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n459), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NOR3_X1   g055(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G112), .B2(new_n459), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n476), .A2(new_n478), .A3(new_n482), .ZN(G162));
  NAND2_X1  g058(.A1(G114), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G102), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n469), .A2(new_n494), .A3(G138), .A4(new_n459), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n460), .B2(new_n461), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(new_n497), .C1(new_n460), .C2(new_n461), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n491), .A2(new_n496), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XOR2_X1   g079(.A(KEYINPUT5), .B(G543), .Z(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OR3_X1    g081(.A1(new_n505), .A2(KEYINPUT70), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT70), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n513), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n505), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G50), .B1(G88), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n511), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n516), .A2(G51), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n514), .A2(G89), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n518), .A2(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n532), .B2(new_n515), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n533), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n535), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT71), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n516), .A2(G43), .B1(G81), .B2(new_n518), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G860), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT72), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OR3_X1    g127(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n515), .B2(new_n552), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n553), .A2(new_n554), .B1(G91), .B2(new_n518), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT73), .B(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n505), .B2(new_n557), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(KEYINPUT74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(KEYINPUT74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(G651), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n555), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND2_X1  g138(.A1(new_n518), .A2(G87), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT75), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n525), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n516), .A2(G49), .B1(G651), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G288));
  AOI22_X1  g143(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n535), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n516), .A2(G48), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n518), .A2(G86), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n535), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT76), .Z(new_n576));
  AOI22_X1  g151(.A1(new_n516), .A2(G47), .B1(G85), .B2(new_n518), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G290));
  INV_X1    g153(.A(G868), .ZN(new_n579));
  NOR2_X1   g154(.A1(G301), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n518), .A2(G92), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT10), .Z(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n505), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n516), .A2(G54), .B1(new_n585), .B2(G651), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n580), .B1(new_n587), .B2(new_n579), .ZN(G284));
  AOI21_X1  g163(.A(new_n580), .B1(new_n587), .B2(new_n579), .ZN(G321));
  MUX2_X1   g164(.A(G286), .B(G299), .S(new_n579), .Z(G297));
  MUX2_X1   g165(.A(G286), .B(G299), .S(new_n579), .Z(G280));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n587), .B1(new_n592), .B2(G860), .ZN(G148));
  INV_X1    g168(.A(new_n543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n579), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n587), .A2(new_n592), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n579), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT11), .Z(G282));
  INV_X1    g173(.A(new_n597), .ZN(G323));
  NAND2_X1  g174(.A1(new_n475), .A2(G2104), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT12), .Z(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(KEYINPUT78), .B2(G2100), .ZN(new_n604));
  NAND2_X1  g179(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n603), .A2(KEYINPUT78), .A3(G2100), .ZN(new_n607));
  MUX2_X1   g182(.A(G99), .B(G111), .S(G2105), .Z(new_n608));
  AOI22_X1  g183(.A1(new_n475), .A2(G135), .B1(G2104), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n477), .A2(new_n610), .A3(G123), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(new_n477), .B2(G123), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G2096), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n606), .A2(new_n607), .A3(new_n615), .ZN(G156));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2438), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2427), .B(G2430), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT14), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT80), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n618), .B2(new_n619), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2443), .B(G2446), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT81), .ZN(new_n631));
  INV_X1    g206(.A(G14), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n628), .B2(new_n629), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(G401));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT82), .ZN(new_n637));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT18), .ZN(new_n642));
  INV_X1    g217(.A(new_n638), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n640), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(KEYINPUT17), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n643), .A2(KEYINPUT17), .A3(new_n639), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n639), .B1(new_n643), .B2(KEYINPUT17), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(new_n637), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n642), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(new_n614), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(G227));
  XOR2_X1   g226(.A(G1971), .B(G1976), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n656), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT20), .Z(new_n660));
  AOI211_X1 g235(.A(new_n658), .B(new_n660), .C1(new_n653), .C2(new_n657), .ZN(new_n661));
  XOR2_X1   g236(.A(G1981), .B(G1986), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT83), .ZN(new_n665));
  XOR2_X1   g240(.A(G1991), .B(G1996), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(G229));
  NAND2_X1  g243(.A1(new_n587), .A2(G16), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(G4), .B2(G16), .ZN(new_n670));
  INV_X1    g245(.A(G1348), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  MUX2_X1   g248(.A(G104), .B(G116), .S(G2105), .Z(new_n674));
  AOI22_X1  g249(.A1(new_n477), .A2(G128), .B1(G2104), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G140), .ZN(new_n676));
  INV_X1    g251(.A(new_n475), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G29), .ZN(new_n679));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G26), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G2067), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n672), .A2(new_n673), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(G29), .A2(G35), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G162), .B2(G29), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n686), .B1(G2090), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G20), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT23), .Z(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G299), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G1956), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n691), .A2(G2090), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(KEYINPUT96), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n701));
  NOR2_X1   g276(.A1(G16), .A2(G19), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n594), .B2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1341), .Z(new_n704));
  NAND4_X1  g279(.A1(new_n692), .A2(new_n700), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(KEYINPUT24), .A2(G34), .ZN(new_n706));
  NAND2_X1  g281(.A1(KEYINPUT24), .A2(G34), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G160), .B2(G29), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(G2084), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n693), .A2(G21), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G168), .B2(new_n693), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G1966), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT92), .ZN(new_n715));
  NOR2_X1   g290(.A1(G27), .A2(G29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G164), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G2078), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT31), .B(G11), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT30), .B(G28), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n680), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n693), .A2(G5), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G301), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n722), .B1(new_n680), .B2(new_n613), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G1966), .B2(new_n713), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n469), .A2(G127), .ZN(new_n729));
  AND2_X1   g304(.A1(G115), .A2(G2104), .ZN(new_n730));
  OAI21_X1  g305(.A(G2105), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n475), .A2(G139), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n463), .A2(G103), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n731), .B(new_n732), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G33), .B(new_n737), .S(G29), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2072), .ZN(new_n739));
  NOR4_X1   g314(.A1(new_n719), .A2(new_n726), .A3(new_n728), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n709), .A2(G2084), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT88), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G32), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n475), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n477), .A2(G129), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT89), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT26), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n743), .B1(new_n750), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT91), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n752), .B(new_n754), .ZN(new_n755));
  AND4_X1   g330(.A1(new_n711), .A2(new_n740), .A3(new_n742), .A4(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n705), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G6), .B(G305), .S(G16), .Z(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT32), .B(G1981), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(G166), .A2(G16), .ZN(new_n764));
  OR2_X1    g339(.A1(G16), .A2(G22), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n763), .B1(G1971), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1971), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n693), .A2(G23), .ZN(new_n771));
  INV_X1    g346(.A(G288), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n693), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT33), .B(G1976), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AND3_X1   g350(.A1(new_n768), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT34), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  MUX2_X1   g354(.A(G24), .B(G290), .S(G16), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G1986), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(G1986), .ZN(new_n782));
  INV_X1    g357(.A(G25), .ZN(new_n783));
  OAI21_X1  g358(.A(KEYINPUT84), .B1(new_n783), .B2(G29), .ZN(new_n784));
  OR3_X1    g359(.A1(new_n783), .A2(KEYINPUT84), .A3(G29), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n475), .A2(G131), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n477), .A2(G119), .ZN(new_n787));
  OAI21_X1  g362(.A(KEYINPUT85), .B1(G95), .B2(G2105), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g364(.A1(KEYINPUT85), .A2(G95), .A3(G2105), .ZN(new_n790));
  OAI221_X1 g365(.A(G2104), .B1(G107), .B2(new_n459), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n786), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n784), .B(new_n785), .C1(new_n793), .C2(new_n680), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  XOR2_X1   g370(.A(new_n794), .B(new_n795), .Z(new_n796));
  NOR2_X1   g371(.A1(new_n782), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n778), .A2(new_n779), .A3(new_n781), .A4(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT36), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(KEYINPUT86), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n760), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(G311));
  XNOR2_X1  g378(.A(new_n802), .B(KEYINPUT97), .ZN(G150));
  NAND2_X1  g379(.A1(new_n516), .A2(G55), .ZN(new_n805));
  INV_X1    g380(.A(new_n518), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT99), .B(G93), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n805), .B1(new_n806), .B2(new_n807), .C1(new_n535), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G860), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT37), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n543), .B(new_n809), .ZN(new_n812));
  INV_X1    g387(.A(new_n587), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n592), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n544), .B1(new_n818), .B2(KEYINPUT39), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n811), .B1(new_n819), .B2(new_n820), .ZN(G145));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n822));
  AND4_X1   g397(.A1(new_n822), .A2(new_n491), .A3(new_n496), .A4(new_n502), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n489), .A2(new_n490), .B1(new_n499), .B2(new_n501), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n824), .B2(new_n496), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(new_n678), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n750), .B(new_n737), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n827), .B(new_n828), .Z(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G106), .B(G118), .S(G2105), .Z(new_n831));
  AOI22_X1  g406(.A1(new_n477), .A2(G130), .B1(G2104), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G142), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n677), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n601), .B(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n792), .B(KEYINPUT101), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n830), .A2(new_n837), .ZN(new_n839));
  XNOR2_X1  g414(.A(G162), .B(G160), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n613), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n837), .A2(KEYINPUT102), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n841), .B1(new_n830), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n830), .B2(new_n843), .ZN(new_n845));
  INV_X1    g420(.A(G37), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n842), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g423(.A1(new_n809), .A2(new_n579), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT106), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n587), .A2(G299), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n587), .A2(G299), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT41), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT104), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n853), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n855), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n812), .B(new_n596), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n857), .A2(new_n862), .ZN(new_n866));
  INV_X1    g441(.A(new_n864), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(KEYINPUT105), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n854), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n772), .B(G290), .ZN(new_n871));
  XOR2_X1   g446(.A(G166), .B(G305), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT42), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n850), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n868), .A2(new_n869), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n877), .A2(KEYINPUT106), .A3(new_n865), .A4(new_n874), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(new_n875), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n849), .B1(new_n880), .B2(new_n579), .ZN(G295));
  OAI21_X1  g456(.A(new_n849), .B1(new_n880), .B2(new_n579), .ZN(G331));
  INV_X1    g457(.A(new_n873), .ZN(new_n883));
  XNOR2_X1  g458(.A(G301), .B(G168), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n812), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n854), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n883), .B(new_n886), .C1(new_n863), .C2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n885), .A2(new_n855), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(new_n854), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n861), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n873), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT107), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n889), .A2(new_n893), .A3(new_n873), .A4(new_n890), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n887), .A2(new_n892), .A3(new_n846), .A4(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n886), .B1(new_n863), .B2(new_n885), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n873), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n899), .A2(KEYINPUT43), .A3(new_n846), .A4(new_n887), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n895), .A2(KEYINPUT43), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n846), .A3(new_n887), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(KEYINPUT43), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(KEYINPUT44), .B2(new_n904), .ZN(G397));
  XNOR2_X1  g480(.A(KEYINPUT108), .B(G1384), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT45), .B1(new_n826), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(KEYINPUT109), .B(G40), .ZN(new_n909));
  AOI211_X1 g484(.A(new_n909), .B(new_n465), .C1(new_n472), .C2(G2105), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n750), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G1996), .ZN(new_n913));
  INV_X1    g488(.A(G1996), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n750), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n678), .B(new_n684), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n793), .A2(new_n795), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n793), .A2(new_n795), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G290), .B(G1986), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G8), .ZN(new_n924));
  NOR2_X1   g499(.A1(G166), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT55), .Z(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT45), .B1(new_n503), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n472), .A2(G2105), .ZN(new_n930));
  INV_X1    g505(.A(new_n465), .ZN(new_n931));
  INV_X1    g506(.A(new_n909), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n500), .B1(new_n469), .B2(new_n497), .ZN(new_n935));
  INV_X1    g510(.A(new_n501), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n486), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT69), .B1(new_n486), .B2(G2104), .ZN(new_n938));
  OAI22_X1  g513(.A1(new_n935), .A2(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n493), .A2(new_n495), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT100), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n824), .A2(new_n822), .A3(new_n496), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT45), .A4(new_n907), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n934), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G2090), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n503), .A2(new_n928), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G1384), .B1(new_n824), .B2(new_n496), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n933), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n947), .A2(new_n769), .B1(new_n948), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n948), .ZN(new_n957));
  INV_X1    g532(.A(new_n934), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n826), .A2(KEYINPUT110), .A3(KEYINPUT45), .A4(new_n907), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n943), .A2(new_n944), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(KEYINPUT111), .B(new_n957), .C1(new_n961), .C2(G1971), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(G8), .B(new_n927), .C1(new_n956), .C2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n926), .B1(new_n955), .B2(new_n924), .ZN(new_n965));
  OAI21_X1  g540(.A(G8), .B1(new_n949), .B2(new_n933), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT112), .Z(new_n967));
  NAND2_X1  g542(.A1(new_n772), .A2(G1976), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G305), .A2(G1981), .ZN(new_n972));
  INV_X1    g547(.A(G1981), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n570), .A2(new_n571), .A3(new_n973), .A4(new_n572), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT113), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n972), .A2(new_n978), .A3(KEYINPUT49), .A4(new_n974), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n977), .A2(new_n979), .B1(new_n976), .B2(new_n975), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n967), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n971), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n967), .A2(new_n968), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(KEYINPUT52), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n964), .A2(new_n965), .A3(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT116), .B(G2084), .Z(new_n986));
  NAND2_X1  g561(.A1(new_n954), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n929), .B2(new_n933), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n952), .A2(KEYINPUT45), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n910), .B(KEYINPUT114), .C1(new_n952), .C2(KEYINPUT45), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1966), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n992), .A2(KEYINPUT115), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT115), .B1(new_n992), .B2(new_n993), .ZN(new_n995));
  OAI211_X1 g570(.A(G168), .B(new_n987), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G8), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT51), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT62), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n987), .B1(new_n994), .B2(new_n995), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(G286), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n998), .B(new_n999), .C1(new_n997), .C2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n947), .B2(G2078), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n954), .A2(G1961), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G2078), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(G301), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1000), .B1(new_n996), .B2(G8), .ZN(new_n1013));
  INV_X1    g588(.A(new_n997), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n1007), .B2(G1966), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n992), .A2(KEYINPUT115), .A3(new_n993), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1016), .A2(new_n1017), .B1(new_n954), .B2(new_n986), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT51), .B1(new_n1018), .B2(G168), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1013), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT125), .B1(new_n1020), .B2(new_n999), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT125), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1002), .A2(new_n997), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1022), .B(KEYINPUT62), .C1(new_n1023), .C2(new_n1013), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1012), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G301), .B(KEYINPUT54), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n472), .B(KEYINPUT124), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G2105), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1029), .A2(G40), .A3(new_n931), .A4(new_n1009), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n908), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n959), .A2(new_n960), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n1027), .B(new_n1006), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1026), .A2(new_n1027), .B1(new_n1033), .B2(new_n1005), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1023), .B2(new_n1013), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT61), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n954), .A2(G1956), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT56), .B(G2072), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n961), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1040), .A2(KEYINPUT119), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(KEYINPUT119), .ZN(new_n1042));
  NOR3_X1   g617(.A1(G299), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(G299), .A2(new_n1042), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n934), .B(new_n1038), .C1(new_n945), .C2(new_n946), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1037), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1036), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n954), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n949), .A2(new_n933), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1052), .A2(new_n671), .B1(new_n684), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(KEYINPUT60), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n684), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT60), .B(new_n1057), .C1(new_n954), .C2(G1348), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1058), .B2(new_n587), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n587), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1056), .A3(new_n587), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT58), .B(G1341), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1053), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n961), .B2(new_n914), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1064), .B1(new_n1067), .B2(new_n543), .ZN(new_n1068));
  AOI211_X1 g643(.A(G1996), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT59), .B(new_n594), .C1(new_n1069), .C2(new_n1066), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1063), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1045), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1036), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1047), .A2(new_n1048), .A3(new_n1045), .A4(new_n1077), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1073), .B(new_n1076), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1049), .A2(KEYINPUT120), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1079), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1073), .B1(new_n1084), .B2(new_n1076), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1051), .B(new_n1072), .C1(new_n1082), .C2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1054), .A2(new_n813), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1049), .B1(new_n1046), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1035), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n985), .B1(new_n1025), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n964), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n981), .A2(new_n969), .A3(new_n772), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n974), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1091), .A2(new_n984), .B1(new_n967), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1018), .A2(new_n924), .A3(G286), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n964), .A2(new_n984), .A3(new_n965), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(KEYINPUT117), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(G8), .B1(new_n956), .B2(new_n963), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n926), .ZN(new_n1100));
  NOR4_X1   g675(.A1(new_n1018), .A2(new_n1097), .A3(new_n924), .A4(G286), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1100), .A2(new_n964), .A3(new_n984), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT117), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT118), .B(new_n1094), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1090), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(new_n1098), .A3(new_n1102), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT118), .B1(new_n1110), .B2(new_n1094), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n923), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(G290), .A2(G1986), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT48), .B1(new_n911), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n911), .A2(KEYINPUT48), .A3(new_n1113), .ZN(new_n1115));
  AOI211_X1 g690(.A(new_n1114), .B(new_n1115), .C1(new_n921), .C2(new_n911), .ZN(new_n1116));
  INV_X1    g691(.A(new_n916), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n911), .B1(new_n912), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n911), .A2(new_n914), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1119), .A2(KEYINPUT46), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(KEYINPUT46), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1123));
  XNOR2_X1  g698(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n917), .A2(new_n920), .B1(G2067), .B2(new_n678), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n1116), .B(new_n1124), .C1(new_n911), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1112), .A2(new_n1126), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g702(.A1(new_n897), .A2(new_n900), .ZN(new_n1129));
  INV_X1    g703(.A(G319), .ZN(new_n1130));
  NOR3_X1   g704(.A1(G229), .A2(new_n1130), .A3(G227), .ZN(new_n1131));
  AND3_X1   g705(.A1(new_n634), .A2(new_n847), .A3(new_n1131), .ZN(new_n1132));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1132), .ZN(G308));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(G225));
endmodule


