//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G469), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n192), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(G104), .A3(new_n196), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n201), .A3(new_n203), .A4(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT4), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n196), .A2(G104), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n204), .A2(G107), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(new_n202), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n201), .B1(new_n210), .B2(new_n200), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n214), .A2(new_n202), .B1(G104), .B2(new_n196), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n205), .B1(new_n197), .B2(new_n198), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n213), .B(G101), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n220), .A2(KEYINPUT64), .A3(G143), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT64), .B1(new_n220), .B2(G143), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT0), .B(G128), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n218), .A2(G146), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT65), .B1(new_n220), .B2(G143), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n218), .A3(G146), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n227), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n217), .A2(new_n226), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT79), .B1(new_n212), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(G101), .B1(new_n215), .B2(new_n216), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n238));
  AOI211_X1 g052(.A(new_n232), .B(new_n227), .C1(new_n228), .C2(new_n230), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n218), .B2(G146), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n220), .A2(KEYINPUT64), .A3(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n224), .B1(new_n243), .B2(new_n219), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT79), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n238), .A2(new_n245), .A3(new_n246), .A4(new_n217), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(G134), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT11), .B1(new_n251), .B2(G137), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(new_n249), .A3(G134), .ZN(new_n254));
  AOI211_X1 g068(.A(G131), .B(new_n250), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n254), .ZN(new_n257));
  INV_X1    g071(.A(new_n250), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G101), .B1(new_n209), .B2(new_n208), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n206), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT1), .B1(new_n218), .B2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G128), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G128), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n223), .A2(new_n265), .B1(new_n231), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT10), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n267), .B(new_n227), .C1(new_n228), .C2(new_n230), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n228), .A2(new_n230), .ZN(new_n273));
  INV_X1    g087(.A(new_n227), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n273), .A2(new_n274), .B1(G128), .B2(new_n264), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n206), .B(new_n261), .C1(new_n272), .C2(new_n275), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n263), .A2(new_n271), .B1(new_n276), .B2(new_n270), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n248), .A2(new_n260), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n260), .B1(new_n248), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n195), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n269), .A2(new_n262), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n257), .A2(new_n258), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G131), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n257), .A2(new_n256), .A3(new_n258), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT12), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n260), .B1(new_n276), .B2(new_n281), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT12), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n195), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n248), .A2(new_n260), .A3(new_n277), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n280), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n191), .B1(new_n296), .B2(new_n189), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n292), .A2(KEYINPUT80), .A3(new_n294), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT80), .B1(new_n292), .B2(new_n294), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n195), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n278), .A2(new_n279), .A3(new_n195), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(G469), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G475), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT87), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(new_n193), .A3(G143), .A4(G214), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n256), .ZN(new_n309));
  NOR2_X1   g123(.A1(G237), .A2(G953), .ZN(new_n310));
  AOI21_X1  g124(.A(G143), .B1(new_n310), .B2(G214), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n307), .A2(new_n193), .A3(G214), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n218), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n314), .A2(KEYINPUT87), .A3(new_n256), .A4(new_n308), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT17), .ZN(new_n316));
  NAND2_X1  g130(.A1(G143), .A2(G214), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n317), .A2(G237), .A3(G953), .ZN(new_n318));
  OAI21_X1  g132(.A(G131), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n312), .A2(new_n315), .A3(new_n316), .A4(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n319), .A2(new_n316), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT16), .ZN(new_n326));
  OR3_X1    g140(.A1(new_n324), .A2(KEYINPUT16), .A3(G140), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n326), .A2(G146), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(G146), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n320), .A2(new_n321), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(KEYINPUT18), .A2(G131), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n311), .A2(new_n318), .A3(KEYINPUT85), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n314), .B2(new_n308), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G214), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n338), .A2(G237), .A3(G953), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n332), .B(new_n308), .C1(new_n339), .C2(G143), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT86), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n314), .A2(new_n342), .A3(new_n332), .A4(new_n308), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n323), .A2(new_n325), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(new_n220), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G113), .B(G122), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(new_n204), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n331), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n312), .A2(new_n315), .A3(new_n319), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT19), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT19), .B1(new_n323), .B2(new_n325), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n220), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT88), .ZN(new_n355));
  INV_X1    g169(.A(new_n328), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(new_n220), .C1(new_n352), .C2(new_n353), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n351), .A2(new_n355), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n349), .B1(new_n359), .B2(new_n347), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n305), .B1(new_n350), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT20), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n363), .B(new_n305), .C1(new_n350), .C2(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT90), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n349), .B1(new_n331), .B2(new_n347), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n350), .A2(new_n367), .A3(KEYINPUT89), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n331), .A2(new_n347), .ZN(new_n369));
  INV_X1    g183(.A(new_n349), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(KEYINPUT89), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n190), .ZN(new_n372));
  OAI21_X1  g186(.A(G475), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n365), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n366), .B1(new_n365), .B2(new_n373), .ZN(new_n375));
  INV_X1    g189(.A(G122), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(G116), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT91), .B(G122), .ZN(new_n379));
  INV_X1    g193(.A(G116), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT14), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G107), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n376), .A2(KEYINPUT91), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G116), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(new_n378), .C1(KEYINPUT14), .C2(new_n196), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n218), .A2(G128), .ZN(new_n390));
  INV_X1    g204(.A(G128), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G143), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT92), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT92), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n390), .B2(new_n392), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n394), .A2(new_n251), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(KEYINPUT92), .ZN(new_n398));
  XNOR2_X1  g212(.A(G128), .B(G143), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n395), .ZN(new_n400));
  AOI21_X1  g214(.A(G134), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n383), .B(new_n389), .C1(new_n397), .C2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n251), .B1(new_n394), .B2(new_n396), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n404), .B(G134), .C1(KEYINPUT13), .C2(new_n390), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n196), .B1(new_n388), .B2(new_n378), .ZN(new_n406));
  AOI211_X1 g220(.A(G107), .B(new_n377), .C1(new_n387), .C2(G116), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n403), .B(new_n405), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G217), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n187), .A2(new_n409), .A3(G953), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n402), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n402), .B2(new_n408), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n190), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT93), .ZN(new_n414));
  INV_X1    g228(.A(G478), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(KEYINPUT15), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(new_n190), .C1(new_n411), .C2(new_n412), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n413), .A2(new_n416), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n193), .A2(G952), .ZN(new_n421));
  INV_X1    g235(.A(G234), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n307), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI211_X1 g238(.A(new_n190), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n419), .A2(new_n420), .A3(new_n428), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n374), .A2(new_n375), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G214), .B1(G237), .B2(G902), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G210), .B1(G237), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(KEYINPUT2), .A2(G113), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT67), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT2), .ZN(new_n438));
  INV_X1    g252(.A(G113), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n436), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G119), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G116), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT69), .B(G119), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(G116), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT68), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n442), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n443), .A2(KEYINPUT69), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G119), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n451), .A3(G116), .ZN(new_n452));
  INV_X1    g266(.A(new_n444), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n441), .ZN(new_n455));
  NOR3_X1   g269(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n435), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n457), .A3(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n238), .A3(new_n217), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n446), .A2(new_n442), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n445), .A2(new_n462), .A3(G116), .ZN(new_n463));
  OAI211_X1 g277(.A(G113), .B(new_n463), .C1(new_n454), .C2(new_n462), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n263), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G122), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n460), .A2(new_n467), .A3(new_n465), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n472), .A3(new_n468), .ZN(new_n473));
  OAI21_X1  g287(.A(G125), .B1(new_n239), .B2(new_n244), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n223), .A2(new_n265), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n231), .A2(new_n268), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n324), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n193), .A2(G224), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n478), .B(new_n479), .Z(new_n480));
  AND3_X1   g294(.A1(new_n471), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n464), .A2(new_n461), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n262), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n465), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT81), .B(KEYINPUT8), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n467), .B(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT7), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n479), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n478), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT83), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT7), .B1(new_n479), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n494), .B2(new_n479), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n474), .A2(new_n477), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n474), .A2(new_n477), .A3(KEYINPUT84), .A4(new_n496), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n488), .A2(new_n493), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n470), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n190), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n434), .B1(new_n481), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n500), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n486), .B1(new_n483), .B2(new_n465), .ZN(new_n506));
  INV_X1    g320(.A(new_n493), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n508), .B2(new_n470), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n471), .A2(new_n473), .A3(new_n480), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n433), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n432), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  AND4_X1   g326(.A1(new_n188), .A2(new_n304), .A3(new_n430), .A4(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G472), .A2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n273), .A2(new_n274), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n241), .A2(new_n242), .B1(new_n218), .B2(G146), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n518), .A2(new_n232), .B1(new_n519), .B2(new_n224), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT66), .B1(new_n249), .B2(G134), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n251), .A3(G137), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n249), .A2(G134), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G131), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n285), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n260), .A2(new_n520), .B1(new_n269), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n459), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n446), .A2(new_n447), .A3(new_n442), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n457), .B1(new_n454), .B2(KEYINPUT68), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n448), .A2(KEYINPUT70), .A3(new_n458), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT28), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n526), .A2(new_n285), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n475), .A2(new_n476), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n245), .A2(new_n286), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n535), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n529), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n310), .A2(G210), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT27), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT26), .B(G101), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n243), .A2(new_n219), .B1(G128), .B2(new_n264), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n285), .B(new_n526), .C1(new_n272), .C2(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n226), .B(new_n234), .C1(new_n255), .C2(new_n259), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n549), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n459), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n535), .A2(new_n539), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n546), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n554), .A2(KEYINPUT31), .A3(new_n555), .A4(new_n546), .ZN(new_n559));
  AOI221_X4 g373(.A(KEYINPUT71), .B1(new_n542), .B2(new_n547), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n559), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n542), .A2(new_n547), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n517), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n535), .A2(new_n539), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n540), .B2(new_n541), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT29), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n547), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(G902), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n554), .A2(new_n555), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n547), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n529), .B(new_n546), .C1(new_n540), .C2(new_n541), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n574), .B(new_n570), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n572), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n528), .B1(new_n534), .B2(new_n533), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n528), .A2(KEYINPUT30), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n584), .B2(new_n459), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT31), .B1(new_n585), .B2(new_n546), .ZN(new_n586));
  INV_X1    g400(.A(new_n559), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n563), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT71), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n562), .A2(new_n561), .A3(new_n563), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n515), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n565), .B(new_n580), .C1(new_n591), .C2(KEYINPUT32), .ZN(new_n592));
  INV_X1    g406(.A(new_n330), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT73), .B(KEYINPUT23), .Z(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(G128), .B2(new_n445), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n445), .A2(G128), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n391), .A2(KEYINPUT23), .A3(G119), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G110), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n596), .B1(new_n443), .B2(G128), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT24), .B(G110), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n593), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n601), .ZN(new_n604));
  INV_X1    g418(.A(G110), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n595), .A2(new_n605), .A3(new_n596), .A4(new_n597), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n328), .B1(new_n220), .B2(new_n345), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT74), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT22), .B(G137), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n603), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n603), .B2(new_n609), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n409), .B1(G234), .B2(new_n190), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(G902), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT77), .Z(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n616), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT75), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n190), .A4(new_n614), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT76), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT25), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n615), .A2(new_n616), .A3(G902), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT75), .B1(new_n625), .B2(KEYINPUT25), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n618), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n621), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n513), .A2(new_n592), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  INV_X1    g447(.A(new_n188), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n634), .B(new_n630), .C1(new_n297), .C2(new_n303), .ZN(new_n635));
  INV_X1    g449(.A(G472), .ZN(new_n636));
  OAI221_X1 g450(.A(new_n190), .B1(KEYINPUT94), .B2(new_n636), .C1(new_n560), .C2(new_n564), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n190), .B1(new_n560), .B2(new_n564), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n636), .A2(KEYINPUT94), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n635), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT96), .B(G478), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n414), .A2(new_n418), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT33), .B1(new_n411), .B2(new_n412), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n402), .A2(new_n408), .ZN(new_n646));
  INV_X1    g460(.A(new_n410), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n402), .A2(new_n408), .A3(new_n410), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n415), .A2(G902), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n644), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n653), .ZN(new_n655));
  AOI211_X1 g469(.A(KEYINPUT95), .B(new_n655), .C1(new_n645), .C2(new_n651), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n643), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n374), .B2(new_n375), .ZN(new_n658));
  INV_X1    g472(.A(new_n511), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n433), .B1(new_n509), .B2(new_n510), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n431), .B(new_n428), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n641), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT97), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n419), .A2(new_n420), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n373), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n362), .A2(KEYINPUT99), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n361), .A2(new_n669), .A3(KEYINPUT20), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n364), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n364), .A2(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n667), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n675), .A2(new_n676), .A3(new_n512), .A4(new_n428), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n671), .ZN(new_n678));
  INV_X1    g492(.A(new_n667), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT100), .B1(new_n680), .B2(new_n661), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n641), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT35), .B(G107), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  NAND2_X1  g498(.A1(new_n603), .A2(new_n609), .ZN(new_n685));
  INV_X1    g499(.A(new_n613), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(KEYINPUT36), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n620), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n626), .B2(new_n629), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n640), .A2(new_n637), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT101), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n640), .A2(new_n637), .A3(new_n693), .A4(new_n690), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n692), .A2(new_n513), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT37), .B(G110), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G12));
  AND3_X1   g511(.A1(new_n304), .A2(new_n188), .A3(new_n512), .ZN(new_n698));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n425), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n423), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n680), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n592), .A2(new_n698), .A3(new_n690), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n705));
  INV_X1    g519(.A(new_n690), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n589), .A2(new_n590), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n707), .A2(new_n517), .B1(G472), .B2(new_n579), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n514), .B1(new_n560), .B2(new_n564), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n516), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n706), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n698), .A4(new_n703), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT103), .B(G128), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G30));
  OAI21_X1  g530(.A(new_n666), .B1(new_n374), .B2(new_n375), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n717), .A2(new_n432), .A3(new_n690), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n504), .A2(KEYINPUT38), .A3(new_n511), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT38), .B1(new_n504), .B2(new_n511), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n591), .A2(KEYINPUT32), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n581), .A2(new_n546), .ZN(new_n725));
  AOI21_X1  g539(.A(G902), .B1(new_n725), .B2(new_n567), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n573), .A2(new_n546), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n636), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n565), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n723), .B1(new_n724), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n710), .A2(KEYINPUT104), .A3(new_n565), .A4(new_n729), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n634), .B1(new_n297), .B2(new_n303), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n701), .B(KEYINPUT39), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n739));
  AOI211_X1 g553(.A(new_n722), .B(new_n734), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n218), .ZN(G45));
  AND3_X1   g555(.A1(new_n592), .A2(new_n698), .A3(new_n690), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n657), .B(new_n701), .C1(new_n374), .C2(new_n375), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT105), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n365), .A2(new_n373), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT90), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n365), .A2(new_n366), .A3(new_n373), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n657), .A4(new_n701), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  AOI21_X1  g567(.A(new_n630), .B1(new_n708), .B2(new_n710), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n661), .A2(new_n658), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n248), .A2(new_n277), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n286), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n293), .B1(new_n757), .B2(new_n294), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n189), .B(new_n190), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n188), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n190), .B1(new_n758), .B2(new_n759), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n189), .B1(new_n762), .B2(KEYINPUT106), .ZN(new_n763));
  AOI211_X1 g577(.A(KEYINPUT106), .B(G902), .C1(new_n280), .C2(new_n295), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n761), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n754), .A2(new_n755), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT41), .B(G113), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G15));
  NAND2_X1  g583(.A1(new_n681), .A2(new_n677), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n754), .A3(new_n766), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G116), .ZN(G18));
  AOI21_X1  g586(.A(new_n634), .B1(new_n296), .B2(new_n189), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n774));
  OAI21_X1  g588(.A(G469), .B1(new_n296), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n775), .B2(new_n764), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n431), .B1(new_n659), .B2(new_n660), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n592), .A2(new_n778), .A3(new_n430), .A4(new_n690), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G119), .ZN(G21));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n777), .B2(new_n717), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n512), .A2(new_n748), .A3(KEYINPUT107), .A4(new_n666), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n568), .A2(new_n547), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n515), .B1(new_n562), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n630), .B(new_n786), .C1(new_n638), .C2(G472), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n787), .A3(new_n428), .A4(new_n766), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G122), .ZN(G24));
  NAND4_X1  g603(.A1(new_n744), .A2(new_n750), .A3(new_n766), .A4(new_n512), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n638), .A2(G472), .ZN(new_n791));
  INV_X1    g605(.A(new_n786), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n690), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT108), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n786), .B(new_n706), .C1(new_n638), .C2(G472), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n751), .A2(new_n795), .A3(new_n796), .A4(new_n778), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G125), .ZN(G27));
  XOR2_X1   g613(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n504), .A2(new_n431), .A3(new_n511), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n304), .A2(new_n188), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n592), .A2(new_n803), .A3(new_n631), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n744), .A2(new_n750), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n754), .A2(new_n751), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G131), .ZN(G33));
  NAND4_X1  g625(.A1(new_n592), .A2(new_n803), .A3(new_n631), .A4(new_n703), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT110), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n754), .A2(new_n814), .A3(new_n703), .A4(new_n803), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G134), .ZN(G36));
  AOI21_X1  g631(.A(new_n706), .B1(new_n640), .B2(new_n637), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n657), .A2(new_n746), .A3(new_n747), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(KEYINPUT43), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(KEYINPUT43), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n818), .A2(new_n822), .A3(KEYINPUT44), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT44), .B1(new_n822), .B2(new_n818), .ZN(new_n824));
  INV_X1    g638(.A(new_n802), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n292), .A2(new_n294), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT80), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n292), .A2(KEYINPUT80), .A3(new_n294), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n293), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n827), .B1(new_n832), .B2(new_n301), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n300), .A2(KEYINPUT45), .A3(new_n302), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n834), .A3(G469), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT111), .A4(G469), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n191), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n760), .B1(new_n839), .B2(KEYINPUT46), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT46), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n841), .B(new_n191), .C1(new_n837), .C2(new_n838), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n188), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  INV_X1    g658(.A(new_n736), .ZN(new_n845));
  OR3_X1    g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n826), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(KEYINPUT113), .B(G137), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(G39));
  OR4_X1    g664(.A1(new_n592), .A2(new_n805), .A3(new_n631), .A4(new_n825), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT47), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(KEYINPUT47), .B(new_n188), .C1(new_n840), .C2(new_n842), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(new_n322), .ZN(G42));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT120), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n820), .A2(new_n821), .A3(new_n423), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n721), .A2(new_n776), .A3(new_n431), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n787), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT50), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n861), .A2(new_n787), .A3(KEYINPUT50), .A4(new_n862), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n825), .A2(new_n776), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n795), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n861), .A2(KEYINPUT118), .A3(new_n795), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n776), .A2(new_n630), .A3(new_n423), .A4(new_n825), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n748), .A2(new_n657), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n734), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n867), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n760), .B1(new_n775), .B2(new_n764), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n878), .A2(new_n188), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n853), .A2(new_n854), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n861), .A2(new_n787), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n881), .A2(new_n802), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n877), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT51), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n861), .A2(new_n754), .A3(new_n868), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT48), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n734), .A2(new_n748), .A3(new_n657), .A4(new_n874), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n881), .A2(new_n778), .ZN(new_n890));
  AND4_X1   g704(.A1(new_n421), .A2(new_n888), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n883), .B2(KEYINPUT51), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n884), .B1(new_n883), .B2(KEYINPUT51), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n886), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n373), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n666), .A2(new_n895), .A3(new_n702), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n592), .A2(new_n678), .A3(new_n690), .A4(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n793), .A2(new_n805), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n803), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n810), .A2(new_n816), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n746), .A2(new_n747), .A3(new_n666), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n661), .B1(new_n658), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(new_n635), .A3(new_n637), .A4(new_n640), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n632), .A2(new_n779), .A3(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n754), .B(new_n766), .C1(new_n770), .C2(new_n755), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n695), .A3(new_n788), .A4(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n713), .A2(new_n705), .B1(new_n794), .B2(new_n797), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n689), .B(new_n701), .C1(new_n626), .C2(new_n629), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n304), .A2(new_n188), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT116), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT116), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n735), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n784), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n916), .A2(new_n733), .B1(new_n742), .B2(new_n751), .ZN(new_n917));
  XNOR2_X1  g731(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n909), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n909), .B2(new_n917), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n907), .B(new_n908), .C1(new_n919), .C2(new_n922), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n806), .A2(new_n809), .B1(new_n813), .B2(new_n815), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n692), .A2(new_n513), .A3(new_n694), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n632), .A2(new_n779), .A3(new_n903), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n905), .A2(new_n788), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n924), .A2(new_n927), .A3(new_n928), .A4(new_n899), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n917), .A2(new_n714), .A3(new_n798), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT52), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n909), .A2(KEYINPUT52), .A3(new_n917), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n923), .B(KEYINPUT54), .C1(new_n934), .C2(new_n908), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n907), .B(KEYINPUT53), .C1(new_n919), .C2(new_n922), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n936), .B(new_n937), .C1(new_n934), .C2(KEYINPUT53), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n860), .B1(new_n894), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n631), .A2(new_n188), .A3(new_n431), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n819), .B(new_n941), .C1(KEYINPUT49), .C2(new_n878), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT114), .ZN(new_n943));
  INV_X1    g757(.A(new_n721), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n878), .A2(KEYINPUT49), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT115), .Z(new_n946));
  NAND4_X1  g760(.A1(new_n943), .A2(new_n734), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n857), .B1(new_n940), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n893), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n883), .A2(KEYINPUT51), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n951), .A3(new_n885), .A4(new_n891), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n935), .A2(new_n938), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n859), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(KEYINPUT121), .A3(new_n947), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n949), .A2(new_n955), .ZN(G75));
  INV_X1    g770(.A(new_n933), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT52), .B1(new_n909), .B2(new_n917), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n907), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n908), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n190), .B1(new_n960), .B2(new_n936), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(G210), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n471), .A2(new_n473), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(new_n480), .Z(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(KEYINPUT123), .A2(KEYINPUT56), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n962), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n967), .B1(new_n962), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n193), .A2(G952), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(G51));
  OAI21_X1  g786(.A(new_n936), .B1(new_n934), .B2(KEYINPUT53), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT54), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n938), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n191), .B(KEYINPUT57), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n758), .B2(new_n759), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n961), .A2(new_n837), .A3(new_n838), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n971), .B1(new_n978), .B2(new_n979), .ZN(G54));
  NAND3_X1  g794(.A1(new_n961), .A2(KEYINPUT58), .A3(G475), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n350), .A2(new_n360), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n983), .A2(new_n984), .A3(new_n971), .ZN(G60));
  NAND2_X1  g799(.A1(G478), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT59), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n652), .B1(new_n953), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n987), .B1(new_n645), .B2(new_n651), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n971), .B(new_n989), .C1(new_n975), .C2(new_n990), .ZN(G63));
  XNOR2_X1  g805(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(G217), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT60), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n973), .A2(KEYINPUT124), .A3(new_n688), .A4(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n971), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n995), .B1(new_n960), .B2(new_n936), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n997), .B(new_n998), .C1(new_n617), .C2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT124), .B1(new_n999), .B2(new_n688), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n993), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n973), .A2(new_n996), .ZN(new_n1003));
  INV_X1    g817(.A(new_n617), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n971), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n973), .A2(new_n688), .A3(new_n996), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT124), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1005), .A2(new_n1008), .A3(new_n997), .A4(new_n992), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1002), .A2(new_n1009), .ZN(G66));
  INV_X1    g824(.A(G224), .ZN(new_n1011));
  OAI21_X1  g825(.A(G953), .B1(new_n426), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n906), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(G953), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n963), .B1(G898), .B2(new_n193), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(G69));
  NOR2_X1   g830(.A1(new_n848), .A2(new_n855), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n846), .A2(new_n847), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1018), .A2(new_n754), .A3(new_n784), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT127), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n924), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n924), .A2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n909), .A2(new_n752), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1017), .A2(new_n1019), .A3(new_n193), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n352), .A2(new_n353), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT126), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n584), .B(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(G900), .B2(G953), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n740), .A2(new_n1023), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT62), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n825), .B1(new_n658), .B2(new_n901), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n754), .A2(new_n737), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1034), .A2(new_n1017), .A3(new_n1036), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n1037), .A2(new_n193), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1028), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1030), .B(new_n1032), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1030), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1039), .B1(new_n1037), .B2(new_n193), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1031), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1040), .A2(new_n1043), .ZN(G72));
  NAND4_X1  g858(.A1(new_n1034), .A2(new_n1013), .A3(new_n1017), .A4(new_n1036), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  AOI21_X1  g861(.A(new_n727), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n725), .A2(new_n554), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n1017), .A2(new_n1019), .A3(new_n1013), .A4(new_n1024), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1049), .B1(new_n1050), .B2(new_n1047), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1047), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1052), .B1(new_n574), .B2(new_n556), .ZN(new_n1053));
  OAI211_X1 g867(.A(new_n923), .B(new_n1053), .C1(new_n934), .C2(new_n908), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(new_n998), .ZN(new_n1055));
  NOR3_X1   g869(.A1(new_n1048), .A2(new_n1051), .A3(new_n1055), .ZN(G57));
endmodule


