

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(KEYINPUT101), .B(n750), .ZN(n773) );
  NOR2_X4 U552 ( .A1(G2105), .A2(n532), .ZN(n989) );
  NOR2_X2 U553 ( .A1(n540), .A2(n539), .ZN(G160) );
  INV_X1 U554 ( .A(KEYINPUT29), .ZN(n771) );
  XNOR2_X1 U555 ( .A(n772), .B(n771), .ZN(n778) );
  NOR2_X1 U556 ( .A1(n821), .A2(n820), .ZN(n823) );
  NOR2_X1 U557 ( .A1(G651), .A2(n630), .ZN(n657) );
  NOR2_X1 U558 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U559 ( .A1(n647), .A2(G89), .ZN(n517) );
  XNOR2_X1 U560 ( .A(n517), .B(KEYINPUT4), .ZN(n519) );
  XOR2_X1 U561 ( .A(G543), .B(KEYINPUT0), .Z(n630) );
  INV_X1 U562 ( .A(G651), .ZN(n521) );
  NOR2_X1 U563 ( .A1(n630), .A2(n521), .ZN(n651) );
  NAND2_X1 U564 ( .A1(G76), .A2(n651), .ZN(n518) );
  NAND2_X1 U565 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U566 ( .A(n520), .B(KEYINPUT5), .ZN(n528) );
  NAND2_X1 U567 ( .A1(G51), .A2(n657), .ZN(n525) );
  NOR2_X1 U568 ( .A1(G543), .A2(n521), .ZN(n522) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n522), .Z(n523) );
  XNOR2_X1 U570 ( .A(KEYINPUT68), .B(n523), .ZN(n648) );
  NAND2_X1 U571 ( .A1(G63), .A2(n648), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U573 ( .A(KEYINPUT6), .B(n526), .Z(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U575 ( .A(n529), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U576 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U577 ( .A(G2104), .ZN(n532) );
  NAND2_X1 U578 ( .A1(G101), .A2(n989), .ZN(n530) );
  XNOR2_X1 U579 ( .A(n530), .B(KEYINPUT23), .ZN(n531) );
  XNOR2_X1 U580 ( .A(KEYINPUT67), .B(n531), .ZN(n535) );
  AND2_X1 U581 ( .A1(n532), .A2(G2105), .ZN(n984) );
  NAND2_X1 U582 ( .A1(G125), .A2(n984), .ZN(n533) );
  XNOR2_X1 U583 ( .A(n533), .B(KEYINPUT66), .ZN(n534) );
  NAND2_X1 U584 ( .A1(n535), .A2(n534), .ZN(n540) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n985) );
  NAND2_X1 U586 ( .A1(G113), .A2(n985), .ZN(n538) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  XOR2_X2 U588 ( .A(KEYINPUT17), .B(n536), .Z(n988) );
  NAND2_X1 U589 ( .A1(G137), .A2(n988), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G85), .A2(n647), .ZN(n542) );
  NAND2_X1 U592 ( .A1(G60), .A2(n648), .ZN(n541) );
  NAND2_X1 U593 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U594 ( .A1(G72), .A2(n651), .ZN(n544) );
  NAND2_X1 U595 ( .A1(G47), .A2(n657), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U597 ( .A1(n546), .A2(n545), .ZN(G290) );
  XNOR2_X1 U598 ( .A(G1341), .B(G2427), .ZN(n556) );
  XOR2_X1 U599 ( .A(G2451), .B(KEYINPUT107), .Z(n548) );
  XNOR2_X1 U600 ( .A(G1348), .B(G2443), .ZN(n547) );
  XNOR2_X1 U601 ( .A(n548), .B(n547), .ZN(n552) );
  XOR2_X1 U602 ( .A(G2438), .B(G2435), .Z(n550) );
  XNOR2_X1 U603 ( .A(G2430), .B(G2454), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U605 ( .A(n552), .B(n551), .Z(n554) );
  XNOR2_X1 U606 ( .A(G2446), .B(KEYINPUT108), .ZN(n553) );
  XNOR2_X1 U607 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U608 ( .A(n556), .B(n555), .ZN(n557) );
  AND2_X1 U609 ( .A1(n557), .A2(G14), .ZN(G401) );
  NAND2_X1 U610 ( .A1(G52), .A2(n657), .ZN(n559) );
  NAND2_X1 U611 ( .A1(G64), .A2(n648), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n559), .A2(n558), .ZN(n564) );
  NAND2_X1 U613 ( .A1(G90), .A2(n647), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G77), .A2(n651), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U617 ( .A1(n564), .A2(n563), .ZN(G171) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G108), .ZN(G238) );
  INV_X1 U620 ( .A(G120), .ZN(G236) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U623 ( .A(n565), .B(KEYINPUT10), .ZN(n566) );
  XNOR2_X1 U624 ( .A(KEYINPUT72), .B(n566), .ZN(G223) );
  INV_X1 U625 ( .A(G567), .ZN(n684) );
  NOR2_X1 U626 ( .A1(n684), .A2(G223), .ZN(n567) );
  XOR2_X1 U627 ( .A(KEYINPUT73), .B(n567), .Z(n568) );
  XNOR2_X1 U628 ( .A(KEYINPUT11), .B(n568), .ZN(G234) );
  INV_X1 U629 ( .A(G860), .ZN(n602) );
  NAND2_X1 U630 ( .A1(G56), .A2(n648), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n569), .B(KEYINPUT14), .ZN(n579) );
  NAND2_X1 U632 ( .A1(n647), .A2(G81), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G68), .A2(n651), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n573) );
  XNOR2_X1 U637 ( .A(n574), .B(n573), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G43), .A2(n657), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT75), .B(n575), .ZN(n576) );
  NOR2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U642 ( .A(n580), .B(KEYINPUT76), .ZN(n956) );
  OR2_X1 U643 ( .A1(n602), .A2(n956), .ZN(G153) );
  INV_X1 U644 ( .A(G868), .ZN(n669) );
  NOR2_X1 U645 ( .A1(n669), .A2(G171), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT77), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G92), .A2(n647), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G66), .A2(n648), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G79), .A2(n651), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G54), .A2(n657), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n588), .Z(n953) );
  INV_X1 U655 ( .A(n953), .ZN(n764) );
  NAND2_X1 U656 ( .A1(n669), .A2(n764), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G53), .A2(n657), .ZN(n591) );
  XOR2_X1 U659 ( .A(KEYINPUT70), .B(n591), .Z(n598) );
  NAND2_X1 U660 ( .A1(G91), .A2(n647), .ZN(n593) );
  NAND2_X1 U661 ( .A1(G78), .A2(n651), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U663 ( .A(n594), .B(KEYINPUT69), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G65), .A2(n648), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U667 ( .A(KEYINPUT71), .B(n599), .ZN(G299) );
  NAND2_X1 U668 ( .A1(G286), .A2(G868), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G299), .A2(n669), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U671 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n603), .A2(n953), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(n956), .A2(G868), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G868), .A2(n953), .ZN(n605) );
  NOR2_X1 U676 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U678 ( .A1(n988), .A2(G135), .ZN(n608) );
  XNOR2_X1 U679 ( .A(KEYINPUT78), .B(n608), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n984), .A2(G123), .ZN(n609) );
  XNOR2_X1 U681 ( .A(KEYINPUT18), .B(n609), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n612), .B(KEYINPUT79), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G99), .A2(n989), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n985), .A2(G111), .ZN(n615) );
  XOR2_X1 U687 ( .A(KEYINPUT80), .B(n615), .Z(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n999) );
  XNOR2_X1 U689 ( .A(n999), .B(G2096), .ZN(n619) );
  INV_X1 U690 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U692 ( .A1(G559), .A2(n953), .ZN(n620) );
  XNOR2_X1 U693 ( .A(n620), .B(n956), .ZN(n666) );
  NOR2_X1 U694 ( .A1(n666), .A2(G860), .ZN(n629) );
  NAND2_X1 U695 ( .A1(G93), .A2(n647), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G67), .A2(n648), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G80), .A2(n651), .ZN(n623) );
  XNOR2_X1 U699 ( .A(KEYINPUT81), .B(n623), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n657), .A2(G55), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n668) );
  XOR2_X1 U703 ( .A(n668), .B(KEYINPUT82), .Z(n628) );
  XNOR2_X1 U704 ( .A(n629), .B(n628), .ZN(G145) );
  NAND2_X1 U705 ( .A1(n657), .A2(G49), .ZN(n635) );
  NAND2_X1 U706 ( .A1(G87), .A2(n630), .ZN(n632) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U709 ( .A1(n648), .A2(n633), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U711 ( .A(KEYINPUT83), .B(n636), .Z(G288) );
  NAND2_X1 U712 ( .A1(n647), .A2(G88), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(KEYINPUT88), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G75), .A2(n651), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U716 ( .A(KEYINPUT89), .B(n640), .ZN(n646) );
  NAND2_X1 U717 ( .A1(G50), .A2(n657), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n641), .B(KEYINPUT87), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G62), .A2(n648), .ZN(n642) );
  XOR2_X1 U720 ( .A(KEYINPUT86), .B(n642), .Z(n643) );
  NOR2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(G303) );
  INV_X1 U723 ( .A(G303), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G86), .A2(n647), .ZN(n650) );
  NAND2_X1 U725 ( .A1(G61), .A2(n648), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n656) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n653) );
  NAND2_X1 U728 ( .A1(G73), .A2(n651), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U730 ( .A(KEYINPUT84), .B(n654), .Z(n655) );
  NOR2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n657), .A2(G48), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(G305) );
  XOR2_X1 U734 ( .A(KEYINPUT90), .B(KEYINPUT19), .Z(n660) );
  XNOR2_X1 U735 ( .A(G290), .B(n660), .ZN(n661) );
  XNOR2_X1 U736 ( .A(G288), .B(n661), .ZN(n663) );
  INV_X1 U737 ( .A(G299), .ZN(n747) );
  XNOR2_X1 U738 ( .A(n747), .B(G166), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n664), .B(G305), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(n668), .ZN(n952) );
  XNOR2_X1 U742 ( .A(n666), .B(n952), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U744 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XNOR2_X1 U747 ( .A(n672), .B(KEYINPUT91), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n673), .B(KEYINPUT20), .ZN(n674) );
  NAND2_X1 U749 ( .A1(n674), .A2(G2090), .ZN(n675) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U753 ( .A1(G132), .A2(G82), .ZN(n677) );
  XNOR2_X1 U754 ( .A(n677), .B(KEYINPUT92), .ZN(n678) );
  XNOR2_X1 U755 ( .A(n678), .B(KEYINPUT22), .ZN(n679) );
  NOR2_X1 U756 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U757 ( .A1(G96), .A2(n680), .ZN(n832) );
  NAND2_X1 U758 ( .A1(G2106), .A2(n832), .ZN(n681) );
  XNOR2_X1 U759 ( .A(n681), .B(KEYINPUT93), .ZN(n686) );
  NOR2_X1 U760 ( .A1(G236), .A2(G238), .ZN(n682) );
  NAND2_X1 U761 ( .A1(G69), .A2(n682), .ZN(n683) );
  NOR2_X1 U762 ( .A1(G237), .A2(n683), .ZN(n831) );
  NOR2_X1 U763 ( .A1(n684), .A2(n831), .ZN(n685) );
  NOR2_X1 U764 ( .A1(n686), .A2(n685), .ZN(G319) );
  INV_X1 U765 ( .A(G319), .ZN(n1009) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U767 ( .A1(n1009), .A2(n687), .ZN(n830) );
  NAND2_X1 U768 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G102), .A2(n989), .ZN(n688) );
  XNOR2_X1 U770 ( .A(n688), .B(KEYINPUT96), .ZN(n691) );
  NAND2_X1 U771 ( .A1(G114), .A2(n985), .ZN(n689) );
  XOR2_X1 U772 ( .A(KEYINPUT95), .B(n689), .Z(n690) );
  NAND2_X1 U773 ( .A1(n691), .A2(n690), .ZN(n696) );
  NAND2_X1 U774 ( .A1(n984), .A2(G126), .ZN(n692) );
  XNOR2_X1 U775 ( .A(n692), .B(KEYINPUT94), .ZN(n694) );
  NAND2_X1 U776 ( .A1(G138), .A2(n988), .ZN(n693) );
  NAND2_X1 U777 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U778 ( .A1(n696), .A2(n695), .ZN(G164) );
  NAND2_X1 U779 ( .A1(G104), .A2(n989), .ZN(n698) );
  NAND2_X1 U780 ( .A1(G140), .A2(n988), .ZN(n697) );
  NAND2_X1 U781 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U782 ( .A(KEYINPUT34), .B(n699), .ZN(n705) );
  NAND2_X1 U783 ( .A1(n984), .A2(G128), .ZN(n700) );
  XOR2_X1 U784 ( .A(KEYINPUT97), .B(n700), .Z(n702) );
  NAND2_X1 U785 ( .A1(n985), .A2(G116), .ZN(n701) );
  NAND2_X1 U786 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U787 ( .A(KEYINPUT35), .B(n703), .Z(n704) );
  NOR2_X1 U788 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U789 ( .A(KEYINPUT36), .B(n706), .ZN(n1005) );
  XNOR2_X1 U790 ( .A(G2067), .B(KEYINPUT37), .ZN(n729) );
  NOR2_X1 U791 ( .A1(n1005), .A2(n729), .ZN(n845) );
  NOR2_X1 U792 ( .A1(G164), .A2(G1384), .ZN(n737) );
  NAND2_X1 U793 ( .A1(G160), .A2(G40), .ZN(n736) );
  NOR2_X1 U794 ( .A1(n737), .A2(n736), .ZN(n733) );
  NAND2_X1 U795 ( .A1(n845), .A2(n733), .ZN(n822) );
  NAND2_X1 U796 ( .A1(G129), .A2(n984), .ZN(n708) );
  NAND2_X1 U797 ( .A1(G141), .A2(n988), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n989), .A2(G105), .ZN(n709) );
  XOR2_X1 U800 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n985), .A2(G117), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n978) );
  NOR2_X1 U804 ( .A1(G1996), .A2(n978), .ZN(n842) );
  NAND2_X1 U805 ( .A1(G1996), .A2(n978), .ZN(n722) );
  NAND2_X1 U806 ( .A1(G95), .A2(n989), .ZN(n715) );
  NAND2_X1 U807 ( .A1(G131), .A2(n988), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n984), .A2(G119), .ZN(n716) );
  XOR2_X1 U810 ( .A(KEYINPUT98), .B(n716), .Z(n717) );
  NOR2_X1 U811 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n985), .A2(G107), .ZN(n719) );
  NAND2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n979) );
  NAND2_X1 U814 ( .A1(G1991), .A2(n979), .ZN(n721) );
  NAND2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n861) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n723) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n979), .ZN(n862) );
  NOR2_X1 U818 ( .A1(n723), .A2(n862), .ZN(n724) );
  NOR2_X1 U819 ( .A1(n861), .A2(n724), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n842), .A2(n725), .ZN(n726) );
  XOR2_X1 U821 ( .A(n726), .B(KEYINPUT105), .Z(n727) );
  XNOR2_X1 U822 ( .A(KEYINPUT39), .B(n727), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n822), .A2(n728), .ZN(n730) );
  NAND2_X1 U824 ( .A1(n1005), .A2(n729), .ZN(n846) );
  NAND2_X1 U825 ( .A1(n730), .A2(n846), .ZN(n731) );
  NAND2_X1 U826 ( .A1(n731), .A2(n733), .ZN(n732) );
  XNOR2_X1 U827 ( .A(n732), .B(KEYINPUT106), .ZN(n825) );
  INV_X1 U828 ( .A(n733), .ZN(n735) );
  XNOR2_X1 U829 ( .A(G1986), .B(G290), .ZN(n905) );
  NOR2_X1 U830 ( .A1(n905), .A2(n861), .ZN(n734) );
  NOR2_X1 U831 ( .A1(n735), .A2(n734), .ZN(n821) );
  XNOR2_X1 U832 ( .A(KEYINPUT99), .B(n736), .ZN(n738) );
  NAND2_X2 U833 ( .A1(n738), .A2(n737), .ZN(n750) );
  NAND2_X1 U834 ( .A1(G8), .A2(n750), .ZN(n814) );
  NOR2_X1 U835 ( .A1(G1981), .A2(G305), .ZN(n739) );
  XOR2_X1 U836 ( .A(n739), .B(KEYINPUT24), .Z(n740) );
  NOR2_X1 U837 ( .A1(n814), .A2(n740), .ZN(n819) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n804) );
  NAND2_X1 U839 ( .A1(n804), .A2(KEYINPUT33), .ZN(n741) );
  NOR2_X1 U840 ( .A1(n814), .A2(n741), .ZN(n809) );
  NAND2_X1 U841 ( .A1(n773), .A2(G2072), .ZN(n742) );
  XNOR2_X1 U842 ( .A(n742), .B(KEYINPUT27), .ZN(n744) );
  XNOR2_X1 U843 ( .A(G1956), .B(KEYINPUT103), .ZN(n921) );
  NOR2_X1 U844 ( .A1(n921), .A2(n773), .ZN(n743) );
  NOR2_X1 U845 ( .A1(n744), .A2(n743), .ZN(n748) );
  NOR2_X1 U846 ( .A1(n748), .A2(n747), .ZN(n746) );
  INV_X1 U847 ( .A(KEYINPUT28), .ZN(n745) );
  XNOR2_X1 U848 ( .A(n746), .B(n745), .ZN(n770) );
  NAND2_X1 U849 ( .A1(n748), .A2(n747), .ZN(n768) );
  XOR2_X1 U850 ( .A(G1996), .B(KEYINPUT104), .Z(n873) );
  XNOR2_X1 U851 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n751) );
  OR2_X1 U852 ( .A1(n873), .A2(n751), .ZN(n749) );
  OR2_X1 U853 ( .A1(n750), .A2(n749), .ZN(n754) );
  OR2_X1 U854 ( .A1(n750), .A2(n873), .ZN(n752) );
  NAND2_X1 U855 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U856 ( .A1(n754), .A2(n753), .ZN(n756) );
  NAND2_X1 U857 ( .A1(n750), .A2(G1341), .ZN(n755) );
  NAND2_X1 U858 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U859 ( .A1(n956), .A2(n757), .ZN(n758) );
  XNOR2_X1 U860 ( .A(KEYINPUT65), .B(n758), .ZN(n762) );
  NAND2_X1 U861 ( .A1(n750), .A2(G1348), .ZN(n760) );
  NAND2_X1 U862 ( .A1(G2067), .A2(n773), .ZN(n759) );
  NAND2_X1 U863 ( .A1(n760), .A2(n759), .ZN(n763) );
  OR2_X1 U864 ( .A1(n764), .A2(n763), .ZN(n761) );
  NAND2_X1 U865 ( .A1(n762), .A2(n761), .ZN(n766) );
  NAND2_X1 U866 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U867 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U868 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U869 ( .A1(n770), .A2(n769), .ZN(n772) );
  XNOR2_X1 U870 ( .A(G2078), .B(KEYINPUT25), .ZN(n875) );
  NAND2_X1 U871 ( .A1(n773), .A2(n875), .ZN(n775) );
  XOR2_X1 U872 ( .A(G1961), .B(KEYINPUT100), .Z(n932) );
  NAND2_X1 U873 ( .A1(n932), .A2(n750), .ZN(n774) );
  NAND2_X1 U874 ( .A1(n775), .A2(n774), .ZN(n782) );
  NAND2_X1 U875 ( .A1(G171), .A2(n782), .ZN(n776) );
  XNOR2_X1 U876 ( .A(n776), .B(KEYINPUT102), .ZN(n777) );
  NAND2_X1 U877 ( .A1(n778), .A2(n777), .ZN(n787) );
  NOR2_X1 U878 ( .A1(G1966), .A2(n814), .ZN(n798) );
  NOR2_X1 U879 ( .A1(G2084), .A2(n750), .ZN(n795) );
  NOR2_X1 U880 ( .A1(n798), .A2(n795), .ZN(n779) );
  NAND2_X1 U881 ( .A1(G8), .A2(n779), .ZN(n780) );
  XNOR2_X1 U882 ( .A(KEYINPUT30), .B(n780), .ZN(n781) );
  NOR2_X1 U883 ( .A1(G168), .A2(n781), .ZN(n784) );
  NOR2_X1 U884 ( .A1(G171), .A2(n782), .ZN(n783) );
  NOR2_X1 U885 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U886 ( .A(KEYINPUT31), .B(n785), .Z(n786) );
  NAND2_X1 U887 ( .A1(n787), .A2(n786), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n796), .A2(G286), .ZN(n792) );
  NOR2_X1 U889 ( .A1(G2090), .A2(n750), .ZN(n789) );
  NOR2_X1 U890 ( .A1(G1971), .A2(n814), .ZN(n788) );
  NOR2_X1 U891 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U892 ( .A1(n790), .A2(G303), .ZN(n791) );
  NAND2_X1 U893 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U894 ( .A1(G8), .A2(n793), .ZN(n794) );
  XNOR2_X1 U895 ( .A(n794), .B(KEYINPUT32), .ZN(n802) );
  NAND2_X1 U896 ( .A1(G8), .A2(n795), .ZN(n800) );
  INV_X1 U897 ( .A(n796), .ZN(n797) );
  NOR2_X1 U898 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U899 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n813) );
  NOR2_X1 U901 ( .A1(G1971), .A2(G303), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n900) );
  NAND2_X1 U903 ( .A1(n813), .A2(n900), .ZN(n805) );
  NAND2_X1 U904 ( .A1(G1976), .A2(G288), .ZN(n906) );
  NAND2_X1 U905 ( .A1(n805), .A2(n906), .ZN(n806) );
  NOR2_X1 U906 ( .A1(n814), .A2(n806), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n807), .A2(KEYINPUT33), .ZN(n808) );
  NOR2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U909 ( .A(G1981), .B(G305), .Z(n896) );
  NAND2_X1 U910 ( .A1(n810), .A2(n896), .ZN(n817) );
  NOR2_X1 U911 ( .A1(G2090), .A2(G303), .ZN(n811) );
  NAND2_X1 U912 ( .A1(G8), .A2(n811), .ZN(n812) );
  NAND2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U919 ( .A(KEYINPUT40), .B(n826), .ZN(G329) );
  INV_X1 U920 ( .A(G223), .ZN(n827) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U923 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U926 ( .A(n831), .ZN(n833) );
  NOR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G325) );
  XNOR2_X1 U928 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  NAND2_X1 U930 ( .A1(G124), .A2(n984), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT44), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n989), .A2(G100), .ZN(n835) );
  NAND2_X1 U933 ( .A1(n836), .A2(n835), .ZN(n840) );
  NAND2_X1 U934 ( .A1(G112), .A2(n985), .ZN(n838) );
  NAND2_X1 U935 ( .A1(G136), .A2(n988), .ZN(n837) );
  NAND2_X1 U936 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U937 ( .A1(n840), .A2(n839), .ZN(G162) );
  INV_X1 U938 ( .A(G171), .ZN(G301) );
  XOR2_X1 U939 ( .A(G2090), .B(G162), .Z(n841) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n843), .B(KEYINPUT51), .ZN(n844) );
  NOR2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n847) );
  NAND2_X1 U943 ( .A1(n847), .A2(n846), .ZN(n860) );
  NAND2_X1 U944 ( .A1(G103), .A2(n989), .ZN(n849) );
  NAND2_X1 U945 ( .A1(G139), .A2(n988), .ZN(n848) );
  NAND2_X1 U946 ( .A1(n849), .A2(n848), .ZN(n854) );
  NAND2_X1 U947 ( .A1(G127), .A2(n984), .ZN(n851) );
  NAND2_X1 U948 ( .A1(G115), .A2(n985), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(KEYINPUT47), .B(n852), .Z(n853) );
  NOR2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n1000) );
  XOR2_X1 U952 ( .A(G2072), .B(n1000), .Z(n856) );
  XOR2_X1 U953 ( .A(G164), .B(G2078), .Z(n855) );
  NOR2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(KEYINPUT118), .B(n857), .Z(n858) );
  XNOR2_X1 U956 ( .A(KEYINPUT50), .B(n858), .ZN(n859) );
  NOR2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n867) );
  XNOR2_X1 U958 ( .A(G160), .B(G2084), .ZN(n864) );
  NOR2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U961 ( .A1(n865), .A2(n999), .ZN(n866) );
  NAND2_X1 U962 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U963 ( .A(KEYINPUT52), .B(n868), .ZN(n869) );
  XNOR2_X1 U964 ( .A(KEYINPUT119), .B(n869), .ZN(n871) );
  INV_X1 U965 ( .A(KEYINPUT55), .ZN(n870) );
  NAND2_X1 U966 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U967 ( .A1(n872), .A2(G29), .ZN(n950) );
  XOR2_X1 U968 ( .A(G29), .B(KEYINPUT122), .Z(n894) );
  XNOR2_X1 U969 ( .A(n873), .B(G32), .ZN(n885) );
  XNOR2_X1 U970 ( .A(KEYINPUT121), .B(G2067), .ZN(n874) );
  XNOR2_X1 U971 ( .A(n874), .B(G26), .ZN(n880) );
  XNOR2_X1 U972 ( .A(G27), .B(n875), .ZN(n876) );
  NAND2_X1 U973 ( .A1(n876), .A2(G28), .ZN(n878) );
  XNOR2_X1 U974 ( .A(G33), .B(G2072), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U976 ( .A1(n880), .A2(n879), .ZN(n883) );
  XNOR2_X1 U977 ( .A(G25), .B(G1991), .ZN(n881) );
  XNOR2_X1 U978 ( .A(KEYINPUT120), .B(n881), .ZN(n882) );
  NOR2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n884) );
  NAND2_X1 U980 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U981 ( .A(n886), .B(KEYINPUT53), .ZN(n889) );
  XOR2_X1 U982 ( .A(G2084), .B(G34), .Z(n887) );
  XNOR2_X1 U983 ( .A(KEYINPUT54), .B(n887), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U985 ( .A(G35), .B(G2090), .ZN(n890) );
  NOR2_X1 U986 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n892), .B(KEYINPUT55), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n895) );
  NAND2_X1 U989 ( .A1(G11), .A2(n895), .ZN(n948) );
  XNOR2_X1 U990 ( .A(G16), .B(KEYINPUT56), .ZN(n917) );
  XNOR2_X1 U991 ( .A(G1966), .B(G168), .ZN(n897) );
  NAND2_X1 U992 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n898), .B(KEYINPUT57), .ZN(n915) );
  NAND2_X1 U994 ( .A1(G1971), .A2(G303), .ZN(n899) );
  NAND2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n902) );
  XNOR2_X1 U996 ( .A(G1961), .B(G301), .ZN(n901) );
  NOR2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n911) );
  XNOR2_X1 U998 ( .A(n953), .B(G1348), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n903), .B(KEYINPUT123), .ZN(n909) );
  XNOR2_X1 U1000 ( .A(G1956), .B(G299), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(n911), .A2(n910), .ZN(n913) );
  XNOR2_X1 U1005 ( .A(G1341), .B(n956), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1007 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1008 ( .A1(n917), .A2(n916), .ZN(n946) );
  INV_X1 U1009 ( .A(G16), .ZN(n944) );
  XNOR2_X1 U1010 ( .A(G1341), .B(G19), .ZN(n919) );
  XNOR2_X1 U1011 ( .A(G1981), .B(G6), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1013 ( .A(KEYINPUT124), .B(n920), .ZN(n923) );
  XNOR2_X1 U1014 ( .A(n921), .B(G20), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(n926) );
  XOR2_X1 U1016 ( .A(KEYINPUT59), .B(G1348), .Z(n924) );
  XNOR2_X1 U1017 ( .A(G4), .B(n924), .ZN(n925) );
  NOR2_X1 U1018 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1019 ( .A(n927), .B(KEYINPUT125), .ZN(n928) );
  XNOR2_X1 U1020 ( .A(n928), .B(KEYINPUT60), .ZN(n930) );
  XNOR2_X1 U1021 ( .A(G21), .B(G1966), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1023 ( .A(KEYINPUT126), .B(n931), .ZN(n934) );
  XNOR2_X1 U1024 ( .A(n932), .B(G5), .ZN(n933) );
  NAND2_X1 U1025 ( .A1(n934), .A2(n933), .ZN(n941) );
  XNOR2_X1 U1026 ( .A(G1971), .B(G22), .ZN(n936) );
  XNOR2_X1 U1027 ( .A(G23), .B(G1976), .ZN(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G1986), .B(G24), .Z(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(KEYINPUT58), .B(n939), .ZN(n940) );
  NOR2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(KEYINPUT61), .B(n942), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1035 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1036 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1037 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1038 ( .A(KEYINPUT62), .B(n951), .Z(G311) );
  XNOR2_X1 U1039 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1040 ( .A(G132), .ZN(G219) );
  INV_X1 U1041 ( .A(G82), .ZN(G220) );
  XOR2_X1 U1042 ( .A(KEYINPUT115), .B(n952), .Z(n955) );
  XNOR2_X1 U1043 ( .A(n953), .B(G171), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(n955), .B(n954), .ZN(n958) );
  XOR2_X1 U1045 ( .A(G286), .B(n956), .Z(n957) );
  XNOR2_X1 U1046 ( .A(n958), .B(n957), .ZN(n959) );
  NOR2_X1 U1047 ( .A1(G37), .A2(n959), .ZN(G397) );
  XOR2_X1 U1048 ( .A(G2100), .B(G2096), .Z(n961) );
  XNOR2_X1 U1049 ( .A(G2090), .B(KEYINPUT43), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(n961), .B(n960), .ZN(n962) );
  XOR2_X1 U1051 ( .A(n962), .B(KEYINPUT110), .Z(n964) );
  XNOR2_X1 U1052 ( .A(G2072), .B(G2678), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(n964), .B(n963), .ZN(n968) );
  XOR2_X1 U1054 ( .A(KEYINPUT42), .B(G2084), .Z(n966) );
  XNOR2_X1 U1055 ( .A(G2067), .B(G2078), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(n966), .B(n965), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(n968), .B(n967), .ZN(G227) );
  XOR2_X1 U1058 ( .A(G1976), .B(G1981), .Z(n970) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G1971), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(n970), .B(n969), .ZN(n971) );
  XOR2_X1 U1061 ( .A(n971), .B(KEYINPUT41), .Z(n973) );
  XNOR2_X1 U1062 ( .A(G1996), .B(G1991), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1064 ( .A(G2474), .B(G1986), .Z(n975) );
  XNOR2_X1 U1065 ( .A(G1956), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n975), .B(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n977), .B(n976), .ZN(G229) );
  XNOR2_X1 U1068 ( .A(G160), .B(n978), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n980), .B(n979), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G164), .B(n981), .ZN(n1004) );
  XOR2_X1 U1071 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n983) );
  XNOR2_X1 U1072 ( .A(G162), .B(KEYINPUT46), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n983), .B(n982), .ZN(n998) );
  NAND2_X1 U1074 ( .A1(G130), .A2(n984), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(G118), .A2(n985), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n996) );
  XNOR2_X1 U1077 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n994) );
  NAND2_X1 U1078 ( .A1(n988), .A2(G142), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n989), .A2(G106), .ZN(n990) );
  XOR2_X1 U1080 ( .A(KEYINPUT111), .B(n990), .Z(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1082 ( .A(n994), .B(n993), .Z(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1084 ( .A(n998), .B(n997), .Z(n1002) );
  XNOR2_X1 U1085 ( .A(n1000), .B(n999), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(n1002), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(n1004), .B(n1003), .ZN(n1006) );
  XOR2_X1 U1088 ( .A(n1006), .B(n1005), .Z(n1007) );
  NOR2_X1 U1089 ( .A1(G37), .A2(n1007), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(KEYINPUT114), .B(n1008), .ZN(G395) );
  NOR2_X1 U1091 ( .A1(G401), .A2(n1009), .ZN(n1014) );
  NOR2_X1 U1092 ( .A1(G227), .A2(G229), .ZN(n1011) );
  XNOR2_X1 U1093 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(n1011), .B(n1010), .ZN(n1012) );
  NOR2_X1 U1095 ( .A1(G397), .A2(n1012), .ZN(n1013) );
  NAND2_X1 U1096 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1097 ( .A1(n1015), .A2(G395), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(n1016), .B(KEYINPUT117), .ZN(G225) );
  INV_X1 U1099 ( .A(G225), .ZN(G308) );
  INV_X1 U1100 ( .A(G69), .ZN(G235) );
  INV_X1 U1101 ( .A(G96), .ZN(G221) );
endmodule

