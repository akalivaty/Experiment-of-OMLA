//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(KEYINPUT27), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT27), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G183gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(G183gat), .ZN(new_n210));
  AOI21_X1  g009(.A(G190gat), .B1(new_n210), .B2(KEYINPUT65), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT28), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(KEYINPUT28), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n203), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT28), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n205), .A2(KEYINPUT27), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT65), .B1(new_n210), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT65), .B1(new_n205), .B2(KEYINPUT27), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n214), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT66), .A3(new_n215), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT26), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR3_X1   g027(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n228), .A2(new_n229), .B1(new_n205), .B2(new_n214), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n217), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n234), .A2(new_n225), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n205), .A2(new_n214), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n235), .B(new_n236), .C1(new_n237), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n237), .A2(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n237), .A2(KEYINPUT64), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(new_n238), .A3(new_n239), .A4(new_n244), .ZN(new_n245));
  AND4_X1   g044(.A1(KEYINPUT25), .A2(new_n236), .A3(new_n234), .A4(new_n225), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n241), .A2(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n202), .B1(new_n232), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n252), .ZN(new_n254));
  INV_X1    g053(.A(G197gat), .ZN(new_n255));
  INV_X1    g054(.A(G204gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G197gat), .A2(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT22), .ZN(new_n259));
  NAND2_X1  g058(.A1(G211gat), .A2(G218gat), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n254), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n261), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n252), .A3(new_n251), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n202), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT29), .B1(new_n232), .B2(new_n248), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n250), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G92gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT73), .B(G64gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n274), .A2(KEYINPUT30), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT72), .B1(new_n268), .B2(new_n267), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n223), .A2(new_n215), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n230), .B1(new_n278), .B2(new_n203), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n247), .B1(new_n279), .B2(new_n224), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n277), .B(new_n202), .C1(new_n280), .C2(KEYINPUT29), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n249), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n265), .B(KEYINPUT71), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n269), .B(new_n275), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT75), .B(KEYINPUT30), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n269), .B1(new_n282), .B2(new_n283), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(new_n273), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n269), .B(new_n274), .C1(new_n282), .C2(new_n283), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  OAI22_X1  g091(.A1(new_n286), .A2(new_n287), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G1gat), .B(G29gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT0), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(G57gat), .ZN(new_n296));
  INV_X1    g095(.A(G85gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G113gat), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT1), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G113gat), .A2(G120gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n300), .A2(new_n305), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT80), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G155gat), .ZN(new_n312));
  INV_X1    g111(.A(G162gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n317), .B2(KEYINPUT2), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT76), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G141gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n323), .A3(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n321), .A2(new_n323), .A3(new_n326), .A4(G148gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT78), .B(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G141gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT79), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n324), .A2(KEYINPUT77), .B1(new_n328), .B2(G141gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n327), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n319), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336));
  INV_X1    g135(.A(G148gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT2), .B1(new_n320), .B2(new_n337), .ZN(new_n338));
  AOI211_X1 g137(.A(new_n316), .B(new_n314), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n311), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  AND4_X1   g139(.A1(new_n333), .A2(new_n325), .A3(new_n327), .A4(new_n329), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n333), .B1(new_n332), .B2(new_n327), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n318), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n339), .ZN(new_n344));
  INV_X1    g143(.A(new_n309), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n335), .A2(new_n339), .A3(new_n309), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n343), .A2(new_n356), .A3(new_n344), .A4(new_n345), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n335), .A2(new_n339), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n361), .A2(KEYINPUT82), .A3(new_n356), .A4(new_n345), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n346), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n357), .A2(new_n360), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(new_n335), .B2(new_n339), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n366), .A3(new_n344), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n367), .A3(new_n311), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n368), .A2(new_n348), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n353), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n358), .ZN(new_n372));
  AND4_X1   g171(.A1(new_n348), .A2(new_n372), .A3(new_n368), .A4(new_n351), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n299), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n348), .B1(new_n372), .B2(new_n368), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n340), .A2(new_n346), .A3(new_n348), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT39), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n376), .B2(KEYINPUT39), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n356), .B1(new_n361), .B2(new_n345), .ZN(new_n381));
  INV_X1    g180(.A(new_n358), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n368), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT39), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n349), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n298), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT40), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n299), .B1(new_n375), .B2(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT40), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n349), .ZN(new_n390));
  INV_X1    g189(.A(new_n379), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n388), .B(new_n389), .C1(new_n392), .C2(new_n378), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n293), .A2(new_n374), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(G50gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT85), .ZN(new_n400));
  INV_X1    g199(.A(G22gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n266), .B1(new_n367), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n343), .A2(new_n344), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n366), .B1(new_n265), .B2(KEYINPUT29), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n402), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(KEYINPUT86), .B(new_n402), .C1(new_n404), .C2(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n283), .B1(new_n367), .B2(new_n403), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n413), .A2(new_n407), .A3(new_n402), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n401), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  AOI211_X1 g215(.A(G22gat), .B(new_n414), .C1(new_n410), .C2(new_n411), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n400), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n405), .A2(new_n406), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT29), .B1(new_n361), .B2(new_n366), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(new_n266), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT86), .B1(new_n421), .B2(new_n402), .ZN(new_n422));
  INV_X1    g221(.A(new_n411), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n415), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(G22gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n412), .A2(new_n401), .A3(new_n415), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n399), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n395), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n289), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n274), .B1(new_n430), .B2(KEYINPUT38), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n364), .A2(new_n369), .ZN(new_n432));
  INV_X1    g231(.A(new_n353), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n373), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .A4(new_n299), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n298), .A2(KEYINPUT6), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n299), .A2(new_n436), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n438), .B(new_n439), .C1(new_n370), .C2(new_n373), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n276), .A2(new_n281), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n283), .B1(new_n443), .B2(new_n250), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT37), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n269), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n232), .A2(new_n248), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n403), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n249), .B1(new_n449), .B2(new_n202), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT37), .B1(new_n450), .B2(new_n266), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n451), .B(KEYINPUT88), .C1(new_n283), .C2(new_n282), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n443), .A2(new_n283), .A3(new_n250), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n450), .A2(new_n266), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n274), .B1(new_n456), .B2(KEYINPUT37), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT38), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n289), .B2(KEYINPUT37), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n441), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n429), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n232), .A2(new_n345), .A3(new_n248), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n345), .B1(new_n232), .B2(new_n248), .ZN(new_n467));
  INV_X1    g266(.A(G227gat), .ZN(new_n468));
  INV_X1    g267(.A(G233gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT68), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT34), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n467), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n280), .A2(new_n345), .ZN(new_n475));
  INV_X1    g274(.A(new_n470), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(KEYINPUT68), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n470), .B1(new_n466), .B2(new_n467), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT32), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT33), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G43gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G71gat), .B(G99gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT67), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490));
  AOI211_X1 g289(.A(new_n490), .B(new_n487), .C1(new_n481), .C2(new_n483), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n482), .B1(new_n488), .B2(KEYINPUT33), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n481), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n465), .B(new_n480), .C1(new_n492), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n484), .A2(new_n488), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n490), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n484), .A2(KEYINPUT67), .A3(new_n488), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n465), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n473), .A2(new_n479), .A3(KEYINPUT69), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n494), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n503), .A3(KEYINPUT36), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n496), .A2(new_n503), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n437), .A2(new_n440), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(new_n293), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n504), .B(new_n507), .C1(new_n509), .C2(new_n428), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n464), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n425), .A2(new_n426), .A3(new_n399), .ZN(new_n513));
  INV_X1    g312(.A(new_n400), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n425), .B2(new_n426), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n505), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n293), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n437), .A2(new_n440), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n512), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n509), .A2(KEYINPUT35), .A3(new_n428), .A4(new_n505), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT89), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n458), .A2(new_n459), .B1(new_n453), .B2(new_n461), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n395), .B(new_n428), .C1(new_n524), .C2(new_n441), .ZN(new_n525));
  INV_X1    g324(.A(new_n428), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n519), .ZN(new_n527));
  INV_X1    g326(.A(new_n504), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT36), .B1(new_n496), .B2(new_n503), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT89), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n520), .A4(new_n521), .ZN(new_n533));
  INV_X1    g332(.A(G8gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(G1gat), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n536), .A2(KEYINPUT94), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n538));
  INV_X1    g337(.A(G1gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT16), .B1(KEYINPUT92), .B2(G1gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT93), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n536), .A2(KEYINPUT94), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n537), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n547), .B2(KEYINPUT93), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n534), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT14), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G29gat), .A2(G36gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G50gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(G43gat), .ZN(new_n556));
  INV_X1    g355(.A(G43gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(G50gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT15), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n553), .B(KEYINPUT91), .Z(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n552), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n558), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT15), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n561), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n536), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n570), .A2(new_n546), .A3(new_n534), .A4(new_n542), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n549), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n569), .B1(new_n549), .B2(new_n572), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(KEYINPUT98), .B(new_n569), .C1(new_n549), .C2(new_n572), .ZN(new_n577));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT97), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT13), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT99), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n576), .A2(KEYINPUT99), .A3(new_n577), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n569), .B(KEYINPUT17), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n549), .A2(new_n572), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT18), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT96), .ZN(new_n590));
  AND4_X1   g389(.A1(new_n575), .A2(new_n588), .A3(new_n578), .A4(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(KEYINPUT96), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n588), .A2(new_n575), .A3(new_n578), .A4(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT11), .ZN(new_n598));
  INV_X1    g397(.A(G169gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G197gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n595), .A3(new_n602), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n596), .A2(KEYINPUT100), .A3(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT21), .ZN(new_n611));
  XNOR2_X1  g410(.A(G57gat), .B(G64gat), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G71gat), .B(G78gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n587), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n617), .A2(KEYINPUT101), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(KEYINPUT101), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n611), .ZN(new_n620));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n618), .B2(new_n619), .ZN(new_n625));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT102), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n627), .B(new_n630), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n624), .A2(new_n625), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n619), .ZN(new_n634));
  INV_X1    g433(.A(new_n622), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(new_n636), .B2(new_n623), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT105), .B(KEYINPUT7), .ZN(new_n639));
  NAND2_X1  g438(.A1(G85gat), .A2(G92gat), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  INV_X1    g442(.A(G92gat), .ZN(new_n644));
  AOI22_X1  g443(.A1(KEYINPUT8), .A2(new_n643), .B1(new_n297), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G99gat), .B(G106gat), .Z(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n586), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  AND2_X1   g451(.A1(G232gat), .A2(G233gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n652), .A2(new_n569), .B1(KEYINPUT41), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n655), .A2(new_n659), .A3(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G134gat), .B(G162gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT103), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n653), .A2(KEYINPUT41), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT104), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n657), .A2(new_n666), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n658), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n638), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(G230gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n469), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n650), .B(new_n616), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(KEYINPUT10), .ZN(new_n677));
  INV_X1    g476(.A(new_n616), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n652), .A2(KEYINPUT10), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n675), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(G120gat), .B(G148gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G176gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n256), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n683), .B(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n523), .A2(new_n533), .A3(new_n610), .A4(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n518), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(new_n539), .ZN(G1324gat));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n293), .B1(new_n694), .B2(new_n695), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT108), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT16), .B(G8gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n700), .A2(new_n699), .A3(new_n702), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n701), .B2(G8gat), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1325gat));
  OAI21_X1  g505(.A(G15gat), .B1(new_n696), .B2(new_n530), .ZN(new_n707));
  INV_X1    g506(.A(new_n505), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(G15gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n696), .B2(new_n709), .ZN(G1326gat));
  NOR2_X1   g509(.A1(new_n696), .A2(new_n428), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  AND2_X1   g512(.A1(new_n523), .A2(new_n533), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n633), .A2(new_n637), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n688), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n672), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n714), .A2(new_n610), .A3(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(G29gat), .A3(new_n518), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT45), .Z(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n464), .B2(new_n510), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n525), .A2(new_n527), .A3(new_n530), .A4(KEYINPUT109), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n522), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n723), .B1(new_n727), .B2(new_n718), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n718), .A2(new_n723), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n523), .A2(new_n533), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n717), .A2(new_n609), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n518), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n722), .A2(new_n734), .ZN(G1328gat));
  OAI21_X1  g534(.A(G36gat), .B1(new_n733), .B2(new_n517), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n517), .A2(G36gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT46), .B1(new_n720), .B2(new_n738), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n720), .A2(KEYINPUT46), .A3(new_n738), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT110), .Z(G1329gat));
  OAI21_X1  g541(.A(G43gat), .B1(new_n733), .B2(new_n530), .ZN(new_n743));
  INV_X1    g542(.A(new_n720), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n557), .A3(new_n505), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT47), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n746), .B(new_n748), .ZN(G1330gat));
  NAND2_X1  g548(.A1(new_n526), .A2(new_n555), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT112), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT48), .B1(new_n720), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n728), .A2(new_n526), .A3(new_n730), .A4(new_n732), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n754), .A2(KEYINPUT113), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n555), .B1(new_n754), .B2(KEYINPUT113), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(KEYINPUT114), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(KEYINPUT114), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n744), .A2(new_n751), .B1(new_n754), .B2(G50gat), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n758), .A2(new_n759), .B1(KEYINPUT48), .B2(new_n760), .ZN(G1331gat));
  NAND3_X1  g560(.A1(new_n673), .A2(new_n609), .A3(new_n688), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n727), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n508), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g564(.A1(new_n727), .A2(new_n517), .A3(new_n762), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  AND2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n766), .B2(new_n767), .ZN(G1333gat));
  INV_X1    g569(.A(new_n530), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n763), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n708), .A2(G71gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(G71gat), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n763), .A2(new_n526), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g576(.A(KEYINPUT115), .B1(new_n609), .B2(new_n638), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n779), .B(new_n715), .C1(new_n607), .C2(new_n608), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n689), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n725), .A2(new_n726), .ZN(new_n783));
  INV_X1    g582(.A(new_n522), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n718), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n730), .B(new_n782), .C1(new_n785), .C2(KEYINPUT44), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n728), .A2(KEYINPUT116), .A3(new_n730), .A4(new_n782), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n518), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  INV_X1    g591(.A(new_n781), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n718), .A4(new_n781), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n689), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n297), .A3(new_n508), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n791), .A2(new_n797), .ZN(G1336gat));
  NOR2_X1   g597(.A1(new_n517), .A2(G92gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  OAI21_X1  g600(.A(G92gat), .B1(new_n786), .B2(new_n517), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n800), .A2(KEYINPUT118), .A3(new_n801), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n293), .A3(new_n789), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G92gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n800), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(KEYINPUT52), .ZN(new_n812));
  INV_X1    g611(.A(new_n799), .ZN(new_n813));
  NOR4_X1   g612(.A1(new_n794), .A2(new_n795), .A3(new_n689), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n809), .B2(G92gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(KEYINPUT117), .A3(new_n801), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n807), .B1(new_n812), .B2(new_n816), .ZN(G1337gat));
  INV_X1    g616(.A(G99gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n790), .A2(new_n818), .A3(new_n530), .ZN(new_n819));
  AOI21_X1  g618(.A(G99gat), .B1(new_n796), .B2(new_n505), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(G1338gat));
  INV_X1    g620(.A(G106gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n796), .A2(new_n822), .A3(new_n526), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824));
  OAI21_X1  g623(.A(G106gat), .B1(new_n786), .B2(new_n428), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G106gat), .B1(new_n790), .B2(new_n428), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n823), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n828), .B2(new_n824), .ZN(G1339gat));
  NAND3_X1  g628(.A1(new_n677), .A2(new_n679), .A3(new_n675), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n681), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n686), .B1(new_n680), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT55), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n683), .A2(new_n687), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n607), .A3(new_n608), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n580), .B1(new_n576), .B2(new_n577), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n578), .B1(new_n588), .B2(new_n575), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n601), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n606), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n688), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n672), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  AND4_X1   g643(.A1(new_n672), .A2(new_n836), .A3(new_n837), .A4(new_n842), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n638), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n691), .A2(new_n609), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n293), .A2(new_n518), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n516), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT119), .Z(new_n853));
  NOR2_X1   g652(.A1(new_n609), .A2(G113gat), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT120), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n852), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n609), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1340gat));
  NAND3_X1  g658(.A1(new_n853), .A2(new_n303), .A3(new_n688), .ZN(new_n860));
  OAI21_X1  g659(.A(G120gat), .B1(new_n857), .B2(new_n689), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1341gat));
  NAND2_X1  g661(.A1(new_n852), .A2(new_n715), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g663(.A1(new_n852), .A2(new_n672), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT56), .B1(new_n865), .B2(G134gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(G134gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n771), .A2(new_n850), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n848), .A2(new_n526), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n320), .A3(new_n610), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n848), .A2(new_n526), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n870), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n609), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n321), .A2(new_n323), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n872), .A2(new_n328), .A3(new_n688), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n689), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(KEYINPUT59), .A3(new_n328), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n847), .A2(KEYINPUT121), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n691), .B2(new_n609), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n846), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT122), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n892), .B(new_n846), .C1(new_n887), .C2(new_n889), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n428), .A2(KEYINPUT57), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n875), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n688), .A3(new_n870), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n886), .B1(new_n897), .B2(G148gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n882), .B1(new_n885), .B2(new_n898), .ZN(G1345gat));
  OAI21_X1  g698(.A(G155gat), .B1(new_n883), .B2(new_n638), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n872), .A2(new_n312), .A3(new_n715), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n883), .B2(new_n718), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n872), .A2(new_n313), .A3(new_n672), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1347gat));
  NAND3_X1  g704(.A1(new_n505), .A2(new_n518), .A3(new_n293), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT123), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n526), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n848), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n599), .A3(new_n609), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n508), .B1(new_n846), .B2(new_n847), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n516), .A2(new_n517), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n610), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n910), .B1(new_n915), .B2(new_n599), .ZN(G1348gat));
  OAI21_X1  g715(.A(G176gat), .B1(new_n909), .B2(new_n689), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n689), .A2(G176gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n913), .B2(new_n918), .ZN(G1349gat));
  OAI21_X1  g718(.A(G183gat), .B1(new_n909), .B2(new_n638), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n715), .A2(new_n213), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n913), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n214), .A3(new_n672), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n848), .A2(new_n672), .A3(new_n908), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n925), .A2(new_n926), .A3(G190gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n925), .B2(G190gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT124), .Z(G1351gat));
  NOR3_X1   g729(.A1(new_n771), .A2(new_n517), .A3(new_n428), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n610), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n771), .A2(new_n508), .A3(new_n517), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n896), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n609), .A2(new_n255), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1352gat));
  NOR3_X1   g737(.A1(new_n932), .A2(G204gat), .A3(new_n689), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(KEYINPUT125), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n896), .A2(new_n688), .A3(new_n935), .ZN(new_n943));
  OAI221_X1 g742(.A(new_n941), .B1(new_n939), .B2(new_n942), .C1(new_n943), .C2(new_n256), .ZN(G1353gat));
  NAND4_X1  g743(.A1(new_n895), .A2(new_n715), .A3(new_n875), .A4(new_n935), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n932), .A2(G211gat), .A3(new_n638), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT126), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n952), .B1(new_n946), .B2(new_n947), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(G1354gat));
  AOI21_X1  g753(.A(G218gat), .B1(new_n933), .B2(new_n672), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n672), .A2(G218gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n936), .B2(new_n956), .ZN(G1355gat));
endmodule


