//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT64), .B1(new_n193), .B2(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(G146), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n197));
  OAI21_X1  g011(.A(G128), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n196), .A2(new_n198), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT10), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n205), .C2(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT79), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT80), .B(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G104), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT81), .B(G101), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G104), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n210), .A2(new_n217), .A3(new_n218), .A4(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n216), .A2(G104), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n205), .A2(G107), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n222), .A2(KEYINPUT82), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT82), .B1(new_n222), .B2(new_n225), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n204), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n208), .A2(new_n209), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n219), .A2(KEYINPUT80), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n232), .A3(G104), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n221), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(G101), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n196), .A2(new_n240), .B1(new_n199), .B2(new_n238), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n242), .B(G101), .C1(new_n229), .C2(new_n235), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n237), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  MUX2_X1   g058(.A(new_n198), .B(new_n201), .S(new_n199), .Z(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n222), .A3(new_n225), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n203), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n248), .A2(new_n249), .B1(G134), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(G134), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G137), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(G131), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n254), .A2(G137), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n250), .A2(G134), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n248), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  INV_X1    g075(.A(new_n249), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n253), .B1(new_n262), .B2(new_n252), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n228), .A2(new_n244), .A3(new_n247), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT84), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n243), .A2(new_n241), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n271), .A2(new_n237), .B1(new_n203), .B2(new_n246), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n272), .A2(KEYINPUT84), .A3(new_n228), .A4(new_n267), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(G227), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n265), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n272), .B2(new_n228), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n270), .A2(new_n273), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n222), .A2(new_n225), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n222), .A2(KEYINPUT82), .A3(new_n225), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n202), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n246), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT12), .B1(new_n291), .B2(new_n265), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT12), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n293), .B(new_n281), .C1(new_n290), .C2(new_n246), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n284), .B1(new_n285), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n196), .A2(new_n198), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n199), .A2(new_n201), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n226), .A2(new_n227), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n246), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n265), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n293), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n291), .A2(KEYINPUT12), .A3(new_n265), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n274), .A3(KEYINPUT85), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n283), .B1(new_n307), .B2(new_n278), .ZN(new_n308));
  OAI21_X1  g122(.A(G469), .B1(new_n308), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT86), .B(G469), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n305), .A2(new_n279), .A3(new_n274), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n282), .B1(new_n270), .B2(new_n273), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(new_n279), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT87), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI22_X1  g131(.A1(new_n280), .A2(new_n295), .B1(new_n313), .B2(new_n279), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(KEYINPUT87), .A3(new_n310), .A4(new_n311), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n189), .B1(new_n309), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(KEYINPUT73), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(G125), .A3(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n323), .B2(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G146), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n191), .B1(new_n327), .B2(new_n329), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G128), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n334), .A2(G128), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G110), .ZN(new_n339));
  XNOR2_X1  g153(.A(G119), .B(G128), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT72), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT24), .B(G110), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT74), .B1(new_n333), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n330), .B(G146), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n340), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n342), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n345), .A2(new_n346), .A3(new_n350), .A4(new_n339), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G137), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n355), .B2(new_n359), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G125), .B(G140), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n332), .B1(new_n191), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n348), .A2(new_n349), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n338), .A2(G110), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n352), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n363), .B1(new_n352), .B2(new_n368), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n310), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n352), .A2(new_n368), .ZN(new_n374));
  INV_X1    g188(.A(new_n363), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n352), .A2(new_n363), .A3(new_n368), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT25), .A3(new_n310), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G217), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(G234), .B2(new_n310), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(G902), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT77), .B1(new_n376), .B2(new_n377), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT67), .ZN(new_n390));
  OAI21_X1  g204(.A(G131), .B1(new_n258), .B2(new_n259), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n299), .A2(new_n264), .A3(new_n391), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n251), .A2(new_n256), .A3(G131), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n261), .B1(new_n260), .B2(new_n263), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n241), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT66), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n265), .A2(KEYINPUT66), .A3(new_n241), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n392), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n390), .B1(new_n399), .B2(KEYINPUT30), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n299), .A2(new_n264), .A3(new_n391), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n265), .A2(KEYINPUT66), .A3(new_n241), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT66), .B1(new_n265), .B2(new_n241), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(KEYINPUT67), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G116), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT68), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT68), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G116), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n410), .A3(G119), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n334), .A2(G116), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT2), .B(G113), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n414), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n411), .A3(new_n412), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n401), .A2(new_n395), .A3(KEYINPUT30), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n400), .A2(new_n406), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n401), .A2(new_n395), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n418), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n423));
  NOR2_X1   g237(.A1(G237), .A2(G953), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G210), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n423), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT26), .B(G101), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n422), .A2(KEYINPUT70), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n420), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT31), .ZN(new_n431));
  INV_X1    g245(.A(new_n428), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT28), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n422), .B(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n404), .A2(new_n418), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT31), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n420), .A2(new_n438), .A3(new_n429), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G472), .A2(G902), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT32), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT32), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n421), .A2(new_n418), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n434), .A2(KEYINPUT29), .A3(new_n432), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n310), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n434), .A2(new_n435), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n432), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n422), .A2(new_n432), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n420), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G472), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n389), .B1(new_n446), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n460), .B(KEYINPUT89), .Z(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n411), .A2(KEYINPUT5), .A3(new_n412), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n412), .A2(KEYINPUT5), .ZN(new_n464));
  INV_X1    g278(.A(G113), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT88), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n463), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n470), .A3(new_n417), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n288), .B2(new_n289), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n473));
  INV_X1    g287(.A(G101), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n230), .A2(new_n232), .A3(G104), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n220), .B1(new_n475), .B2(new_n215), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n476), .B2(new_n210), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n243), .A2(new_n418), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n462), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n468), .A2(new_n470), .A3(new_n417), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n227), .B2(new_n226), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n243), .A2(new_n418), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n237), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n461), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(KEYINPUT6), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n488), .B(new_n462), .C1(new_n472), .C2(new_n480), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n299), .A2(G125), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n241), .A2(new_n323), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n276), .A2(G224), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT90), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n489), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n202), .A2(new_n323), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT7), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n498), .B2(new_n493), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n497), .B(new_n500), .C1(new_n323), .C2(new_n241), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT91), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n493), .A2(KEYINPUT7), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n503), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n501), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n288), .A2(new_n289), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n507), .A2(new_n482), .B1(new_n237), .B2(new_n484), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n508), .B2(new_n461), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n461), .B(KEYINPUT8), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n467), .A2(new_n417), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n288), .B2(new_n289), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n471), .A2(new_n286), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(G902), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G210), .B1(G237), .B2(G902), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n496), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n496), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n459), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G237), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n276), .A3(G214), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(new_n193), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G131), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n521), .A2(new_n193), .ZN(new_n524));
  AOI21_X1  g338(.A(G143), .B1(new_n424), .B2(G214), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n261), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(KEYINPUT17), .A3(G131), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n333), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G113), .B(G122), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(new_n205), .ZN(new_n533));
  AND2_X1   g347(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G131), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n364), .A2(new_n191), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n324), .A2(G146), .A3(new_n326), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n526), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT94), .ZN(new_n539));
  OAI211_X1 g353(.A(G131), .B(new_n534), .C1(new_n524), .C2(new_n525), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n531), .B(new_n533), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT19), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n364), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n324), .A2(KEYINPUT19), .A3(new_n326), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT95), .B1(new_n549), .B2(G146), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n547), .A2(new_n548), .A3(new_n551), .A4(new_n191), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n332), .B1(new_n523), .B2(new_n527), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n542), .B2(new_n543), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n533), .B1(new_n556), .B2(KEYINPUT96), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n526), .A2(new_n535), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n536), .A2(new_n537), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n540), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT94), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n561), .A2(new_n541), .B1(new_n553), .B2(new_n554), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n545), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G475), .A2(G902), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT20), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n533), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n562), .B2(new_n563), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n556), .A2(KEYINPUT96), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n544), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(new_n566), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n561), .A2(new_n541), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n533), .B1(new_n575), .B2(new_n531), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n310), .B1(new_n545), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n568), .A2(new_n574), .B1(G475), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n408), .A2(new_n410), .A3(G122), .ZN(new_n579));
  INV_X1    g393(.A(G122), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G116), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n582), .A2(KEYINPUT97), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(KEYINPUT97), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n216), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n216), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n193), .A2(G128), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n200), .A2(G143), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n254), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n592), .B(KEYINPUT99), .Z(new_n593));
  NAND3_X1  g407(.A1(new_n193), .A2(KEYINPUT13), .A3(G128), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n591), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT13), .B1(new_n193), .B2(G128), .ZN(new_n596));
  OAI21_X1  g410(.A(G134), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n597), .A2(KEYINPUT98), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(KEYINPUT98), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n593), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n589), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n582), .A2(KEYINPUT14), .ZN(new_n603));
  INV_X1    g417(.A(new_n579), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n219), .B1(new_n604), .B2(KEYINPUT14), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n590), .A2(new_n591), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G134), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n603), .A2(new_n605), .B1(new_n592), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n588), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n187), .A2(new_n381), .A3(G953), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n602), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n610), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n600), .B1(new_n587), .B2(new_n588), .ZN(new_n613));
  INV_X1    g427(.A(new_n609), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G478), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(KEYINPUT15), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(KEYINPUT15), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  AOI211_X1 g438(.A(G902), .B(new_n622), .C1(new_n611), .C2(new_n615), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n578), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(G234), .A2(G237), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(G952), .A3(new_n276), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(G902), .A3(G953), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT21), .B(G898), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n519), .A2(new_n627), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n321), .A2(new_n458), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(new_n218), .Z(G3));
  INV_X1    g451(.A(new_n442), .ZN(new_n638));
  INV_X1    g452(.A(G472), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n440), .B2(new_n310), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n638), .A2(new_n640), .A3(new_n389), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n321), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT101), .Z(new_n643));
  INV_X1    g457(.A(new_n578), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n611), .A2(new_n615), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT33), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n611), .A2(new_n615), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(G478), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n617), .A2(new_n310), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n616), .B2(new_n617), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n519), .A3(new_n634), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n643), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  INV_X1    g471(.A(new_n626), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n578), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n659), .A2(new_n519), .A3(new_n634), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n643), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NAND2_X1  g477(.A1(new_n309), .A2(new_n320), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n188), .A3(new_n635), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n420), .A2(new_n438), .A3(new_n429), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n438), .B1(new_n420), .B2(new_n429), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n666), .A2(new_n667), .A3(new_n436), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n668), .B2(G902), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(new_n374), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n384), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n383), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n442), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n669), .A2(new_n673), .A3(KEYINPUT102), .A4(new_n442), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n665), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT37), .B(G110), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  NAND2_X1  g495(.A1(new_n446), .A2(new_n457), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n321), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n684));
  OR3_X1    g498(.A1(new_n631), .A2(new_n684), .A3(G900), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n684), .B1(new_n631), .B2(G900), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n629), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n659), .A2(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n380), .A2(new_n382), .B1(new_n384), .B2(new_n671), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n519), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  OR2_X1    g508(.A1(new_n421), .A2(new_n418), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n428), .B1(new_n420), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(G902), .B1(new_n454), .B2(new_n447), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n446), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n517), .A2(new_n518), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT105), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n701), .B(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n644), .A2(new_n658), .ZN(new_n706));
  INV_X1    g520(.A(new_n459), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n706), .A2(new_n673), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n700), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n687), .B(KEYINPUT39), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n321), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n709), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n193), .ZN(G45));
  NAND2_X1  g531(.A1(new_n649), .A2(new_n651), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n578), .A2(new_n718), .A3(new_n688), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n691), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n683), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  NAND2_X1  g536(.A1(new_n458), .A2(new_n654), .ZN(new_n723));
  INV_X1    g537(.A(G469), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n318), .B2(new_n310), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n189), .B(new_n725), .C1(new_n317), .C2(new_n319), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT41), .B(G113), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND2_X1  g544(.A1(new_n458), .A2(new_n660), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n727), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n407), .ZN(G18));
  NOR2_X1   g547(.A1(new_n627), .A2(new_n634), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n682), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n725), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n320), .A2(new_n188), .A3(new_n691), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n334), .ZN(G21));
  OR2_X1    g553(.A1(new_n517), .A2(new_n518), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n459), .A3(new_n658), .A4(new_n644), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n634), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n726), .ZN(new_n743));
  INV_X1    g557(.A(new_n389), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n434), .A2(new_n447), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n428), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n431), .A2(new_n439), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n747), .A2(new_n748), .A3(new_n441), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n747), .B2(new_n441), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n744), .B(new_n669), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n580), .ZN(G24));
  OAI211_X1 g567(.A(new_n719), .B(new_n669), .C1(new_n749), .C2(new_n750), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n726), .A3(new_n756), .A4(new_n691), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT107), .B1(new_n737), .B2(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n701), .A2(new_n188), .A3(new_n459), .ZN(new_n762));
  NAND2_X1  g576(.A1(G469), .A2(G902), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT108), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n308), .B2(G469), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n762), .B1(new_n765), .B2(new_n320), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n719), .ZN(new_n767));
  INV_X1    g581(.A(new_n458), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n761), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n458), .A3(KEYINPUT42), .A4(new_n719), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n458), .A3(new_n689), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  NAND2_X1  g588(.A1(new_n701), .A2(new_n459), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n652), .A2(new_n578), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n669), .A2(new_n442), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n673), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n775), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n779), .A4(new_n673), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT109), .ZN(new_n785));
  INV_X1    g599(.A(new_n320), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n305), .A2(KEYINPUT85), .A3(new_n274), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT85), .B1(new_n305), .B2(new_n274), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n278), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n283), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n724), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  INV_X1    g608(.A(new_n764), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n786), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n188), .A3(new_n710), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n785), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  NAND2_X1  g617(.A1(new_n719), .A2(new_n389), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n682), .A2(new_n775), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT47), .B1(new_n800), .B2(new_n188), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n807), .B(new_n189), .C1(new_n798), .C2(new_n799), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NOR2_X1   g624(.A1(new_n775), .A2(new_n629), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n726), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n700), .A2(new_n389), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(KEYINPUT115), .A3(new_n813), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n578), .A3(new_n718), .A4(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n669), .B(new_n673), .C1(new_n749), .C2(new_n750), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n778), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n751), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n630), .A3(new_n778), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n704), .A2(new_n707), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n727), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(KEYINPUT50), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n823), .A2(new_n827), .A3(new_n727), .A4(new_n824), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n818), .B(new_n821), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n800), .A2(new_n188), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n807), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n800), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n786), .A2(new_n725), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n189), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n823), .A2(new_n775), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n831), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n812), .A2(new_n458), .A3(new_n778), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT48), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n816), .A2(new_n644), .A3(new_n652), .A4(new_n817), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n823), .A2(new_n727), .A3(new_n519), .ZN(new_n846));
  INV_X1    g660(.A(G952), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n846), .A2(new_n847), .A3(G953), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n837), .A2(new_n840), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n826), .A2(new_n828), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n818), .A4(new_n821), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n854));
  AOI22_X1  g668(.A1(KEYINPUT114), .A2(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n850), .A2(KEYINPUT114), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n842), .B(new_n849), .C1(new_n857), .C2(KEYINPUT51), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n321), .B(new_n682), .C1(new_n692), .C2(new_n720), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n741), .B1(new_n446), .B2(new_n699), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n690), .A2(new_n188), .A3(new_n687), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n765), .B2(new_n320), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g679(.A(KEYINPUT112), .B(new_n862), .C1(new_n765), .C2(new_n320), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n757), .A2(new_n758), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n859), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n765), .A2(new_n320), .ZN(new_n870));
  INV_X1    g684(.A(new_n862), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT112), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n863), .A2(new_n864), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n861), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n759), .A3(KEYINPUT52), .A4(new_n860), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT113), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n869), .A2(KEYINPUT113), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n773), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n769), .B2(new_n770), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n727), .B1(new_n723), .B2(new_n731), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n743), .A2(new_n751), .B1(new_n735), .B2(new_n737), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n767), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n775), .A2(new_n627), .A3(new_n690), .A4(new_n688), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n887), .A2(new_n820), .B1(new_n683), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n883), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n321), .A2(new_n654), .A3(new_n641), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n636), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT110), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n664), .A2(new_n188), .A3(new_n641), .A4(new_n660), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n665), .B2(new_n678), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n895), .B(KEYINPUT110), .C1(new_n665), .C2(new_n678), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT111), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n896), .A2(new_n894), .ZN(new_n900));
  INV_X1    g714(.A(new_n893), .ZN(new_n901));
  AND4_X1   g715(.A1(KEYINPUT111), .A2(new_n900), .A3(new_n898), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n891), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT53), .B1(new_n881), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n900), .A2(new_n901), .A3(new_n898), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n897), .A2(KEYINPUT111), .A3(new_n898), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n890), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n877), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n904), .A2(KEYINPUT54), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n910), .B1(new_n881), .B2(new_n903), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n877), .A2(KEYINPUT53), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT54), .B1(new_n915), .B2(new_n909), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n858), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n835), .B(KEYINPUT49), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n744), .A2(new_n188), .A3(new_n459), .ZN(new_n921));
  NOR4_X1   g735(.A1(new_n705), .A2(new_n700), .A3(new_n776), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n919), .A2(new_n923), .ZN(G75));
  NAND2_X1  g738(.A1(new_n847), .A2(G953), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT120), .Z(new_n926));
  NAND2_X1  g740(.A1(new_n915), .A2(new_n909), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n310), .B1(new_n913), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(G210), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n487), .A2(new_n489), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT118), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n495), .B(KEYINPUT55), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n926), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n913), .A2(new_n927), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(G902), .ZN(new_n937));
  INV_X1    g751(.A(G210), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n935), .B(new_n933), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n929), .A2(KEYINPUT119), .A3(new_n933), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n934), .B1(new_n941), .B2(new_n942), .ZN(G51));
  INV_X1    g757(.A(new_n926), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n869), .A2(KEYINPUT113), .A3(new_n876), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT113), .B1(new_n869), .B2(new_n876), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT53), .B1(new_n947), .B2(new_n909), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n903), .A2(new_n914), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT54), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT54), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n903), .B2(new_n914), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n913), .A2(KEYINPUT121), .A3(new_n916), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n764), .B(KEYINPUT57), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n318), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n937), .A2(new_n794), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n944), .B1(new_n959), .B2(new_n960), .ZN(G54));
  INV_X1    g775(.A(KEYINPUT122), .ZN(new_n962));
  AND2_X1   g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n928), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n964), .B2(new_n565), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n944), .B1(new_n964), .B2(new_n565), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n928), .A2(KEYINPUT122), .A3(new_n572), .A4(new_n963), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(G60));
  XNOR2_X1  g782(.A(new_n650), .B(KEYINPUT59), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n912), .B2(new_n917), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n646), .A2(new_n648), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n926), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n646), .B2(new_n648), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n956), .B2(new_n973), .ZN(G63));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT61), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n386), .A2(new_n387), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n948), .A2(new_n949), .ZN(new_n979));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT60), .Z(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n978), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n936), .A2(new_n671), .A3(new_n981), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n926), .B1(new_n975), .B2(KEYINPUT61), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n976), .A2(new_n983), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n936), .A2(new_n981), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n985), .B1(new_n988), .B2(new_n978), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n976), .B1(new_n989), .B2(new_n984), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n987), .A2(new_n990), .ZN(G66));
  OAI21_X1  g805(.A(new_n886), .B1(new_n899), .B2(new_n902), .ZN(new_n992));
  NAND2_X1  g806(.A1(G224), .A2(G953), .ZN(new_n993));
  OAI22_X1  g807(.A1(new_n992), .A2(G953), .B1(new_n633), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n931), .B1(G898), .B2(new_n276), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n994), .B(new_n995), .Z(G69));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n400), .A2(new_n406), .A3(new_n419), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n549), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(G900), .B2(G953), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n768), .A2(new_n741), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n800), .A2(new_n188), .A3(new_n710), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT125), .Z(new_n1004));
  NAND3_X1  g818(.A1(new_n883), .A2(new_n759), .A3(new_n860), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n785), .B2(new_n801), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1004), .A2(new_n809), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1001), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n653), .A2(new_n659), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT124), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n775), .B1(new_n1009), .B2(KEYINPUT124), .ZN(new_n1011));
  AND4_X1   g825(.A1(new_n458), .A2(new_n712), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n785), .B2(new_n801), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n759), .A2(new_n860), .ZN(new_n1014));
  OAI21_X1  g828(.A(KEYINPUT62), .B1(new_n716), .B2(new_n1014), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n716), .A2(KEYINPUT62), .A3(new_n1014), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1013), .A2(new_n809), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n276), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n1000), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n997), .B1(new_n1008), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1008), .A2(new_n1019), .A3(new_n997), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1023), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1022), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n1026), .B2(new_n1020), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1024), .A2(new_n1027), .ZN(G72));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  OAI21_X1  g844(.A(new_n1030), .B1(new_n1007), .B2(new_n992), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1031), .A2(new_n420), .A3(new_n454), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1030), .B1(new_n1017), .B2(new_n992), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n696), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1032), .A2(new_n1034), .A3(new_n926), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n455), .A2(new_n1030), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1036), .A2(new_n696), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n904), .A2(new_n911), .A3(new_n1037), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n1038), .A2(KEYINPUT127), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(KEYINPUT127), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(G57));
endmodule


