//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n561, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g030(.A1(G113), .A2(G2104), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n459), .A2(G2105), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n463), .A2(G2105), .B1(G101), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n457), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n460), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT68), .ZN(G160));
  NAND4_X1  g048(.A1(new_n468), .A2(new_n469), .A3(G2105), .A4(new_n460), .ZN(new_n474));
  INV_X1    g049(.A(G124), .ZN(new_n475));
  AND2_X1   g050(.A1(G112), .A2(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n476), .B1(G100), .B2(new_n470), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n474), .A2(new_n475), .B1(new_n477), .B2(new_n459), .ZN(new_n478));
  INV_X1    g053(.A(new_n471), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G136), .ZN(G162));
  AND3_X1   g055(.A1(new_n468), .A2(new_n469), .A3(new_n460), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G138), .A4(new_n470), .ZN(new_n483));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT70), .B1(new_n471), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(KEYINPUT4), .A3(new_n485), .ZN(new_n486));
  NOR4_X1   g061(.A1(new_n461), .A2(KEYINPUT4), .A3(new_n484), .A4(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT67), .B1(new_n457), .B2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n457), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n492), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G102), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT69), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI211_X1 g074(.A(KEYINPUT69), .B(new_n497), .C1(new_n474), .C2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n489), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(new_n509), .B1(new_n506), .B2(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(new_n514), .A3(new_n511), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(new_n510), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n511), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(G651), .B1(G50), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n522), .A2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n511), .A2(new_n528), .A3(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(G51), .B1(new_n510), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n513), .A2(G89), .A3(new_n515), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n533), .A2(KEYINPUT74), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT74), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g115(.A(KEYINPUT75), .B(new_n532), .C1(new_n536), .C2(new_n537), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(G168));
  NAND2_X1  g117(.A1(new_n516), .A2(G90), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n530), .A2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  AOI22_X1  g124(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(G651), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n516), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n530), .A2(G43), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT77), .Z(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  XOR2_X1   g135(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G188));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n522), .A2(KEYINPUT9), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n522), .B2(new_n565), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n519), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n516), .A2(G91), .B1(G651), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G299));
  AND2_X1   g151(.A1(new_n540), .A2(new_n541), .ZN(G286));
  NAND2_X1  g152(.A1(new_n516), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n523), .A2(G49), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n516), .A2(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n519), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G48), .B2(new_n523), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n530), .A2(G47), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n513), .A2(new_n515), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n592), .A2(KEYINPUT81), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(KEYINPUT81), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n593), .A2(new_n594), .B1(new_n545), .B2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n516), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n590), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n519), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(new_n530), .B2(G54), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT82), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G168), .B2(new_n611), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(G168), .B2(new_n611), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND3_X1  g191(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n608), .A2(new_n615), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n617), .B(new_n618), .S(G868), .Z(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g195(.A(new_n464), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n461), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n479), .A2(G135), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  AND2_X1   g202(.A1(G111), .A2(G2105), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G99), .B2(new_n470), .ZN(new_n629));
  OAI22_X1  g204(.A1(new_n474), .A2(new_n627), .B1(new_n629), .B2(new_n459), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(G2096), .B1(new_n626), .B2(new_n630), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n625), .A2(new_n633), .A3(new_n634), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2427), .ZN(new_n639));
  INV_X1    g214(.A(G2430), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n642), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  INV_X1    g235(.A(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n657), .B1(new_n663), .B2(new_n654), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n655), .B2(new_n662), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n655), .A2(new_n658), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n661), .B1(new_n666), .B2(KEYINPUT17), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n660), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n632), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(G2100), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(G2100), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n674), .A2(new_n679), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n679), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n682));
  AOI211_X1 g257(.A(new_n678), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n681), .B2(new_n682), .ZN(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT85), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT86), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT89), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G305), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  NAND2_X1  g280(.A1(G166), .A2(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G16), .B2(G22), .ZN(new_n707));
  INV_X1    g282(.A(G1971), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NOR4_X1   g285(.A1(new_n700), .A2(new_n705), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(G16), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT88), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1986), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n479), .A2(G131), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT87), .ZN(new_n719));
  INV_X1    g294(.A(new_n474), .ZN(new_n720));
  MUX2_X1   g295(.A(G95), .B(G107), .S(G2105), .Z(new_n721));
  AOI22_X1  g296(.A1(new_n720), .A2(G119), .B1(G2104), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(KEYINPUT36), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n711), .B2(new_n712), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n727), .A2(KEYINPUT36), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n717), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G29), .A2(G33), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n479), .A2(G139), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT92), .Z(new_n734));
  INV_X1    g309(.A(G127), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n461), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G115), .B2(G2104), .ZN(new_n737));
  AOI21_X1  g312(.A(KEYINPUT25), .B1(new_n464), .B2(G103), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT25), .ZN(new_n739));
  INV_X1    g314(.A(G103), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n621), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n734), .B1(new_n470), .B2(new_n737), .C1(new_n738), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT93), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n732), .B1(new_n743), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT94), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2072), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G19), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n556), .B2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G1341), .Z(new_n749));
  NAND2_X1  g324(.A1(G164), .A2(G29), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G27), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n749), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G29), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT98), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n758), .A2(new_n757), .A3(G28), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n757), .B2(G28), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n756), .B1(new_n757), .B2(G28), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G11), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n631), .B2(G29), .ZN(new_n764));
  NOR2_X1   g339(.A1(G29), .A2(G35), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G162), .B2(G29), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT29), .Z(new_n767));
  INV_X1    g342(.A(G2090), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n694), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n694), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n764), .B1(new_n767), .B2(new_n768), .C1(G1961), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT26), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n774), .A2(new_n775), .B1(G105), .B2(new_n464), .ZN(new_n776));
  INV_X1    g351(.A(G129), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n474), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n479), .B2(G141), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT95), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n756), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n756), .B2(G32), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n771), .B(new_n784), .C1(new_n768), .C2(new_n767), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT96), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n694), .A2(G20), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT23), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G299), .B2(G16), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1956), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n756), .A2(G26), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT28), .ZN(new_n793));
  MUX2_X1   g368(.A(G104), .B(G116), .S(G2105), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G2104), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT91), .Z(new_n796));
  INV_X1    g371(.A(G140), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n471), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n720), .A2(G128), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(new_n756), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2067), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n770), .A2(G1961), .ZN(new_n803));
  NAND2_X1  g378(.A1(G160), .A2(G29), .ZN(new_n804));
  AND2_X1   g379(.A1(KEYINPUT24), .A2(G34), .ZN(new_n805));
  NOR2_X1   g380(.A1(KEYINPUT24), .A2(G34), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n756), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n804), .A2(G2084), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(G2084), .B1(new_n804), .B2(new_n807), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n791), .A2(new_n802), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n785), .A2(new_n787), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n694), .A2(G4), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n608), .B2(new_n694), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1348), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n746), .A2(new_n755), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n730), .B1(new_n717), .B2(new_n729), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n694), .A2(G21), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G168), .B2(new_n694), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  INV_X1    g395(.A(G1966), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n731), .A2(new_n816), .A3(new_n817), .A4(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  NAND2_X1  g399(.A1(new_n608), .A2(G559), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT38), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT101), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT99), .B(G55), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n530), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  OAI221_X1 g407(.A(new_n830), .B1(new_n545), .B2(new_n831), .C1(new_n590), .C2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n617), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n833), .B1(new_n556), .B2(KEYINPUT100), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n617), .A2(new_n828), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n827), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n840));
  AOI21_X1  g415(.A(G860), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n833), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  XNOR2_X1  g420(.A(new_n723), .B(new_n623), .ZN(new_n846));
  INV_X1    g421(.A(G130), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT104), .B1(new_n470), .B2(G118), .ZN(new_n848));
  OR2_X1    g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(G2104), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n470), .A2(KEYINPUT104), .A3(G118), .ZN(new_n851));
  OAI22_X1  g426(.A1(new_n474), .A2(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n479), .B2(G142), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT105), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n846), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n497), .B1(new_n474), .B2(new_n499), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n486), .B2(new_n488), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n779), .ZN(new_n858));
  INV_X1    g433(.A(new_n800), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n855), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n743), .A2(KEYINPUT95), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(KEYINPUT103), .B2(new_n743), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n861), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G160), .B(G162), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n631), .B(KEYINPUT102), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n864), .A2(new_n867), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g448(.A(new_n618), .B(new_n838), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n607), .A2(G299), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n607), .A2(G299), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  INV_X1    g456(.A(new_n877), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n875), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT41), .B1(new_n882), .B2(new_n875), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(G288), .ZN(new_n889));
  XOR2_X1   g464(.A(G303), .B(G305), .Z(new_n890));
  XOR2_X1   g465(.A(new_n889), .B(new_n890), .Z(new_n891));
  AOI21_X1  g466(.A(new_n881), .B1(new_n880), .B2(new_n886), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n880), .A2(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT42), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n896), .B2(new_n887), .ZN(new_n897));
  OAI21_X1  g472(.A(G868), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n898), .B(KEYINPUT106), .C1(G868), .C2(new_n833), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n891), .B1(new_n888), .B2(new_n892), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n894), .A3(new_n887), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n611), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n833), .A2(G868), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n899), .A2(new_n905), .ZN(G295));
  NOR2_X1   g481(.A1(new_n903), .A2(new_n904), .ZN(G331));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  NAND2_X1  g483(.A1(G168), .A2(G171), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n836), .A2(new_n837), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n834), .ZN(new_n912));
  NOR2_X1   g487(.A1(G168), .A2(G171), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(G286), .A2(G301), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n838), .B1(new_n915), .B2(new_n909), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n885), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n912), .B1(new_n910), .B2(new_n913), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n838), .A3(new_n909), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n878), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n891), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n869), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(KEYINPUT107), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n918), .A2(KEYINPUT108), .A3(new_n878), .A4(new_n919), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n927), .B(new_n885), .C1(new_n914), .C2(new_n916), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n923), .A2(new_n925), .A3(new_n926), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n922), .B1(new_n929), .B2(new_n894), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n922), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n917), .A2(new_n920), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n894), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n908), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n931), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n930), .A2(KEYINPUT109), .A3(new_n931), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(new_n935), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n940), .A2(new_n941), .B1(KEYINPUT43), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n937), .B1(new_n943), .B2(new_n908), .ZN(G397));
  XOR2_X1   g519(.A(KEYINPUT110), .B(G1384), .Z(new_n945));
  NOR2_X1   g520(.A1(new_n857), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(G40), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n472), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G2067), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n800), .B(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT113), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n954), .B2(new_n779), .ZN(new_n955));
  INV_X1    g530(.A(new_n951), .ZN(new_n956));
  INV_X1    g531(.A(G1996), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT112), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n955), .B1(new_n959), .B2(KEYINPUT46), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(KEYINPUT46), .B2(new_n959), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT47), .Z(new_n962));
  OAI21_X1  g537(.A(new_n954), .B1(new_n957), .B2(new_n779), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n963), .A2(new_n956), .B1(new_n959), .B2(new_n780), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n723), .B(new_n725), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT114), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n956), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(G290), .A2(G1986), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(new_n951), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n970), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n719), .A2(new_n722), .A3(new_n725), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n964), .A2(new_n975), .B1(new_n952), .B2(new_n800), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n951), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n962), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(G305), .B(G1981), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  INV_X1    g557(.A(G8), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n857), .A2(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n984), .B2(new_n950), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n696), .A2(G1976), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n988), .A3(new_n987), .ZN(new_n990));
  OR3_X1    g565(.A1(new_n696), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n986), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(G303), .A2(G8), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT115), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT115), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(new_n998), .C1(new_n995), .C2(new_n994), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n489), .B2(new_n502), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n949), .B1(new_n946), .B2(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n708), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n857), .B2(G1384), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT4), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n471), .A2(new_n484), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n482), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n487), .B1(new_n1012), .B2(new_n485), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT69), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n856), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n500), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT50), .B(new_n1009), .C1(new_n1013), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1008), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(new_n768), .A3(new_n950), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n983), .B1(new_n1006), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n999), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n993), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n986), .A2(new_n1023), .A3(new_n696), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(G1981), .B2(G305), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n985), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n993), .A2(KEYINPUT118), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n986), .B(new_n1028), .C1(new_n989), .C2(new_n992), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1029), .A3(new_n1021), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n950), .B1(new_n984), .B2(new_n1007), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT117), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(KEYINPUT50), .B2(new_n1001), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1031), .A2(KEYINPUT117), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1006), .B1(new_n1036), .B2(G2090), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n999), .B1(new_n1037), .B2(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1030), .A2(new_n1038), .ZN(new_n1039));
  AOI211_X1 g614(.A(G2084), .B(new_n949), .C1(new_n1008), .C2(new_n1017), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1002), .B(new_n1009), .C1(new_n1013), .C2(new_n856), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1966), .B1(new_n1042), .B2(new_n950), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1002), .B1(new_n503), .B2(new_n1009), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n857), .A2(KEYINPUT45), .A3(G1384), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n950), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n821), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT119), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n983), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G168), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT63), .B1(new_n1039), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1021), .A2(KEYINPUT63), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n999), .A2(new_n1020), .ZN(new_n1056));
  NOR4_X1   g631(.A1(new_n1055), .A2(new_n1052), .A3(new_n993), .A4(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1026), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n1005), .B2(G2078), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n949), .B1(new_n1008), .B2(new_n1017), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1061), .A2(G1961), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n752), .A2(KEYINPUT53), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1048), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(new_n1064), .B2(KEYINPUT123), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(KEYINPUT123), .B2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G301), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n540), .A2(G8), .A3(new_n541), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT121), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1051), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1048), .A2(new_n1044), .A3(new_n821), .ZN(new_n1072));
  INV_X1    g647(.A(G2084), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1018), .A2(new_n1073), .A3(new_n950), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1069), .B(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(KEYINPUT51), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1070), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1071), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1071), .A2(new_n1080), .A3(KEYINPUT122), .A4(new_n1081), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(KEYINPUT62), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT62), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1067), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n947), .A2(new_n1063), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1004), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT124), .ZN(new_n1091));
  XOR2_X1   g666(.A(G301), .B(KEYINPUT54), .Z(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1062), .A3(new_n1060), .A4(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1066), .B2(new_n1092), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1061), .A2(G1348), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n950), .A2(new_n984), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(G2067), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n607), .B(KEYINPUT60), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n607), .ZN(new_n1101));
  OAI211_X1 g676(.A(KEYINPUT60), .B(new_n1101), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT120), .B(G1996), .Z(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1005), .B2(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1107), .A2(KEYINPUT59), .A3(new_n556), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT59), .B1(new_n1107), .B2(new_n556), .ZN(new_n1109));
  NOR4_X1   g684(.A1(new_n1103), .A2(new_n1108), .A3(new_n1109), .A4(KEYINPUT61), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1098), .A2(new_n607), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n566), .B2(new_n568), .ZN(new_n1112));
  AOI22_X1  g687(.A1(G299), .A2(KEYINPUT57), .B1(new_n575), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT56), .B(G2072), .Z(new_n1115));
  OAI22_X1  g690(.A1(new_n1035), .A2(G1956), .B1(new_n1005), .B2(new_n1115), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1110), .A2(new_n1111), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1116), .A2(new_n1118), .A3(new_n1114), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1103), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1119), .A2(new_n1120), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1094), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1088), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1058), .B1(new_n1125), .B2(new_n1039), .ZN(new_n1126));
  NAND2_X1  g701(.A1(G290), .A2(G1986), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n969), .A2(KEYINPUT111), .A3(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(new_n956), .C1(KEYINPUT111), .C2(new_n1127), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n968), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n978), .B1(new_n1126), .B2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g706(.A1(new_n692), .A2(new_n652), .ZN(new_n1133));
  NAND3_X1  g707(.A1(new_n670), .A2(G319), .A3(new_n671), .ZN(new_n1134));
  XNOR2_X1  g708(.A(new_n1134), .B(KEYINPUT127), .ZN(new_n1135));
  NOR3_X1   g709(.A1(new_n872), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g710(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g711(.A1(new_n943), .A2(new_n1137), .ZN(G308));
  AND2_X1   g712(.A1(new_n940), .A2(new_n941), .ZN(new_n1139));
  AOI21_X1  g713(.A(new_n931), .B1(new_n933), .B2(new_n935), .ZN(new_n1140));
  OAI21_X1  g714(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(G225));
endmodule


