//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1167,
    new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n460), .A2(new_n462), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n463), .A2(new_n469), .ZN(G160));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT67), .Z(G162));
  OR2_X1    g055(.A1(G102), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n483), .B2(new_n484), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n488), .B(new_n491), .C1(new_n484), .C2(new_n483), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n486), .B1(new_n490), .B2(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT6), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(KEYINPUT68), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT6), .A3(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT69), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(KEYINPUT69), .A2(KEYINPUT5), .A3(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n496), .B2(new_n498), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n506), .A2(G88), .B1(G50), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n509), .A2(new_n495), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  NAND2_X1  g087(.A1(new_n506), .A2(G89), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(KEYINPUT70), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n502), .A2(new_n515), .A3(new_n503), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n514), .A2(G63), .A3(G651), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(G51), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n513), .A2(new_n517), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n521), .B(new_n522), .ZN(G168));
  NAND3_X1  g098(.A1(new_n514), .A2(G64), .A3(new_n516), .ZN(new_n524));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n495), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n507), .A2(G52), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n505), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G171));
  NAND3_X1  g105(.A1(new_n514), .A2(G56), .A3(new_n516), .ZN(new_n531));
  NAND2_X1  g106(.A1(G68), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n495), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n507), .A2(G43), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n505), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(new_n533), .B2(new_n536), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n504), .A2(G65), .ZN(new_n548));
  NAND2_X1  g123(.A1(G78), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n495), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT74), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT74), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n551), .A2(new_n552), .B1(G91), .B2(new_n506), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n507), .A2(new_n554), .A3(G53), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n554), .B1(new_n507), .B2(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT73), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OR3_X1    g133(.A1(new_n556), .A2(KEYINPUT73), .A3(new_n557), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n553), .A2(new_n558), .A3(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  XNOR2_X1  g136(.A(new_n521), .B(KEYINPUT71), .ZN(G286));
  NAND2_X1  g137(.A1(new_n514), .A2(new_n516), .ZN(new_n563));
  INV_X1    g138(.A(G74), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n495), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n507), .A2(G49), .ZN(new_n566));
  INV_X1    g141(.A(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n567), .B2(new_n505), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G288));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n505), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n499), .A2(new_n504), .A3(new_n573), .A4(G86), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n572), .A2(new_n574), .B1(G48), .B2(new_n507), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n504), .A2(G61), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n495), .B1(new_n576), .B2(new_n577), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT75), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n575), .A2(new_n581), .A3(new_n583), .ZN(G305));
  NAND3_X1  g159(.A1(new_n514), .A2(G60), .A3(new_n516), .ZN(new_n585));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n495), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n499), .A2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(KEYINPUT77), .B(G47), .Z(new_n590));
  OAI22_X1  g165(.A1(new_n505), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G301), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n504), .A2(G66), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT78), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n507), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n506), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT10), .B1(new_n506), .B2(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(KEYINPUT79), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(KEYINPUT79), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(new_n594), .ZN(G284));
  AOI21_X1  g182(.A(new_n595), .B1(new_n606), .B2(new_n594), .ZN(G321));
  MUX2_X1   g183(.A(G286), .B(G299), .S(new_n594), .Z(G297));
  XOR2_X1   g184(.A(G297), .B(KEYINPUT80), .Z(G280));
  XNOR2_X1  g185(.A(KEYINPUT81), .B(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n606), .B1(G860), .B2(new_n611), .ZN(G148));
  NOR2_X1   g187(.A1(new_n542), .A2(G868), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n604), .A2(new_n605), .A3(new_n611), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(G868), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n475), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n462), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G135), .B2(new_n473), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT84), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND2_X1  g199(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n460), .A2(new_n465), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  NOR2_X1   g203(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n624), .B(new_n630), .C1(new_n628), .C2(new_n625), .ZN(G156));
  XOR2_X1   g206(.A(KEYINPUT15), .B(G2435), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT86), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT87), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n641), .A2(new_n644), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n641), .A2(new_n644), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n651), .A3(G14), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT17), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n657), .B2(new_n654), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n658), .B1(KEYINPUT88), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(KEYINPUT88), .B2(new_n660), .ZN(new_n662));
  INV_X1    g237(.A(new_n654), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n659), .A3(new_n656), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n655), .A2(new_n659), .A3(new_n657), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT89), .ZN(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n680), .C1(new_n671), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n686), .A2(new_n689), .A3(new_n687), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(G229));
  MUX2_X1   g268(.A(G6), .B(G305), .S(G16), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT91), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n569), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n699), .B2(G23), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT33), .B(G1976), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n699), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G1971), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(G1971), .ZN(new_n709));
  NOR4_X1   g284(.A1(new_n704), .A2(new_n705), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n697), .A2(new_n698), .A3(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n592), .A2(new_n699), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n699), .B2(G24), .ZN(new_n715));
  INV_X1    g290(.A(G1986), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT90), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n473), .A2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n475), .A2(G119), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n462), .A2(G107), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n721), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n717), .A2(new_n718), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n712), .A2(new_n713), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n732));
  OR2_X1    g307(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n732), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n712), .A2(new_n735), .A3(new_n713), .A4(new_n730), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n719), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  INV_X1    g314(.A(G139), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n467), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n460), .A2(G127), .ZN(new_n742));
  INV_X1    g317(.A(G115), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n464), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(G2105), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n737), .B1(new_n745), .B2(new_n719), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G2072), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n699), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n606), .B2(new_n699), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT93), .B(G1348), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n699), .A2(G5), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G171), .B2(new_n699), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1961), .ZN(new_n756));
  OR3_X1    g331(.A1(new_n749), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n747), .A2(G2072), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT95), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT29), .ZN(new_n762));
  INV_X1    g337(.A(G2090), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n473), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n475), .A2(G129), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT26), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G32), .B(new_n769), .S(G29), .Z(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n719), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n473), .A2(G140), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n475), .A2(G128), .ZN(new_n776));
  OR2_X1    g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(new_n719), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT30), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n784), .A2(G28), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n719), .B1(new_n784), .B2(G28), .ZN(new_n786));
  AND2_X1   g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  NOR2_X1   g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  OAI22_X1  g363(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT24), .ZN(new_n790));
  INV_X1    g365(.A(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n790), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G160), .B2(new_n719), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(G2084), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n772), .A2(new_n783), .A3(new_n795), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n623), .A2(new_n719), .B1(new_n794), .B2(G2084), .ZN(new_n797));
  NOR2_X1   g372(.A1(G27), .A2(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n796), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n759), .A2(new_n764), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n699), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n542), .B2(new_n699), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1341), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n699), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT23), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n551), .A2(new_n552), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n506), .A2(G91), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n559), .A2(new_n558), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n807), .B1(new_n812), .B2(new_n699), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1956), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n805), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G21), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G168), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT97), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1966), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n757), .A2(new_n802), .A3(new_n815), .A4(new_n819), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n734), .A2(new_n736), .A3(new_n820), .ZN(G311));
  NAND3_X1  g396(.A1(new_n734), .A2(new_n736), .A3(new_n820), .ZN(G150));
  NAND2_X1  g397(.A1(new_n507), .A2(G55), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n505), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT99), .ZN(new_n826));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n563), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G651), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n606), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n538), .A2(new_n540), .B1(new_n826), .B2(new_n830), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n826), .A2(new_n537), .A3(new_n830), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n836), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n841), .A2(KEYINPUT100), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT100), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G860), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n841), .B2(new_n842), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n833), .B1(new_n845), .B2(new_n847), .ZN(G145));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n780), .B(G164), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n769), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n745), .Z(new_n852));
  XOR2_X1   g427(.A(new_n726), .B(KEYINPUT101), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n627), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n473), .A2(G142), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n475), .A2(G130), .ZN(new_n856));
  OR2_X1    g431(.A1(G106), .A2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n857), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n854), .A2(new_n860), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT102), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n861), .B2(new_n862), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n852), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n852), .A2(new_n863), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n623), .B(G160), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(G162), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n849), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n852), .ZN(new_n873));
  INV_X1    g448(.A(new_n866), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n861), .A2(new_n862), .A3(new_n865), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n864), .A2(new_n866), .A3(new_n852), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(G395));
  NAND2_X1  g456(.A1(new_n831), .A2(new_n594), .ZN(new_n882));
  XNOR2_X1  g457(.A(G305), .B(new_n592), .ZN(new_n883));
  XNOR2_X1  g458(.A(G166), .B(new_n569), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT42), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n606), .A2(new_n887), .A3(new_n611), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n614), .A2(KEYINPUT103), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n840), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n840), .A3(new_n889), .ZN(new_n892));
  NAND2_X1  g467(.A1(G299), .A2(new_n603), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(G299), .A2(new_n603), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(KEYINPUT104), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT41), .B1(new_n894), .B2(new_n895), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  INV_X1    g476(.A(new_n603), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n812), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n898), .A3(new_n893), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n892), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n899), .B(new_n905), .C1(new_n906), .C2(new_n890), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n905), .A2(new_n899), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n891), .A2(new_n892), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT105), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n886), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(new_n908), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT105), .ZN(new_n915));
  INV_X1    g490(.A(new_n886), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n897), .A4(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n882), .B1(new_n918), .B2(new_n594), .ZN(G295));
  OAI21_X1  g494(.A(new_n882), .B1(new_n918), .B2(new_n594), .ZN(G331));
  NAND2_X1  g495(.A1(G286), .A2(G301), .ZN(new_n921));
  NAND2_X1  g496(.A1(G168), .A2(G171), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n837), .B2(new_n839), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n840), .A2(new_n921), .A3(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n905), .A2(new_n926), .A3(new_n899), .ZN(new_n927));
  INV_X1    g502(.A(new_n885), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n896), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n925), .A2(new_n924), .B1(new_n900), .B2(new_n904), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n924), .A2(new_n925), .A3(new_n896), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n885), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n933), .A3(new_n849), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n927), .A2(new_n929), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n885), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n849), .A3(new_n930), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n935), .B(KEYINPUT44), .C1(new_n938), .C2(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  AND4_X1   g515(.A1(new_n940), .A2(new_n930), .A3(new_n933), .A4(new_n849), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(KEYINPUT43), .B2(new_n938), .ZN(new_n942));
  XNOR2_X1  g517(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(G397));
  NOR2_X1   g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G164), .B2(G1384), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n948), .B(G40), .C1(new_n462), .C2(new_n461), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n769), .B(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n779), .B(new_n782), .ZN(new_n957));
  INV_X1    g532(.A(new_n728), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n726), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n726), .A2(new_n958), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n956), .A2(new_n957), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n953), .B(new_n954), .C1(new_n950), .C2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n957), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n950), .B1(new_n963), .B2(new_n769), .ZN(new_n964));
  INV_X1    g539(.A(new_n950), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n965), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n950), .B2(new_n955), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT47), .Z(new_n970));
  NAND2_X1  g545(.A1(new_n956), .A2(new_n957), .ZN(new_n971));
  OAI22_X1  g546(.A1(new_n971), .A2(new_n959), .B1(G2067), .B2(new_n779), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n962), .B(new_n970), .C1(new_n950), .C2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n569), .A2(G1976), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n463), .A2(new_n469), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n490), .A2(new_n492), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n482), .A2(new_n485), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G8), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT113), .B(G1976), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(G288), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(new_n982), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n575), .A2(new_n581), .A3(new_n988), .A4(new_n583), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n507), .A2(G48), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n571), .B2(new_n505), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n991), .B2(new_n582), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n981), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(KEYINPUT114), .A3(new_n996), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n987), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1971), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n979), .A2(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n979), .A2(KEYINPUT108), .A3(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n979), .B2(KEYINPUT45), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT107), .B(new_n946), .C1(G164), .C2(G1384), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n976), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1002), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT109), .B(new_n1002), .C1(new_n1007), .C2(new_n1011), .ZN(new_n1015));
  INV_X1    g590(.A(G1384), .ZN(new_n1016));
  INV_X1    g591(.A(new_n492), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n491), .B1(new_n460), .B2(new_n488), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1016), .B1(new_n1019), .B2(new_n486), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n949), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n1022));
  NOR4_X1   g597(.A1(G164), .A2(new_n1022), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT110), .B1(new_n979), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(G2090), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1014), .A2(new_n1015), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n947), .A2(new_n1003), .A3(new_n976), .ZN(new_n1031));
  INV_X1    g606(.A(G1966), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2084), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1021), .B(new_n1034), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1030), .B(G286), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1001), .A2(new_n1029), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n1038));
  OAI22_X1  g613(.A1(G166), .A2(new_n1030), .B1(KEYINPUT111), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(KEYINPUT111), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n1040), .B(KEYINPUT112), .Z(new_n1041));
  XNOR2_X1  g616(.A(new_n1039), .B(new_n1041), .ZN(new_n1042));
  AOI211_X1 g617(.A(KEYINPUT116), .B(new_n1042), .C1(new_n1028), .C2(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT63), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1028), .A2(G8), .A3(new_n1042), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT63), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n979), .A2(new_n1024), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1021), .A2(new_n763), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1030), .B1(new_n1012), .B2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1036), .B(new_n1046), .C1(new_n1049), .C2(new_n1042), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G288), .A2(G1976), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n995), .A2(KEYINPUT114), .A3(new_n996), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT114), .B1(new_n995), .B2(new_n996), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n989), .B(KEYINPUT115), .Z(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n981), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1051), .A2(new_n1001), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1030), .B1(new_n1035), .B2(new_n1033), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT51), .B1(new_n1060), .B2(KEYINPUT124), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1035), .A2(new_n1033), .A3(G168), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1062), .A2(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(G8), .ZN(new_n1065));
  AOI21_X1  g640(.A(G168), .B1(new_n1035), .B2(new_n1033), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1064), .B1(new_n1067), .B2(new_n1061), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT62), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT62), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1064), .B(new_n1070), .C1(new_n1067), .C2(new_n1061), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NOR4_X1   g648(.A1(G164), .A2(new_n1004), .A3(new_n946), .A4(G1384), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT108), .B1(new_n979), .B2(KEYINPUT45), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n979), .A2(KEYINPUT45), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n949), .B1(new_n1077), .B2(KEYINPUT107), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1078), .A3(new_n1009), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1073), .B1(new_n1079), .B2(G2078), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1026), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1961), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1021), .B(KEYINPUT118), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1073), .A2(G2078), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n947), .A2(new_n1003), .A3(new_n976), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1080), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1049), .A2(new_n1042), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(new_n1045), .A3(new_n1001), .A4(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1044), .B(new_n1059), .C1(new_n1072), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1348), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1082), .A2(new_n1093), .A3(new_n1084), .ZN(new_n1094));
  INV_X1    g669(.A(new_n980), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n782), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT60), .B1(new_n603), .B2(KEYINPUT122), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n603), .A2(KEYINPUT122), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1099), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1097), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n557), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n1109), .B2(new_n555), .ZN(new_n1110));
  AOI22_X1  g685(.A1(G299), .A2(KEYINPUT57), .B1(new_n553), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1021), .A2(new_n1047), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1076), .A2(new_n1078), .A3(new_n1116), .A4(new_n1009), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT117), .B1(new_n1120), .B2(new_n1116), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1112), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(KEYINPUT117), .A3(new_n1116), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1111), .A4(new_n1115), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT120), .B(new_n1112), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1124), .A2(KEYINPUT61), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  AOI22_X1  g707(.A1(new_n1120), .A2(new_n955), .B1(new_n980), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(KEYINPUT121), .ZN(new_n1135));
  OR3_X1    g710(.A1(new_n1133), .A2(new_n541), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n1133), .B2(new_n541), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1130), .A2(new_n1131), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT123), .B(new_n1100), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1108), .A2(new_n1129), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1102), .A2(new_n902), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT119), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1127), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1001), .A2(new_n1090), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n461), .A2(KEYINPUT125), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n461), .A2(KEYINPUT125), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n1149), .A3(G2105), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1150), .A2(G40), .A3(new_n948), .A4(new_n1086), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1007), .A2(new_n1077), .A3(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(G171), .B(KEYINPUT54), .Z(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1147), .A2(new_n1154), .B1(new_n1088), .B2(new_n1153), .ZN(new_n1155));
  AND4_X1   g730(.A1(new_n1045), .A2(new_n1146), .A3(new_n1155), .A4(new_n1068), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1092), .B1(new_n1145), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n961), .A2(new_n945), .ZN(new_n1158));
  NAND2_X1  g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n965), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n973), .B1(new_n1157), .B2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g736(.A1(G227), .A2(new_n458), .ZN(new_n1163));
  AOI21_X1  g737(.A(new_n1163), .B1(new_n691), .B2(new_n692), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n1164), .B(new_n652), .C1(new_n878), .C2(new_n872), .ZN(new_n1165));
  NOR2_X1   g739(.A1(new_n942), .A2(new_n1165), .ZN(G308));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n652), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n1167), .A2(new_n879), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n1169));
  OAI21_X1  g743(.A(new_n1169), .B1(KEYINPUT43), .B2(new_n934), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1170), .ZN(G225));
endmodule


