//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT79), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n191), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n191), .B2(new_n195), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n192), .A2(KEYINPUT67), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n191), .A2(new_n200), .A3(new_n202), .A4(new_n195), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n193), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT3), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT78), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT78), .A2(G107), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G107), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n216));
  NAND2_X1  g030(.A1(G104), .A2(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(G101), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n189), .B1(new_n204), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n215), .A2(new_n218), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n191), .A2(new_n195), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G128), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n191), .A2(new_n195), .A3(new_n196), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n203), .ZN(new_n225));
  INV_X1    g039(.A(new_n193), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n221), .A2(KEYINPUT79), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n191), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n200), .A3(new_n202), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n220), .A2(new_n228), .B1(new_n232), .B2(new_n219), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT12), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G137), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT11), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(G137), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT65), .B(new_n240), .C1(new_n235), .C2(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G131), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT66), .B(G131), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n238), .A2(new_n244), .A3(new_n239), .A4(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n233), .A2(new_n234), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n232), .A2(new_n219), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n204), .A2(new_n189), .A3(new_n219), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT79), .B1(new_n221), .B2(new_n227), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n246), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n220), .A2(new_n228), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n249), .B1(new_n255), .B2(new_n250), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n234), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT81), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n259), .B(new_n234), .C1(new_n254), .C2(new_n256), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n248), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT10), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n199), .A2(KEYINPUT0), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n223), .A2(KEYINPUT0), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n267));
  INV_X1    g081(.A(new_n208), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT78), .A2(G107), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n213), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G107), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n211), .B1(new_n206), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n267), .B(G101), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G101), .B1(new_n270), .B2(new_n272), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n266), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n231), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n263), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n246), .ZN(new_n279));
  XNOR2_X1  g093(.A(G110), .B(G140), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n281), .A2(G227), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n280), .B(new_n282), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n261), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n279), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n278), .A2(new_n246), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n283), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n187), .B(new_n188), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n187), .A2(new_n188), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n284), .B1(new_n261), .B2(new_n279), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(new_n283), .A3(new_n289), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(G469), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G221), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT9), .B(G234), .Z(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n188), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(G125), .ZN(new_n305));
  INV_X1    g119(.A(G125), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT74), .B1(new_n306), .B2(G140), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(G140), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n309), .A2(KEYINPUT16), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(KEYINPUT16), .ZN(new_n311));
  OAI21_X1  g125(.A(G146), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n309), .B2(KEYINPUT16), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n194), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(KEYINPUT90), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G237), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n281), .A3(G214), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT88), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G143), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n321), .B(G214), .C1(new_n318), .C2(G143), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n320), .A2(new_n322), .A3(new_n244), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n244), .B1(new_n320), .B2(new_n322), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT17), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(KEYINPUT17), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT90), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n313), .A2(new_n194), .ZN(new_n329));
  AOI211_X1 g143(.A(G146), .B(new_n311), .C1(new_n309), .C2(KEYINPUT16), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n315), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G113), .B(G122), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(new_n205), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n320), .A2(new_n322), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT18), .A3(G131), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n337), .ZN(new_n339));
  INV_X1    g153(.A(new_n309), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(new_n194), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n304), .A2(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n306), .A2(G140), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n342), .A2(new_n343), .A3(new_n194), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n338), .B(new_n339), .C1(new_n341), .C2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n332), .A2(new_n334), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n334), .B1(new_n332), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n188), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G475), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n312), .B1(new_n324), .B2(new_n323), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT19), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n342), .A2(new_n343), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n340), .B2(new_n352), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(G146), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n345), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n334), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(G475), .B1(new_n346), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n359), .A2(new_n360), .A3(new_n188), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n359), .B2(new_n188), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n350), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n268), .A2(new_n269), .ZN(new_n364));
  XNOR2_X1  g178(.A(G116), .B(G122), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT14), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G116), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT14), .A3(G122), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n196), .B2(G143), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n190), .A2(KEYINPUT91), .A3(G128), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n196), .A2(G143), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n375), .A2(new_n235), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n235), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  OAI221_X1 g192(.A(new_n366), .B1(new_n368), .B2(new_n371), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT13), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n375), .A2(new_n380), .B1(new_n196), .B2(G143), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n380), .B2(new_n375), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G134), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n364), .B(new_n365), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n377), .B(KEYINPUT92), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n379), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n299), .A2(G217), .A3(new_n281), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n388), .B(KEYINPUT93), .Z(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n391));
  INV_X1    g205(.A(new_n389), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n392), .B(new_n379), .C1(new_n385), .C2(new_n386), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n387), .A2(new_n391), .A3(new_n389), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n188), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n394), .A2(new_n395), .A3(new_n188), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n363), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G952), .ZN(new_n404));
  AOI211_X1 g218(.A(G953), .B(new_n404), .C1(G234), .C2(G237), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT21), .B(G898), .Z(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n188), .B(new_n281), .C1(G234), .C2(G237), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n302), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n413));
  INV_X1    g227(.A(G119), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G116), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n369), .A2(G119), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT2), .B(G113), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT69), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT69), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT2), .B(G113), .Z(new_n421));
  XNOR2_X1  g235(.A(G116), .B(G119), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n417), .B1(new_n421), .B2(KEYINPUT68), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT68), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n419), .A2(new_n423), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n273), .A3(new_n275), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n421), .A2(new_n420), .A3(new_n422), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT69), .B1(new_n417), .B2(new_n418), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n432));
  INV_X1    g246(.A(G113), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n422), .A2(KEYINPUT5), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n221), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT82), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n439), .A3(new_n437), .ZN(new_n442));
  AND4_X1   g256(.A1(new_n413), .A2(new_n441), .A3(KEYINPUT6), .A4(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n438), .B2(new_n440), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n413), .B1(new_n445), .B2(new_n442), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n231), .A2(new_n306), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n264), .A2(new_n265), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n306), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G224), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n450), .B1(new_n452), .B2(G953), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n438), .A2(new_n444), .A3(new_n440), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n447), .A2(KEYINPUT84), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n442), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT83), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n445), .A2(new_n413), .A3(new_n442), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n460), .A2(new_n456), .A3(new_n457), .A4(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n455), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n439), .B(KEYINPUT8), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n219), .A2(new_n431), .A3(new_n436), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n435), .B(KEYINPUT85), .Z(new_n470));
  XNOR2_X1  g284(.A(new_n434), .B(KEYINPUT86), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n470), .A2(new_n471), .B1(new_n429), .B2(new_n430), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n468), .B(new_n469), .C1(new_n472), .C2(new_n219), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n451), .B1(new_n466), .B2(new_n453), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n467), .A2(new_n473), .A3(new_n474), .A4(new_n442), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n188), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n465), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G210), .B1(G237), .B2(G902), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n465), .A2(new_n479), .A3(new_n477), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n479), .B1(new_n465), .B2(new_n477), .ZN(new_n487));
  AOI211_X1 g301(.A(new_n480), .B(new_n476), .C1(new_n458), .C2(new_n464), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT87), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n239), .ZN(new_n492));
  OAI21_X1  g306(.A(G131), .B1(new_n492), .B2(new_n236), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n231), .A2(new_n245), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n266), .A2(KEYINPUT64), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n264), .A2(KEYINPUT64), .A3(new_n265), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n246), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n266), .A2(new_n246), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n494), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n427), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT29), .ZN(new_n504));
  INV_X1    g318(.A(new_n427), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n505), .A3(new_n494), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT26), .B(G101), .Z(new_n507));
  NAND2_X1  g321(.A1(new_n321), .A2(G210), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n509), .B(new_n510), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n503), .A2(new_n504), .A3(new_n506), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(KEYINPUT28), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n501), .A2(new_n515), .A3(new_n505), .A4(new_n494), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n501), .A2(new_n494), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n514), .A2(new_n516), .B1(new_n427), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n511), .B1(new_n518), .B2(new_n504), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n516), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n498), .A2(new_n427), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n520), .A2(new_n504), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n513), .B(new_n188), .C1(new_n519), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G472), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n525));
  NOR2_X1   g339(.A1(G472), .A2(G902), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n506), .A2(new_n511), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT71), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n506), .A2(new_n530), .A3(new_n511), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n503), .A2(new_n527), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n520), .A2(new_n521), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n512), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n529), .A2(new_n531), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n527), .B1(new_n536), .B2(new_n503), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n526), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT32), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n503), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n529), .A2(new_n531), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT31), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n532), .A3(new_n534), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(KEYINPUT32), .A3(new_n526), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n523), .A2(new_n546), .A3(G472), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n525), .A2(new_n540), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n329), .A2(new_n330), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT23), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n414), .B2(G128), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n414), .A2(G128), .ZN(new_n552));
  MUX2_X1   g366(.A(new_n551), .B(new_n550), .S(new_n552), .Z(new_n553));
  INV_X1    g367(.A(G110), .ZN(new_n554));
  OR3_X1    g368(.A1(new_n414), .A2(KEYINPUT73), .A3(G128), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT73), .B1(new_n414), .B2(G128), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT24), .B(G110), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n553), .A2(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n553), .A2(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n563), .A2(new_n329), .A3(new_n344), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT76), .B1(new_n560), .B2(new_n564), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT75), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT22), .B(G137), .Z(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n561), .A2(new_n565), .A3(new_n562), .A4(new_n571), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT25), .B1(new_n576), .B2(G902), .ZN(new_n577));
  INV_X1    g391(.A(G217), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(G234), .B2(new_n188), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n580), .A3(new_n188), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n575), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT77), .Z(new_n586));
  NOR2_X1   g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n548), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n412), .A2(new_n491), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n394), .A2(new_n395), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n390), .A2(KEYINPUT33), .A3(new_n393), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(G478), .A3(new_n188), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n396), .A2(new_n397), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n363), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT95), .ZN(new_n599));
  INV_X1    g413(.A(new_n489), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n599), .A2(new_n600), .A3(new_n410), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n188), .B1(new_n535), .B2(new_n537), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n602), .A2(G472), .B1(new_n544), .B2(new_n526), .ZN(new_n603));
  AND4_X1   g417(.A1(new_n587), .A2(new_n297), .A3(new_n301), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT96), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  INV_X1    g422(.A(new_n362), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n359), .A2(new_n360), .A3(new_n188), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n609), .A2(new_n610), .B1(G475), .B2(new_n349), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n402), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n489), .A2(new_n409), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NAND2_X1  g430(.A1(new_n561), .A2(new_n565), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n571), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n584), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n582), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n603), .A2(KEYINPUT97), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT97), .B1(new_n603), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n412), .A2(new_n624), .A3(new_n491), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n554), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(G12));
  AND3_X1   g442(.A1(new_n548), .A2(new_n297), .A3(new_n301), .ZN(new_n629));
  INV_X1    g443(.A(G900), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n405), .B1(new_n408), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n612), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n621), .B(new_n485), .C1(new_n487), .C2(new_n488), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n629), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT99), .B(G128), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G30));
  AND2_X1   g451(.A1(new_n297), .A2(new_n301), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n631), .B(KEYINPUT39), .Z(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n640), .A2(KEYINPUT40), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(KEYINPUT40), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n641), .A2(new_n402), .A3(new_n363), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n483), .A2(KEYINPUT100), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n487), .A2(new_n488), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n644), .A2(new_n647), .A3(new_n649), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n485), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n540), .A2(new_n545), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n517), .A2(new_n427), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n511), .B1(new_n657), .B2(new_n506), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n536), .B2(new_n503), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n659), .B2(G902), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n621), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n643), .A2(new_n654), .A3(new_n655), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n190), .ZN(G45));
  INV_X1    g478(.A(new_n631), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n597), .A2(new_n363), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n638), .A2(new_n548), .A3(new_n634), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  INV_X1    g483(.A(new_n248), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n247), .B1(new_n233), .B2(new_n249), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n255), .A2(new_n250), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT80), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n259), .B1(new_n674), .B2(new_n234), .ZN(new_n675));
  INV_X1    g489(.A(new_n260), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n670), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n290), .B1(new_n677), .B2(new_n285), .ZN(new_n678));
  OAI21_X1  g492(.A(G469), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n301), .A3(new_n291), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n679), .A2(new_n291), .A3(KEYINPUT102), .A4(new_n301), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n682), .A2(KEYINPUT103), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT103), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n601), .B(new_n588), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  OAI211_X1 g502(.A(new_n613), .B(new_n588), .C1(new_n684), .C2(new_n685), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NAND2_X1  g504(.A1(new_n682), .A2(new_n683), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n691), .A2(new_n411), .A3(new_n633), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n548), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  XOR2_X1   g508(.A(KEYINPUT104), .B(G472), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n602), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n532), .B1(new_n511), .B2(new_n518), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n526), .B1(new_n697), .B2(new_n537), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n587), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n363), .A2(new_n402), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n363), .A2(KEYINPUT105), .A3(new_n402), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT106), .B1(new_n489), .B2(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n363), .A2(KEYINPUT105), .A3(new_n402), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT105), .B1(new_n363), .B2(new_n402), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n483), .A2(new_n710), .A3(new_n711), .A4(new_n485), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n701), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n410), .B(new_n713), .C1(new_n684), .C2(new_n685), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NOR2_X1   g529(.A1(new_n699), .A2(new_n666), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n682), .A2(new_n634), .A3(new_n683), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  XNOR2_X1  g532(.A(new_n545), .B(KEYINPUT108), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n525), .A2(new_n547), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n540), .A3(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n721), .A2(KEYINPUT42), .A3(new_n587), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n678), .A2(G902), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n292), .B1(new_n723), .B2(new_n187), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n294), .A2(KEYINPUT107), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n726), .B(new_n284), .C1(new_n261), .C2(new_n279), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n725), .A2(G469), .A3(new_n295), .A4(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n300), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n483), .A2(new_n655), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n667), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n588), .A3(new_n667), .A4(new_n730), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n722), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(G131), .Z(G33));
  NAND4_X1  g550(.A1(new_n729), .A2(new_n588), .A3(new_n632), .A4(new_n730), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  NAND2_X1  g552(.A1(new_n597), .A2(new_n611), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT43), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n597), .A2(new_n741), .A3(new_n611), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n603), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n621), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  INV_X1    g562(.A(new_n730), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n291), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n294), .A2(new_n295), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n187), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n725), .A2(KEYINPUT45), .A3(new_n295), .A4(new_n727), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT109), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n292), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n751), .B1(new_n760), .B2(KEYINPUT46), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT109), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT109), .B1(new_n754), .B2(new_n755), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n293), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n300), .B1(new_n761), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT110), .B1(new_n767), .B2(new_n639), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT46), .B(new_n293), .C1(new_n762), .C2(new_n763), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n291), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n758), .A2(new_n759), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT46), .B1(new_n771), .B2(new_n293), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n301), .B(new_n639), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n750), .B1(new_n768), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  NOR3_X1   g591(.A1(new_n548), .A2(new_n587), .A3(new_n666), .ZN(new_n778));
  OAI211_X1 g592(.A(KEYINPUT47), .B(new_n301), .C1(new_n770), .C2(new_n772), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n766), .A2(new_n291), .A3(new_n769), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT47), .B1(new_n781), .B2(new_n301), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n730), .B(new_n778), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT111), .B(G140), .Z(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G42));
  NAND2_X1  g599(.A1(new_n679), .A2(new_n291), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT49), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n739), .A2(new_n655), .A3(new_n300), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n587), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT112), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n653), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n656), .A2(new_n660), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n791), .B(new_n792), .C1(KEYINPUT49), .C2(new_n786), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n686), .A2(new_n693), .A3(new_n689), .A4(new_n714), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n707), .A2(new_n712), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n665), .A3(new_n661), .A4(new_n729), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n629), .B(new_n634), .C1(new_n632), .C2(new_n667), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n717), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n796), .A2(KEYINPUT52), .A3(new_n797), .A4(new_n717), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n700), .A2(new_n621), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n731), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n412), .B(new_n491), .C1(new_n624), .C2(new_n588), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n598), .A2(new_n612), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n604), .A2(new_n491), .A3(new_n410), .A4(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n621), .A2(new_n403), .A3(new_n665), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n629), .A2(new_n730), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n809), .A3(new_n737), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n735), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n794), .A2(new_n802), .A3(new_n806), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n804), .B(KEYINPUT113), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n686), .A2(new_n693), .A3(new_n689), .A4(new_n714), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n635), .A2(new_n668), .A3(new_n717), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT52), .A4(new_n796), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n800), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n820), .A2(new_n825), .A3(KEYINPUT53), .A4(new_n813), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n816), .A2(new_n817), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n794), .A2(new_n806), .A3(new_n813), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n823), .A2(new_n824), .A3(new_n800), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n815), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n814), .A2(new_n815), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT115), .B(new_n815), .C1(new_n828), .C2(new_n829), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n827), .B1(new_n835), .B2(KEYINPUT54), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n301), .B1(new_n770), .B2(new_n772), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT47), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n839), .B(new_n779), .C1(new_n301), .C2(new_n786), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n740), .A2(new_n405), .A3(new_n742), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n701), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n730), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n651), .A2(new_n842), .A3(new_n655), .A4(new_n652), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(new_n691), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n844), .B(KEYINPUT50), .C1(new_n845), .C2(new_n691), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n843), .A2(KEYINPUT51), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n691), .A2(new_n749), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n405), .A3(new_n743), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n803), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n792), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n587), .A2(new_n405), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n363), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n597), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n848), .A2(new_n862), .A3(new_n850), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n843), .B(new_n860), .C1(new_n861), .C2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n852), .A2(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n721), .A2(new_n587), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n854), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT48), .Z(new_n869));
  NAND4_X1  g683(.A1(new_n842), .A2(new_n600), .A3(new_n682), .A4(new_n683), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(G952), .A3(new_n281), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n856), .A2(new_n857), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n872), .B2(new_n599), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT118), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n836), .A2(new_n866), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n793), .B1(new_n876), .B2(new_n877), .ZN(G75));
  NAND2_X1  g692(.A1(new_n447), .A2(new_n457), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(new_n456), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT55), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(KEYINPUT119), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(G210), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n884), .B(new_n188), .C1(new_n816), .C2(new_n826), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n188), .B1(new_n816), .B2(new_n826), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(G210), .ZN(new_n888));
  INV_X1    g702(.A(new_n883), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n882), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n404), .A2(G953), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT120), .Z(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n886), .A2(new_n890), .A3(new_n895), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(G51));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n188), .B(new_n771), .C1(new_n816), .C2(new_n826), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n292), .B(KEYINPUT57), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n817), .B1(new_n816), .B2(new_n826), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n827), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n678), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n892), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n816), .A2(new_n826), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n816), .A2(new_n826), .A3(new_n817), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n678), .B1(new_n910), .B2(new_n900), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT122), .B(new_n892), .C1(new_n911), .C2(new_n899), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n887), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n346), .A2(new_n358), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n905), .B1(new_n916), .B2(new_n917), .ZN(G60));
  XNOR2_X1  g732(.A(new_n594), .B(KEYINPUT123), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n836), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n921), .ZN(new_n923));
  INV_X1    g737(.A(new_n919), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n910), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n922), .A2(new_n892), .A3(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n907), .A2(new_n619), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n907), .A2(new_n928), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n892), .B(new_n929), .C1(new_n930), .C2(new_n575), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT61), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G66));
  NAND3_X1  g748(.A1(new_n794), .A2(new_n807), .A3(new_n809), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n281), .ZN(new_n936));
  OAI21_X1  g750(.A(G953), .B1(new_n407), .B2(new_n452), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n879), .B1(G898), .B2(new_n281), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  NAND2_X1  g754(.A1(new_n500), .A2(new_n502), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n354), .ZN(new_n942));
  NAND2_X1  g756(.A1(G900), .A2(G953), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n776), .A2(new_n783), .ZN(new_n944));
  INV_X1    g758(.A(new_n821), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n735), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n867), .B1(new_n712), .B2(new_n707), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n768), .B2(new_n775), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n944), .A2(new_n737), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n942), .B(new_n943), .C1(new_n949), .C2(G953), .ZN(new_n950));
  INV_X1    g764(.A(new_n663), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n821), .A3(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n663), .B2(new_n945), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n954), .A2(new_n776), .A3(new_n783), .A4(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n640), .A2(new_n749), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n958), .A2(new_n588), .A3(new_n808), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n281), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n942), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n950), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n964), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n950), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(G72));
  NAND2_X1  g782(.A1(new_n503), .A2(new_n506), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(new_n511), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n776), .A2(new_n948), .A3(new_n737), .A4(new_n783), .ZN(new_n971));
  INV_X1    g785(.A(new_n946), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n935), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n970), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n969), .ZN(new_n979));
  OAI22_X1  g793(.A1(new_n979), .A2(new_n511), .B1(new_n541), .B2(new_n542), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n835), .A2(new_n976), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(new_n892), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n979), .A2(new_n512), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n957), .A2(new_n935), .A3(new_n959), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n977), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g801(.A(KEYINPUT127), .B(new_n983), .C1(new_n984), .C2(new_n977), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n987), .B2(new_n988), .ZN(G57));
endmodule


