//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(KEYINPUT64), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(KEYINPUT64), .B2(new_n457), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  INV_X1    g043(.A(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(G2104), .ZN(new_n470));
  OAI22_X1  g045(.A1(new_n467), .A2(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n472), .B1(new_n465), .B2(G125), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n466), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n471), .B1(new_n474), .B2(KEYINPUT66), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n476), .B1(new_n473), .B2(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(G160));
  INV_X1    g054(.A(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  MUX2_X1   g059(.A(G100), .B(G112), .S(G2105), .Z(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2104), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n489), .B(new_n490), .C1(new_n463), .C2(new_n464), .ZN(new_n491));
  AND2_X1   g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n466), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n463), .B2(new_n464), .ZN(new_n495));
  AND2_X1   g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n489), .B1(new_n467), .B2(new_n490), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n493), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI211_X1 g077(.A(KEYINPUT69), .B(new_n501), .C1(new_n502), .C2(KEYINPUT68), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(G543), .B1(new_n502), .B2(KEYINPUT69), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n511), .A2(new_n520), .ZN(G166));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n517), .A2(KEYINPUT70), .A3(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n512), .A2(new_n513), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n501), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT69), .B1(new_n502), .B2(KEYINPUT68), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n527), .B1(new_n530), .B2(new_n503), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n508), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n526), .A2(new_n532), .A3(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n540));
  AND2_X1   g115(.A1(G77), .A2(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n508), .B2(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n542), .B2(new_n510), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n530), .B2(new_n503), .ZN(new_n545));
  OAI211_X1 g120(.A(KEYINPUT71), .B(G651), .C1(new_n545), .C2(new_n541), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(G52), .A2(new_n525), .B1(new_n531), .B2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(G43), .A2(new_n525), .B1(new_n531), .B2(G81), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n530), .B2(new_n503), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  NAND3_X1  g139(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n518), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n531), .A2(KEYINPUT72), .A3(G91), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n530), .B2(new_n503), .ZN(new_n575));
  AND2_X1   g150(.A1(G78), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n508), .A2(G65), .ZN(new_n578));
  INV_X1    g153(.A(new_n576), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(KEYINPUT73), .A3(new_n579), .ZN(new_n580));
  AND4_X1   g155(.A1(KEYINPUT74), .A2(new_n577), .A3(G651), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n576), .B1(new_n508), .B2(G65), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n510), .B1(new_n582), .B2(KEYINPUT73), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT74), .B1(new_n583), .B2(new_n577), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n572), .B1(new_n581), .B2(new_n584), .ZN(G299));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n547), .A2(new_n586), .A3(new_n548), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n586), .B1(new_n547), .B2(new_n548), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(G301));
  OR2_X1    g164(.A1(new_n511), .A2(new_n520), .ZN(G303));
  NAND2_X1  g165(.A1(new_n531), .A2(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n515), .A2(G49), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  NAND2_X1  g169(.A1(new_n515), .A2(G48), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  OAI221_X1 g172(.A(new_n595), .B1(new_n518), .B2(new_n596), .C1(new_n597), .C2(new_n510), .ZN(G305));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n525), .A2(G47), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n531), .A2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g177(.A1(G72), .A2(G543), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n508), .B2(G60), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n510), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n604), .A2(new_n510), .ZN(new_n607));
  AOI22_X1  g182(.A1(G47), .A2(new_n525), .B1(new_n531), .B2(G85), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT76), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  AOI21_X1  g186(.A(KEYINPUT10), .B1(new_n531), .B2(G92), .ZN(new_n612));
  AND4_X1   g187(.A1(KEYINPUT10), .A2(new_n508), .A3(G92), .A4(new_n517), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT77), .B(G66), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n530), .B2(new_n503), .ZN(new_n616));
  AND2_X1   g191(.A1(G79), .A2(G543), .ZN(new_n617));
  OAI21_X1  g192(.A(G651), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n525), .A2(G54), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n611), .B1(G868), .B2(new_n621), .ZN(G284));
  XOR2_X1   g197(.A(G284), .B(KEYINPUT78), .Z(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT79), .ZN(new_n625));
  INV_X1    g200(.A(G299), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n621), .B1(new_n629), .B2(G860), .ZN(G148));
  NOR2_X1   g205(.A1(new_n557), .A2(G868), .ZN(new_n631));
  INV_X1    g206(.A(new_n621), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(G559), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n631), .B1(new_n633), .B2(G868), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n480), .A2(G2104), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OAI22_X1  g214(.A1(new_n637), .A2(new_n638), .B1(KEYINPUT80), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n638), .B2(new_n637), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n641), .A2(KEYINPUT80), .A3(new_n639), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(KEYINPUT80), .B2(new_n639), .ZN(new_n643));
  MUX2_X1   g218(.A(G99), .B(G111), .S(G2105), .Z(new_n644));
  AOI22_X1  g219(.A1(new_n480), .A2(G135), .B1(G2104), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n483), .A2(KEYINPUT81), .A3(G123), .ZN(new_n646));
  AOI21_X1  g221(.A(KEYINPUT81), .B1(new_n483), .B2(G123), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2096), .ZN(new_n649));
  OR3_X1    g224(.A1(new_n642), .A2(new_n643), .A3(new_n649), .ZN(G156));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  INV_X1    g227(.A(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2427), .ZN(new_n655));
  INV_X1    g230(.A(G2430), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n658), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(new_n672), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n675), .B2(new_n676), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n670), .A2(new_n672), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n671), .B1(new_n680), .B2(KEYINPUT17), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n674), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G2096), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n639), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n691), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT20), .Z(new_n695));
  AOI211_X1 g270(.A(new_n693), .B(new_n695), .C1(new_n688), .C2(new_n692), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT83), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT84), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n698), .B(new_n703), .ZN(G229));
  XOR2_X1   g279(.A(KEYINPUT85), .B(G16), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G23), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT88), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(G288), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT33), .B(G1976), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT89), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G6), .A2(G16), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n597), .A2(new_n510), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n595), .B1(new_n518), .B2(new_n596), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n719), .B1(new_n722), .B2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT87), .B(KEYINPUT34), .Z(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT90), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n705), .A2(G24), .ZN(new_n730));
  XNOR2_X1  g305(.A(G290), .B(KEYINPUT86), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n705), .ZN(new_n732));
  INV_X1    g307(.A(G1986), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G131), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n483), .A2(G119), .ZN(new_n736));
  AND2_X1   g311(.A1(G107), .A2(G2105), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G95), .B2(new_n466), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n736), .C1(new_n462), .C2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G25), .B(new_n739), .S(G29), .Z(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n726), .B2(new_n727), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n729), .A2(new_n734), .A3(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n748));
  INV_X1    g323(.A(G103), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n470), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n470), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n751), .A2(KEYINPUT25), .A3(G103), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n480), .A2(G139), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n466), .B2(new_n754), .ZN(new_n755));
  MUX2_X1   g330(.A(G33), .B(new_n755), .S(G29), .Z(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G2072), .Z(new_n757));
  NAND2_X1  g332(.A1(G164), .A2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G27), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n648), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n759), .A2(new_n760), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n757), .A2(new_n761), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G29), .A2(G35), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G162), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT29), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2090), .ZN(new_n772));
  INV_X1    g347(.A(G141), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n751), .B2(G105), .ZN(new_n775));
  INV_X1    g350(.A(G105), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n470), .A2(KEYINPUT93), .A3(new_n776), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n467), .A2(new_n773), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT26), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G129), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n482), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n784));
  OR3_X1    g359(.A1(new_n778), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n778), .B2(new_n783), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G32), .B(new_n787), .S(G29), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n772), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G1348), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n621), .A2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G4), .B2(G16), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n768), .B(new_n791), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(G168), .A2(G16), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT95), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT95), .B1(G16), .B2(G21), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G1966), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n763), .A2(G26), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT28), .ZN(new_n804));
  MUX2_X1   g379(.A(G104), .B(G116), .S(G2105), .Z(new_n805));
  AOI22_X1  g380(.A1(new_n483), .A2(G128), .B1(G2104), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G140), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n467), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G29), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(KEYINPUT92), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(KEYINPUT92), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n804), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G2067), .Z(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n792), .B2(new_n794), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n706), .A2(G19), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n558), .B2(new_n706), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1341), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n800), .A2(G1966), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n814), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n795), .A2(new_n802), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n705), .A2(G20), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT97), .B(KEYINPUT23), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G299), .B2(G16), .ZN(new_n824));
  INV_X1    g399(.A(G1956), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(G160), .A2(G29), .ZN(new_n827));
  AND2_X1   g402(.A1(KEYINPUT24), .A2(G34), .ZN(new_n828));
  NOR2_X1   g403(.A1(KEYINPUT24), .A2(G34), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n763), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(G2084), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G1961), .ZN(new_n832));
  NOR2_X1   g407(.A1(G171), .A2(new_n713), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G5), .B2(new_n713), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n827), .A2(G2084), .A3(new_n830), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n835), .B(new_n836), .C1(new_n832), .C2(new_n834), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n820), .A2(new_n826), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n745), .A2(new_n746), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n747), .A2(new_n838), .A3(new_n839), .ZN(G150));
  INV_X1    g415(.A(G150), .ZN(G311));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n842));
  AND2_X1   g417(.A1(G80), .A2(G543), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n508), .B2(G67), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n844), .B2(new_n510), .ZN(new_n845));
  INV_X1    g420(.A(G67), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n530), .B2(new_n503), .ZN(new_n847));
  OAI211_X1 g422(.A(KEYINPUT98), .B(G651), .C1(new_n847), .C2(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n525), .A2(G55), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n531), .A2(G93), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n851), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n845), .B2(new_n848), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n525), .A2(G43), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n531), .A2(G81), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n508), .A2(G56), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n510), .B1(new_n862), .B2(new_n554), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT99), .B1(new_n551), .B2(new_n556), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n857), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n861), .B1(new_n860), .B2(new_n863), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n551), .A2(KEYINPUT99), .A3(new_n556), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n853), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n629), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(G860), .B1(new_n874), .B2(KEYINPUT39), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n875), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n855), .B1(new_n877), .B2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(new_n787), .B(new_n499), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n808), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n637), .B(new_n739), .ZN(new_n883));
  MUX2_X1   g458(.A(G106), .B(G118), .S(G2105), .Z(new_n884));
  AOI22_X1  g459(.A1(new_n483), .A2(G130), .B1(G2104), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G142), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n886), .B2(new_n467), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n883), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n882), .A2(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n755), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(KEYINPUT102), .B2(new_n755), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n892), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n895), .B1(new_n898), .B2(new_n890), .ZN(new_n899));
  XNOR2_X1  g474(.A(G160), .B(new_n487), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n648), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n897), .B2(new_n899), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g484(.A1(G290), .A2(G288), .ZN(new_n910));
  INV_X1    g485(.A(G288), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n606), .A2(new_n609), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G303), .A2(G305), .ZN(new_n914));
  NAND2_X1  g489(.A1(G166), .A2(new_n722), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT103), .B1(new_n913), .B2(new_n916), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n606), .A2(new_n609), .A3(new_n911), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n911), .B1(new_n606), .B2(new_n609), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n916), .B(KEYINPUT103), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n870), .B(new_n633), .Z(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(G299), .A2(new_n632), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n621), .B(new_n572), .C1(new_n581), .C2(new_n584), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n926), .A3(new_n928), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n927), .A2(new_n928), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n925), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT104), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n934), .B2(new_n924), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n935), .A2(KEYINPUT104), .ZN(new_n938));
  OAI21_X1  g513(.A(G868), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(G868), .B2(new_n857), .ZN(G295));
  OAI21_X1  g515(.A(new_n939), .B1(G868), .B2(new_n857), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n587), .A2(new_n588), .A3(G286), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n549), .A2(G168), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n943), .A2(new_n870), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n547), .A2(new_n586), .A3(new_n548), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(G168), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n944), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n948), .A2(new_n949), .B1(new_n866), .B2(new_n869), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n927), .A2(new_n926), .A3(new_n928), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n945), .A2(new_n950), .B1(new_n951), .B2(new_n929), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n870), .B1(new_n943), .B2(new_n944), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n948), .A2(new_n949), .A3(new_n866), .A4(new_n869), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n933), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n923), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n923), .A3(new_n955), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n913), .A2(new_n916), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n913), .A2(new_n916), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n960), .B1(new_n963), .B2(new_n921), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n930), .A2(new_n931), .B1(new_n953), .B2(new_n954), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n953), .A2(new_n933), .A3(new_n954), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n964), .B(new_n957), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n903), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT43), .B1(new_n959), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(new_n903), .A3(new_n958), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n942), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n967), .A2(new_n903), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n958), .A2(new_n957), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n970), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n976), .A2(new_n978), .A3(KEYINPUT106), .A4(new_n979), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n975), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n973), .B1(new_n984), .B2(new_n942), .ZN(G397));
  NAND4_X1  g560(.A1(new_n475), .A2(KEYINPUT107), .A3(G40), .A4(new_n477), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n470), .A2(new_n469), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n480), .B2(G137), .ZN(new_n988));
  INV_X1    g563(.A(G125), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n463), .B2(new_n464), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT66), .B(G2105), .C1(new_n990), .C2(new_n472), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n988), .A2(new_n477), .A3(G40), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n986), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT45), .B1(new_n499), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(G1996), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n787), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n998), .B(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n808), .B(G2067), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(G1996), .A3(new_n787), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n739), .B(new_n742), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n1002), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n998), .A2(G1986), .A3(G290), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n999), .B1(KEYINPUT124), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(KEYINPUT124), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1014), .B(new_n1015), .Z(new_n1016));
  OAI21_X1  g591(.A(new_n1002), .B1(new_n787), .B2(new_n1003), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n739), .A2(new_n742), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n1006), .A2(new_n1021), .B1(G2067), .B2(new_n808), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n1012), .B(new_n1020), .C1(new_n1002), .C2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n499), .A2(new_n996), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n995), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1026), .B2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  AOI211_X1 g603(.A(KEYINPUT110), .B(new_n1028), .C1(new_n995), .C2(new_n1025), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G288), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G303), .A2(G8), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n1034), .B(KEYINPUT55), .Z(new_n1035));
  AND3_X1   g610(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n996), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(new_n997), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1971), .B1(new_n1037), .B2(new_n995), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1025), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n499), .A2(new_n996), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n995), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1038), .A2(KEYINPUT109), .B1(new_n1043), .B2(G2090), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1037), .A2(new_n995), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1045), .A2(KEYINPUT109), .A3(new_n709), .ZN(new_n1046));
  OAI211_X1 g621(.A(G8), .B(new_n1035), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1048));
  OAI221_X1 g623(.A(new_n1048), .B1(new_n1031), .B2(G288), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT111), .B1(G305), .B2(G1981), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n720), .A2(new_n721), .A3(G1981), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(G305), .A2(KEYINPUT111), .A3(G1981), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT49), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(new_n1056), .A3(new_n1053), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1055), .B(new_n1057), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1033), .A2(new_n1047), .A3(new_n1049), .A4(new_n1058), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1035), .B1(new_n1060), .B2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(G1966), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1045), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n986), .A2(new_n994), .B1(KEYINPUT50), .B2(new_n1041), .ZN(new_n1064));
  INV_X1    g639(.A(G2084), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(new_n1040), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1028), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1068));
  OR3_X1    g643(.A1(new_n1059), .A2(new_n1061), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1064), .A2(new_n1070), .B1(new_n1039), .B2(new_n1025), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n995), .A2(new_n1042), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1045), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1074), .A2(G2090), .B1(G1971), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1035), .B1(new_n1076), .B2(G8), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1066), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1966), .B1(new_n1037), .B2(new_n995), .ZN(new_n1079));
  OAI21_X1  g654(.A(G8), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR4_X1   g655(.A1(new_n1059), .A2(new_n1077), .A3(G286), .A4(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1069), .B1(new_n1081), .B2(KEYINPUT63), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G288), .A2(G1976), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1058), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1030), .B1(new_n1084), .B2(new_n1051), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1033), .A2(new_n1049), .A3(new_n1058), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1086), .B(KEYINPUT112), .C1(new_n1047), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1047), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1085), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1059), .A2(new_n1077), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1037), .A2(new_n760), .A3(new_n995), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1043), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1064), .A2(KEYINPUT115), .A3(new_n1040), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n832), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1063), .A2(new_n1102), .A3(new_n1066), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1104));
  OAI21_X1  g679(.A(G8), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G286), .A2(G8), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1101), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1080), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT120), .B1(new_n1067), .B2(new_n1109), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1107), .A2(new_n1113), .B1(G168), .B2(new_n1105), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1093), .B(new_n1100), .C1(new_n1114), .C2(KEYINPUT62), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1114), .A2(KEYINPUT62), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1082), .B(new_n1092), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1026), .A2(G2067), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(G1348), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n621), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n632), .B(new_n1119), .C1(new_n1120), .C2(G1348), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT118), .B(KEYINPUT61), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1074), .A2(new_n825), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n1127));
  NAND2_X1  g702(.A1(G299), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT57), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1075), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1128), .B(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1956), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1075), .A2(new_n1130), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1125), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1026), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(G1996), .B2(new_n1045), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1141), .A2(new_n558), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1141), .B2(new_n558), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n621), .A2(new_n1118), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1143), .A2(new_n1144), .B1(new_n1121), .B2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1124), .A2(new_n1138), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT116), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1135), .A2(new_n1136), .A3(KEYINPUT116), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1134), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(KEYINPUT61), .A3(new_n1132), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1122), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1147), .A2(new_n1152), .B1(new_n1153), .B2(new_n1132), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1113), .B1(new_n1155), .B2(KEYINPUT51), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1105), .A2(G168), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT53), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n760), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n474), .A2(new_n471), .A3(new_n1160), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1094), .A2(new_n1159), .B1(new_n1037), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1099), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1158), .B1(new_n1163), .B2(G171), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1095), .A2(G301), .A3(new_n1099), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1168));
  OAI22_X1  g743(.A1(new_n1156), .A2(new_n1157), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1099), .A2(G301), .A3(new_n1162), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1158), .B1(new_n1100), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(KEYINPUT121), .B(new_n1158), .C1(new_n1100), .C2(new_n1170), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1173), .A2(new_n1093), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1154), .B1(new_n1176), .B2(KEYINPUT123), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1117), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G290), .B(new_n733), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1008), .B1(new_n998), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1023), .B1(new_n1180), .B2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n1185));
  NOR2_X1   g759(.A1(new_n959), .A2(new_n968), .ZN(new_n1186));
  AOI21_X1  g760(.A(KEYINPUT106), .B1(new_n1186), .B2(new_n979), .ZN(new_n1187));
  INV_X1    g761(.A(new_n983), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n974), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n685), .A2(new_n459), .A3(new_n668), .ZN(new_n1190));
  XOR2_X1   g764(.A(new_n1190), .B(KEYINPUT126), .Z(new_n1191));
  NOR2_X1   g765(.A1(new_n1191), .A2(G229), .ZN(new_n1192));
  OAI21_X1  g766(.A(new_n1192), .B1(new_n904), .B2(new_n906), .ZN(new_n1193));
  INV_X1    g767(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g768(.A(new_n1185), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g769(.A1(new_n984), .A2(KEYINPUT127), .A3(new_n1193), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1195), .A2(new_n1196), .ZN(G308));
  NAND2_X1  g771(.A1(new_n1189), .A2(new_n1194), .ZN(G225));
endmodule


