//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT89), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT89), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT15), .A3(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT14), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT90), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n206), .B(KEYINPUT14), .Z(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT91), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT91), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n209), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n205), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n211), .A2(new_n217), .A3(KEYINPUT17), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(KEYINPUT93), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n211), .A2(new_n217), .A3(KEYINPUT92), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT92), .B1(new_n211), .B2(new_n217), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G1gat), .B2(new_n224), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n227), .B(G8gat), .Z(new_n228));
  NAND2_X1  g027(.A1(new_n218), .A2(KEYINPUT93), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n219), .A2(new_n223), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n221), .A2(new_n222), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(new_n228), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT18), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n231), .B(new_n228), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n234), .B(KEYINPUT13), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G169gat), .B(G197gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT88), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n235), .A2(new_n249), .A3(new_n238), .A4(new_n241), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G230gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G85gat), .A2(G92gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT96), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT7), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT96), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n258), .B(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT7), .ZN(new_n264));
  INV_X1    g063(.A(G85gat), .ZN(new_n265));
  INV_X1    g064(.A(G92gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G99gat), .ZN(new_n268));
  INV_X1    g067(.A(G106gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT8), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n261), .A2(new_n264), .A3(new_n267), .A4(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G99gat), .B(G106gat), .Z(new_n272));
  OR2_X1    g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n272), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT97), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G57gat), .B(G64gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT94), .ZN(new_n279));
  NAND2_X1  g078(.A1(G71gat), .A2(G78gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(G71gat), .A2(G78gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(KEYINPUT9), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  AOI211_X1 g083(.A(new_n281), .B(new_n282), .C1(new_n278), .C2(KEYINPUT9), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT97), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n277), .A2(KEYINPUT10), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n286), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n275), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT10), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(new_n273), .A3(new_n274), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n257), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n257), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(new_n290), .B2(new_n292), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G120gat), .B(G148gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT100), .ZN(new_n299));
  INV_X1    g098(.A(G176gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G204gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n297), .A2(new_n304), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n254), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G8gat), .B(G36gat), .Z(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(G64gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(new_n266), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT27), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n320));
  INV_X1    g119(.A(G190gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT67), .A4(new_n321), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT68), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT27), .B(G183gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT28), .A3(new_n321), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n324), .A2(new_n331), .A3(new_n325), .A4(new_n326), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT26), .ZN(new_n335));
  NAND2_X1  g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n335), .A2(new_n336), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G183gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n321), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341));
  NAND2_X1  g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT64), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n342), .A2(new_n343), .A3(new_n341), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n342), .B2(new_n341), .ZN(new_n345));
  OAI221_X1 g144(.A(new_n340), .B1(new_n341), .B2(new_n342), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n336), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT65), .ZN(new_n353));
  OAI211_X1 g152(.A(G183gat), .B(G190gat), .C1(new_n353), .C2(KEYINPUT24), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n342), .A2(KEYINPUT65), .A3(new_n341), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n354), .A2(new_n355), .A3(new_n340), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT25), .B1(new_n349), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n316), .B1(new_n338), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n333), .B2(new_n337), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n315), .B1(new_n360), .B2(KEYINPUT29), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT22), .ZN(new_n364));
  NAND2_X1  g163(.A1(G211gat), .A2(G218gat), .ZN(new_n365));
  INV_X1    g164(.A(G211gat), .ZN(new_n366));
  INV_X1    g165(.A(G218gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT73), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT73), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n364), .A2(new_n371), .A3(new_n365), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT22), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n365), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n363), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT74), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n378), .A3(new_n363), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n362), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n359), .A2(new_n361), .A3(new_n381), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n314), .B1(new_n385), .B2(KEYINPUT37), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n359), .A2(new_n361), .A3(new_n381), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n359), .B2(new_n361), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT37), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT85), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND4_X1   g190(.A1(KEYINPUT85), .A2(new_n383), .A3(new_n390), .A4(new_n384), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT38), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n383), .A2(new_n384), .A3(new_n314), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396));
  INV_X1    g195(.A(G120gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G113gat), .ZN(new_n398));
  INV_X1    g197(.A(G113gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G120gat), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT69), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT1), .ZN(new_n403));
  XNOR2_X1  g202(.A(G127gat), .B(G134gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n407));
  AND2_X1   g206(.A1(G127gat), .A2(G134gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(G127gat), .A2(G134gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G113gat), .B(G120gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(KEYINPUT1), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n406), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n407), .B1(new_n406), .B2(new_n412), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n416));
  INV_X1    g215(.A(G148gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G141gat), .ZN(new_n418));
  INV_X1    g217(.A(G141gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G148gat), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n416), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n420), .A3(new_n416), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT2), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G155gat), .B(G162gat), .Z(new_n426));
  INV_X1    g225(.A(G155gat), .ZN(new_n427));
  INV_X1    g226(.A(G162gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n418), .A2(new_n420), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n425), .A2(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n396), .B1(new_n415), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n406), .A2(new_n412), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(KEYINPUT76), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n406), .A2(new_n407), .A3(new_n412), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n425), .A2(new_n426), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n430), .A2(new_n431), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(KEYINPUT78), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n433), .A2(new_n436), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G225gat), .A2(G233gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n445), .B(KEYINPUT77), .Z(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n436), .A2(KEYINPUT4), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n449), .A3(new_n435), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n446), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n442), .A2(KEYINPUT3), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT3), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n455), .A3(new_n439), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n451), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT5), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(KEYINPUT84), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n447), .B2(new_n457), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n457), .A2(new_n460), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G57gat), .B(G85gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(G1gat), .B(G29gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n462), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n459), .A2(new_n461), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT6), .B1(new_n474), .B2(new_n471), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n471), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n473), .A2(new_n475), .B1(new_n476), .B2(KEYINPUT6), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n478), .B(new_n386), .C1(new_n391), .C2(new_n392), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n394), .A2(new_n395), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT29), .B1(new_n432), .B2(new_n454), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT29), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT3), .B1(new_n381), .B2(new_n484), .ZN(new_n485));
  OAI221_X1 g284(.A(new_n482), .B1(new_n381), .B2(new_n483), .C1(new_n485), .C2(new_n432), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n481), .B(KEYINPUT81), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n380), .A2(new_n369), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n484), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n432), .B1(new_n489), .B2(new_n454), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n381), .B1(new_n484), .B2(new_n455), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(G22gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n486), .A2(new_n495), .A3(new_n492), .ZN(new_n496));
  XNOR2_X1  g295(.A(G78gat), .B(G106gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT31), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(G50gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n495), .B1(new_n486), .B2(new_n492), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT82), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n486), .A2(KEYINPUT82), .A3(new_n492), .A4(new_n495), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n499), .B(KEYINPUT80), .Z(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n462), .A2(new_n466), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n433), .A2(new_n443), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT83), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n452), .A4(new_n436), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n451), .A2(new_n456), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n446), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT83), .B1(new_n444), .B2(new_n446), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n512), .A2(new_n514), .A3(new_n515), .A4(KEYINPUT39), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n452), .B1(new_n451), .B2(new_n456), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT39), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n472), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT40), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT40), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n509), .A2(new_n472), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n313), .B1(new_n387), .B2(new_n388), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n395), .A3(KEYINPUT30), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n389), .A2(new_n527), .A3(new_n314), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n508), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n480), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT86), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n464), .A2(new_n465), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n472), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n471), .B1(new_n464), .B2(new_n465), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n529), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n508), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n360), .B(new_n434), .ZN(new_n543));
  NAND2_X1  g342(.A1(G227gat), .A2(G233gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT32), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n543), .B2(new_n544), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G43gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G71gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(new_n268), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n360), .A2(new_n434), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n360), .A2(new_n434), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n553), .A2(new_n554), .A3(new_n544), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n551), .B1(new_n555), .B2(new_n546), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT32), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n544), .B1(new_n553), .B2(new_n554), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n544), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  OAI221_X1 g363(.A(new_n544), .B1(new_n562), .B2(new_n561), .C1(new_n553), .C2(new_n554), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n564), .A2(KEYINPUT72), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT72), .B1(new_n564), .B2(new_n565), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n552), .B(new_n559), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT72), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n556), .A2(new_n558), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n545), .B1(new_n548), .B2(new_n551), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT36), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n568), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n542), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n480), .A2(new_n531), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n533), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n568), .A2(new_n572), .ZN(new_n581));
  INV_X1    g380(.A(new_n508), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT35), .B1(new_n583), .B2(new_n541), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n573), .A2(new_n508), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586));
  INV_X1    g385(.A(new_n477), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n529), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n366), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n289), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G127gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n228), .B1(new_n289), .B2(new_n594), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n598), .A2(KEYINPUT95), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(KEYINPUT95), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g403(.A(G155gat), .B(G183gat), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n604), .B(new_n605), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n600), .B2(new_n603), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n593), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(new_n592), .A3(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n277), .A2(new_n287), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n615), .A2(new_n219), .A3(new_n223), .A4(new_n229), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n277), .B(new_n287), .C1(new_n222), .C2(new_n221), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n618));
  NAND3_X1  g417(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n618), .B1(new_n617), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G190gat), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n321), .B(new_n616), .C1(new_n620), .C2(new_n621), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n623), .A2(G218gat), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(G218gat), .B1(new_n623), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT99), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n367), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n623), .A2(G218gat), .A3(new_n624), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n635), .ZN(new_n637));
  OAI211_X1 g436(.A(KEYINPUT99), .B(new_n637), .C1(new_n625), .C2(new_n626), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AND4_X1   g438(.A1(new_n310), .A2(new_n590), .A3(new_n614), .A4(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n540), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT101), .B(G1gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1324gat));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n530), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT16), .B(G8gat), .ZN(new_n647));
  OR3_X1    g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n645), .B(KEYINPUT102), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n649), .B2(new_n647), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n649), .A2(KEYINPUT103), .A3(G8gat), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT103), .B1(new_n649), .B2(G8gat), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n648), .B(new_n650), .C1(new_n651), .C2(new_n652), .ZN(G1325gat));
  AOI21_X1  g452(.A(G15gat), .B1(new_n640), .B2(new_n581), .ZN(new_n654));
  INV_X1    g453(.A(new_n574), .ZN(new_n655));
  INV_X1    g454(.A(new_n576), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(G15gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT104), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n654), .B1(new_n640), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT105), .ZN(G1326gat));
  NAND2_X1  g461(.A1(new_n640), .A2(new_n508), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  AND2_X1   g464(.A1(new_n636), .A2(new_n638), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n480), .A2(new_n578), .A3(new_n531), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n578), .B1(new_n480), .B2(new_n531), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n542), .A2(new_n574), .A3(new_n576), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n584), .A2(new_n588), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n611), .A2(new_n613), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n310), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(G29gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n641), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(KEYINPUT44), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n639), .B1(new_n580), .B2(new_n589), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n674), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n641), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n678), .B1(new_n685), .B2(new_n676), .ZN(G1328gat));
  INV_X1    g485(.A(G36gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n675), .A2(new_n687), .A3(new_n530), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT46), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(new_n530), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n691), .B2(new_n687), .ZN(G1329gat));
  NAND2_X1  g491(.A1(new_n683), .A2(new_n658), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT47), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(G43gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n675), .A2(new_n697), .A3(new_n581), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n696), .B(new_n699), .ZN(G1330gat));
  INV_X1    g499(.A(KEYINPUT48), .ZN(new_n701));
  INV_X1    g500(.A(G50gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n675), .A2(new_n702), .A3(new_n508), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT107), .Z(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n683), .B2(new_n508), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n683), .A2(new_n508), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n508), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(G50gat), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n703), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n675), .A2(KEYINPUT108), .A3(new_n702), .A4(new_n508), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n701), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n711), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n712), .B1(new_n711), .B2(new_n716), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n706), .B1(new_n717), .B2(new_n718), .ZN(G1331gat));
  AOI211_X1 g518(.A(new_n253), .B(new_n673), .C1(new_n636), .C2(new_n638), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n590), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n309), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n641), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g524(.A1(new_n722), .A2(new_n529), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  AND2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n726), .B2(new_n727), .ZN(G1333gat));
  OAI21_X1  g529(.A(G71gat), .B1(new_n722), .B2(new_n657), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n722), .A2(G71gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n573), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g533(.A1(new_n723), .A2(new_n508), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g535(.A1(new_n673), .A2(new_n254), .A3(KEYINPUT111), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n614), .B2(new_n253), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n309), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n679), .B2(new_n682), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n540), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n672), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n680), .A2(KEYINPUT113), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n740), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT51), .A4(new_n740), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n265), .A3(new_n641), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n746), .B1(new_n755), .B2(new_n308), .ZN(G1336gat));
  NOR3_X1   g555(.A1(new_n308), .A2(new_n529), .A3(G92gat), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT113), .B1(new_n590), .B2(new_n666), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n747), .B(new_n639), .C1(new_n580), .C2(new_n589), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(new_n740), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n749), .A3(new_n740), .A4(new_n759), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n757), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n266), .B1(new_n744), .B2(new_n530), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT115), .B1(new_n769), .B2(KEYINPUT52), .ZN(new_n770));
  INV_X1    g569(.A(new_n757), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n758), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(new_n764), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT115), .B(KEYINPUT52), .C1(new_n773), .C2(new_n767), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(new_n754), .B2(new_n757), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n768), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n771), .B1(new_n752), .B2(new_n753), .ZN(new_n779));
  NOR4_X1   g578(.A1(new_n779), .A2(new_n767), .A3(KEYINPUT116), .A4(KEYINPUT52), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n770), .A2(new_n775), .B1(new_n778), .B2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n745), .B2(new_n657), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n754), .A2(new_n268), .A3(new_n581), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n308), .ZN(G1338gat));
  AOI21_X1  g583(.A(new_n269), .B1(new_n744), .B2(new_n508), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n582), .A2(G106gat), .A3(new_n308), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n754), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n786), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n772), .B2(new_n764), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT53), .B1(new_n791), .B2(new_n785), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1339gat));
  NAND4_X1  g592(.A1(new_n288), .A2(new_n293), .A3(KEYINPUT118), .A4(new_n257), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n288), .A2(new_n293), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n295), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n295), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT54), .B(new_n794), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n304), .B1(new_n294), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n801), .A3(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n305), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n799), .B2(new_n801), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT119), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n801), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n808), .A2(new_n809), .A3(new_n305), .A4(new_n802), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n233), .A2(new_n234), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n236), .A2(new_n237), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n248), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n252), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n636), .A2(new_n811), .A3(new_n638), .A4(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n811), .A2(new_n253), .B1(new_n309), .B2(new_n815), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n666), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n818), .A2(new_n673), .B1(new_n308), .B2(new_n720), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n540), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n583), .A2(new_n530), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n254), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(new_n399), .ZN(G1340gat));
  NOR2_X1   g623(.A1(new_n822), .A2(new_n308), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(new_n397), .ZN(G1341gat));
  INV_X1    g625(.A(new_n822), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(G127gat), .A3(new_n614), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(KEYINPUT120), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(KEYINPUT120), .ZN(new_n830));
  AOI21_X1  g629(.A(G127gat), .B1(new_n827), .B2(new_n614), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(G1342gat));
  NOR2_X1   g631(.A1(new_n822), .A2(new_n639), .ZN(new_n833));
  NOR2_X1   g632(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n834));
  AND2_X1   g633(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n833), .B2(new_n834), .ZN(G1343gat));
  NOR4_X1   g636(.A1(new_n666), .A2(new_n309), .A3(new_n253), .A4(new_n673), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n815), .A2(new_n309), .ZN(new_n839));
  XOR2_X1   g638(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n840));
  NAND2_X1  g639(.A1(new_n806), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n253), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n842), .B2(new_n803), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n639), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n614), .B1(new_n844), .B2(new_n816), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n508), .B1(new_n838), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT57), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n811), .A2(new_n253), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n839), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n639), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n614), .B1(new_n851), .B2(new_n816), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n848), .B(new_n508), .C1(new_n852), .C2(new_n838), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n658), .A2(new_n540), .A3(new_n530), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G141gat), .B1(new_n855), .B2(new_n254), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n819), .A2(new_n582), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n854), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n253), .A2(new_n419), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n862), .B(G148gat), .C1(new_n855), .C2(new_n308), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT57), .B1(new_n819), .B2(new_n582), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n803), .A2(new_n804), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n636), .A2(new_n638), .A3(new_n866), .A4(new_n815), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n614), .B1(new_n844), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n848), .B(new_n508), .C1(new_n838), .C2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n865), .A2(new_n309), .A3(new_n854), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G148gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n864), .B1(new_n871), .B2(KEYINPUT59), .ZN(new_n872));
  AOI211_X1 g671(.A(KEYINPUT122), .B(new_n862), .C1(new_n870), .C2(G148gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n863), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n858), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n417), .A3(new_n309), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1345gat));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n427), .A3(new_n614), .ZN(new_n878));
  OAI21_X1  g677(.A(G155gat), .B1(new_n855), .B2(new_n673), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n875), .B2(new_n666), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n855), .A2(new_n428), .A3(new_n639), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n819), .A2(new_n583), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n641), .A2(new_n529), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n253), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n309), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(G176gat), .ZN(new_n892));
  XOR2_X1   g691(.A(KEYINPUT123), .B(G176gat), .Z(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n890), .B2(new_n893), .ZN(G1349gat));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n329), .B1(KEYINPUT124), .B2(G183gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n887), .A2(new_n614), .A3(new_n898), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n886), .A2(new_n673), .B1(KEYINPUT124), .B2(new_n339), .ZN(new_n900));
  AOI211_X1 g699(.A(new_n896), .B(new_n897), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AND4_X1   g700(.A1(KEYINPUT125), .A2(new_n899), .A3(new_n895), .A4(new_n900), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1350gat));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G190gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n886), .A2(new_n639), .ZN(new_n906));
  MUX2_X1   g705(.A(new_n904), .B(new_n905), .S(new_n906), .Z(G1351gat));
  AND2_X1   g706(.A1(new_n865), .A2(new_n869), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n657), .A2(new_n885), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n253), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g709(.A(KEYINPUT126), .B(G197gat), .Z(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n857), .A2(new_n909), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n254), .A2(new_n911), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  NAND4_X1  g714(.A1(new_n857), .A2(new_n302), .A3(new_n309), .A4(new_n909), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT62), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n916), .A2(KEYINPUT62), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n908), .A2(new_n309), .A3(new_n909), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n302), .ZN(G1353gat));
  NOR3_X1   g719(.A1(new_n913), .A2(G211gat), .A3(new_n673), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT127), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n908), .A2(new_n614), .A3(new_n909), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G211gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT63), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n926), .A3(G211gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n922), .A2(new_n925), .A3(new_n927), .ZN(G1354gat));
  NAND4_X1  g727(.A1(new_n908), .A2(G218gat), .A3(new_n666), .A4(new_n909), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n367), .B1(new_n913), .B2(new_n639), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(G1355gat));
endmodule


