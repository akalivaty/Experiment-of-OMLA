//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT82), .ZN(new_n207));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT80), .B1(new_n209), .B2(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(G141gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n219), .B2(KEYINPUT2), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n216), .ZN(new_n222));
  NOR2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G141gat), .B(G148gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n224), .B(KEYINPUT79), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n209), .A2(G141gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n212), .A2(G148gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n229), .B(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT79), .B1(new_n233), .B2(new_n224), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n221), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G113gat), .ZN(new_n236));
  INV_X1    g035(.A(G120gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT1), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G134gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G127gat), .ZN(new_n240));
  INV_X1    g039(.A(G127gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G134gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(KEYINPUT73), .A2(G113gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT73), .A2(G113gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n237), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(G113gat), .B2(G120gat), .ZN(new_n248));
  AND2_X1   g047(.A1(G113gat), .A2(G120gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  OAI22_X1  g050(.A1(new_n243), .A2(new_n246), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n240), .A2(new_n242), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(new_n248), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n244), .A2(new_n245), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G120gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n238), .B1(new_n236), .B2(new_n237), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n254), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n221), .B(new_n259), .C1(new_n228), .C2(new_n234), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n208), .B1(new_n253), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT5), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n207), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n208), .ZN(new_n264));
  INV_X1    g063(.A(new_n260), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT79), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n227), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n259), .B1(new_n269), .B2(new_n221), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n264), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n215), .A2(new_n220), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n268), .B2(new_n227), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT81), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n235), .A2(new_n277), .A3(KEYINPUT3), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n275), .B(new_n221), .C1(new_n228), .C2(new_n234), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .A4(new_n252), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n274), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n282), .A2(new_n283), .A3(new_n208), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n263), .A2(new_n272), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT83), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n282), .A2(new_n287), .A3(new_n283), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n282), .B2(new_n283), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n280), .B(new_n286), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n206), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n284), .A2(new_n280), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n261), .A2(new_n207), .A3(new_n262), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT82), .B1(new_n271), .B2(KEYINPUT5), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(new_n290), .A3(new_n205), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n290), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT6), .A3(new_n206), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G197gat), .B(G204gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT22), .ZN(new_n305));
  INV_X1    g104(.A(G211gat), .ZN(new_n306));
  INV_X1    g105(.A(G218gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n304), .A3(new_n308), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT27), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G183gat), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n323), .B1(new_n321), .B2(new_n322), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n315), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n324), .ZN(new_n329));
  INV_X1    g128(.A(G169gat), .ZN(new_n330));
  INV_X1    g129(.A(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333));
  NAND2_X1  g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n336), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n335), .B2(new_n337), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n327), .A2(new_n329), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n343));
  NOR2_X1   g142(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n332), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n332), .B(KEYINPUT68), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n334), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(KEYINPUT23), .B2(new_n336), .ZN(new_n351));
  NAND2_X1  g150(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n352));
  MUX2_X1   g151(.A(G183gat), .B(new_n352), .S(G190gat), .Z(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT24), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT66), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT66), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n358), .A3(new_n355), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n351), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n362));
  INV_X1    g161(.A(new_n351), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n347), .B2(new_n348), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n355), .A2(KEYINPUT69), .B1(G183gat), .B2(G190gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(KEYINPUT69), .B2(new_n355), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n366), .B2(new_n353), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n361), .A2(new_n362), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G226gat), .ZN(new_n369));
  INV_X1    g168(.A(G233gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n342), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(KEYINPUT29), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n361), .A2(new_n362), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n364), .A2(new_n367), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n327), .A2(new_n329), .A3(new_n341), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n314), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n371), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n312), .A2(new_n313), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n342), .A2(new_n368), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(new_n373), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n381), .B1(new_n383), .B2(new_n373), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT75), .A3(new_n314), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(KEYINPUT37), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(KEYINPUT37), .A3(new_n388), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT38), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n386), .A2(new_n388), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n391), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n379), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT87), .A3(new_n314), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n384), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT38), .B1(new_n404), .B2(KEYINPUT37), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n395), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n303), .A2(new_n398), .A3(new_n400), .A4(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n408));
  NAND2_X1  g207(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT76), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n393), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n391), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n280), .B1(new_n288), .B2(new_n289), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n264), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n253), .A2(new_n260), .A3(new_n208), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT39), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT39), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(new_n421), .A3(new_n264), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n420), .A2(KEYINPUT40), .A3(new_n205), .A4(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n423), .A2(new_n292), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n412), .A2(new_n410), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n420), .A2(new_n205), .A3(new_n422), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT40), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n413), .A2(new_n424), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT85), .B(G22gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n275), .B1(new_n314), .B2(KEYINPUT29), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n235), .ZN(new_n433));
  XNOR2_X1  g232(.A(G78gat), .B(G106gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT29), .B1(new_n274), .B2(new_n275), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n433), .B(new_n435), .C1(new_n382), .C2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n382), .B1(new_n279), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT3), .B1(new_n382), .B2(new_n438), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n274), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n434), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT31), .B(G50gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G228gat), .A2(G233gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(new_n442), .A3(new_n444), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n431), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n448), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n444), .B1(new_n437), .B2(new_n442), .ZN(new_n453));
  OAI211_X1 g252(.A(G228gat), .B(G233gat), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n430), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n407), .A2(new_n429), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n412), .A2(new_n410), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n412), .A2(new_n410), .A3(new_n393), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(new_n409), .ZN(new_n462));
  INV_X1    g261(.A(new_n301), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n299), .A2(KEYINPUT84), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n292), .A2(new_n465), .A3(new_n298), .A4(new_n293), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n457), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n259), .B1(new_n342), .B2(new_n368), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n376), .A2(new_n252), .A3(new_n377), .ZN(new_n470));
  NAND2_X1  g269(.A1(G227gat), .A2(G233gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n471), .B(KEYINPUT64), .Z(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT65), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G15gat), .B(G43gat), .Z(new_n479));
  XNOR2_X1  g278(.A(G71gat), .B(G99gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n481), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n475), .B(KEYINPUT32), .C1(new_n477), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n472), .B1(new_n469), .B2(new_n470), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI211_X1 g287(.A(KEYINPUT34), .B(new_n474), .C1(new_n469), .C2(new_n470), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n485), .B(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n491), .A2(KEYINPUT36), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT74), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n490), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n488), .A2(new_n489), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n485), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(KEYINPUT36), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n459), .A2(new_n468), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n464), .A2(new_n466), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n502), .A2(new_n301), .B1(new_n413), .B2(new_n425), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n485), .A2(new_n493), .A3(new_n496), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n496), .B1(new_n485), .B2(new_n493), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n457), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n413), .A2(new_n425), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n491), .A4(new_n302), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n500), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT14), .B(G29gat), .Z(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(G36gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n520), .B1(new_n517), .B2(KEYINPUT88), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(KEYINPUT88), .B2(new_n517), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n516), .B(new_n521), .C1(KEYINPUT88), .C2(new_n517), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n523), .A2(new_n524), .A3(new_n525), .A4(KEYINPUT17), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  INV_X1    g330(.A(G1gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT16), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n533), .B(new_n534), .C1(new_n532), .C2(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n535), .B(new_n536), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n525), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(KEYINPUT91), .A2(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n540), .B1(new_n537), .B2(new_n530), .ZN(new_n546));
  INV_X1    g345(.A(new_n544), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(new_n542), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n537), .A2(new_n539), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(new_n540), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n545), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(G197gat), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT11), .B(G169gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT12), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n545), .A2(new_n548), .A3(new_n558), .A4(new_n552), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n512), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT41), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT7), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n571), .B1(new_n570), .B2(new_n575), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT97), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n530), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n566), .A2(KEYINPUT41), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n582), .B2(new_n539), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n320), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n577), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n580), .A3(new_n579), .ZN(new_n589));
  INV_X1    g388(.A(new_n581), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n528), .B2(new_n529), .ZN(new_n592));
  OAI21_X1  g391(.A(G190gat), .B1(new_n592), .B2(new_n585), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT96), .B1(new_n594), .B2(new_n307), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(G218gat), .A3(new_n593), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n568), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n320), .B1(new_n583), .B2(new_n586), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n592), .A2(new_n585), .A3(G190gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n307), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND4_X1   g400(.A1(new_n598), .A2(new_n601), .A3(new_n568), .A4(new_n596), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n565), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n598), .A3(new_n596), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n567), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n595), .A2(new_n568), .A3(new_n596), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n564), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G71gat), .A2(G78gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT9), .ZN(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G64gat), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n613), .B2(KEYINPUT94), .ZN(new_n614));
  OR2_X1    g413(.A1(G71gat), .A2(G78gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT95), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n616), .A3(new_n610), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n610), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT95), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n614), .A2(new_n617), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n610), .B(KEYINPUT93), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n622), .B(new_n615), .C1(new_n612), .C2(new_n613), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G127gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n537), .B1(new_n625), .B2(new_n624), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n217), .ZN(new_n633));
  XOR2_X1   g432(.A(G183gat), .B(G211gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n624), .B1(new_n578), .B2(new_n581), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n621), .B(new_n623), .C1(new_n576), .C2(new_n577), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT98), .Z(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT99), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n589), .A2(new_n590), .B1(new_n621), .B2(new_n623), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n576), .A2(new_n577), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n624), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n623), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n591), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n643), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G120gat), .B(G148gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n645), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n645), .B2(new_n654), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n609), .A2(new_n639), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n563), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT6), .B1(new_n300), .B2(new_n206), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n465), .B1(new_n667), .B2(new_n298), .ZN(new_n668));
  INV_X1    g467(.A(new_n466), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n301), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n532), .ZN(G1324gat));
  OR3_X1    g471(.A1(new_n666), .A2(KEYINPUT101), .A3(new_n508), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT101), .B1(new_n666), .B2(new_n508), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(G8gat), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n666), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(KEYINPUT42), .A3(new_n462), .A4(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n673), .B2(new_n674), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n675), .B(new_n678), .C1(new_n680), .C2(KEYINPUT42), .ZN(G1325gat));
  AOI21_X1  g480(.A(G15gat), .B1(new_n676), .B2(new_n491), .ZN(new_n682));
  INV_X1    g481(.A(new_n499), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G15gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT102), .Z(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n676), .B2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n666), .A2(new_n458), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT103), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n639), .A2(new_n662), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n608), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n563), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n670), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n562), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n507), .A2(new_n511), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n506), .A2(new_n670), .A3(new_n508), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT35), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT105), .B1(new_n701), .B2(new_n510), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n500), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n608), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n512), .B2(new_n608), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n697), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n709), .A2(new_n467), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n696), .B1(new_n710), .B2(new_n513), .ZN(G1328gat));
  NOR3_X1   g510(.A1(new_n694), .A2(G36gat), .A3(new_n508), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(KEYINPUT107), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n709), .A2(new_n462), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G36gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n717), .A2(new_n718), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n714), .B(new_n716), .C1(new_n720), .C2(new_n721), .ZN(G1329gat));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  AND4_X1   g523(.A1(new_n724), .A2(new_n563), .A3(new_n491), .A4(new_n693), .ZN(new_n725));
  INV_X1    g524(.A(new_n697), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n459), .A2(new_n499), .A3(new_n468), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n698), .B1(new_n507), .B2(new_n511), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n701), .A2(KEYINPUT105), .A3(new_n510), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n704), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n730), .A2(new_n609), .A3(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n683), .B(new_n726), .C1(new_n732), .C2(new_n707), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n725), .B1(new_n733), .B2(G43gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n723), .B1(new_n734), .B2(KEYINPUT109), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n724), .B1(new_n709), .B2(new_n683), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n736), .B(KEYINPUT47), .C1(new_n737), .C2(new_n725), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n735), .A2(new_n738), .ZN(G1330gat));
  NAND3_X1  g538(.A1(new_n709), .A2(G50gat), .A3(new_n457), .ZN(new_n740));
  INV_X1    g539(.A(G50gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n694), .B2(new_n458), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1331gat));
  INV_X1    g544(.A(new_n562), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n609), .A2(new_n746), .A3(new_n639), .A4(new_n662), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n467), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n462), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT49), .B(G64gat), .Z(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n751), .B2(new_n753), .ZN(G1333gat));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755));
  INV_X1    g554(.A(G71gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n499), .A2(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n748), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n755), .B1(new_n748), .B2(new_n757), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n748), .A2(new_n491), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(G71gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n748), .A2(new_n457), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n639), .A2(new_n562), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n703), .A2(new_n608), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n768), .A2(KEYINPUT112), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n608), .A4(new_n765), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(KEYINPUT112), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n670), .A2(G85gat), .A3(new_n663), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n765), .A2(new_n662), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n705), .B2(new_n708), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(new_n467), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n573), .B2(new_n776), .ZN(G1336gat));
  AOI21_X1  g576(.A(new_n574), .B1(new_n775), .B2(new_n462), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n462), .A2(new_n574), .A3(new_n662), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n768), .B2(new_n770), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT52), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n778), .A2(KEYINPUT52), .ZN(new_n782));
  INV_X1    g581(.A(new_n779), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n769), .A2(new_n771), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n782), .B2(new_n784), .ZN(G1337gat));
  XOR2_X1   g584(.A(KEYINPUT114), .B(G99gat), .Z(new_n786));
  NAND2_X1  g585(.A1(new_n775), .A2(new_n683), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(KEYINPUT113), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(KEYINPUT113), .B2(new_n787), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n491), .A2(new_n662), .A3(new_n786), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n769), .A2(new_n771), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1338gat));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n775), .B2(new_n457), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n458), .A2(new_n663), .A3(G106gat), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n768), .B2(new_n770), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n794), .A2(KEYINPUT53), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n769), .A2(new_n771), .A3(new_n795), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n746), .A2(new_n256), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  INV_X1    g602(.A(new_n643), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n652), .B2(new_n591), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n650), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT10), .B1(new_n640), .B2(new_n641), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n582), .A2(new_n651), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n803), .B(new_n804), .C1(new_n807), .C2(new_n808), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n658), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT55), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n658), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n806), .A2(new_n809), .A3(new_n812), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n812), .B1(new_n806), .B2(new_n809), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n660), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT116), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n659), .B1(new_n814), .B2(new_n819), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(new_n562), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n546), .A2(new_n542), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n551), .A2(new_n540), .A3(new_n550), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n557), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n662), .A2(new_n561), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n609), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n561), .A2(new_n834), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n603), .B2(new_n607), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n824), .A2(new_n830), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n639), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n609), .A2(new_n746), .A3(new_n639), .A4(new_n663), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT117), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n639), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n839), .A2(new_n840), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n608), .B1(new_n831), .B2(new_n835), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n850), .A3(new_n843), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n495), .A2(new_n497), .A3(new_n456), .A4(new_n451), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n462), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n845), .A2(new_n851), .A3(new_n467), .A4(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n802), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n845), .A2(new_n458), .A3(new_n851), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n851), .A3(new_n860), .A4(new_n458), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n462), .A2(new_n670), .ZN(new_n863));
  AND4_X1   g662(.A1(new_n491), .A2(new_n862), .A3(new_n562), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n857), .B1(new_n864), .B2(new_n236), .ZN(G1340gat));
  OAI211_X1 g664(.A(new_n237), .B(new_n662), .C1(new_n855), .C2(new_n856), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n491), .A2(new_n862), .A3(new_n662), .A4(new_n863), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n237), .ZN(G1341gat));
  AND3_X1   g667(.A1(new_n862), .A2(new_n491), .A3(new_n863), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n846), .A2(new_n241), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n854), .B2(new_n846), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n854), .A2(KEYINPUT120), .A3(new_n846), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(G127gat), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n869), .A2(new_n870), .B1(new_n871), .B2(new_n873), .ZN(G1342gat));
  NAND2_X1  g673(.A1(new_n608), .A2(new_n239), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT56), .B1(new_n854), .B2(new_n875), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n854), .A2(KEYINPUT56), .A3(new_n875), .ZN(new_n877));
  AND4_X1   g676(.A1(new_n491), .A2(new_n862), .A3(new_n608), .A4(new_n863), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n876), .B(new_n877), .C1(new_n878), .C2(new_n239), .ZN(G1343gat));
  NAND2_X1  g678(.A1(new_n499), .A2(new_n863), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n845), .A2(new_n457), .A3(new_n851), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n816), .B1(new_n811), .B2(new_n813), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(KEYINPUT55), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n826), .A2(KEYINPUT121), .A3(new_n827), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n562), .A3(new_n887), .A4(new_n825), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(KEYINPUT122), .A3(new_n835), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT122), .B1(new_n888), .B2(new_n835), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n609), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n841), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n843), .B1(new_n892), .B2(new_n639), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n458), .A2(new_n882), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n880), .B1(new_n883), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n212), .B1(new_n896), .B2(new_n562), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n845), .A2(new_n467), .A3(new_n851), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n683), .A2(new_n462), .A3(new_n458), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n898), .A2(new_n212), .A3(new_n562), .A4(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT58), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n881), .A2(new_n882), .B1(new_n893), .B2(new_n894), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n746), .A3(new_n880), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n900), .B(new_n903), .C1(new_n905), .C2(new_n212), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n902), .A2(new_n906), .ZN(G1344gat));
  NAND2_X1  g706(.A1(new_n898), .A2(new_n899), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT59), .B1(new_n908), .B2(new_n663), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n209), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n911), .A3(new_n662), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n839), .A2(new_n825), .A3(new_n828), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n891), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n844), .B1(new_n914), .B2(new_n846), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n882), .B1(new_n915), .B2(new_n458), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n845), .A2(new_n851), .A3(new_n894), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n663), .B(new_n880), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n910), .B(new_n912), .C1(new_n918), .C2(new_n919), .ZN(G1345gat));
  AOI21_X1  g719(.A(new_n217), .B1(new_n896), .B2(new_n639), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n898), .A2(new_n217), .A3(new_n639), .A4(new_n899), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT123), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n904), .A2(new_n846), .A3(new_n880), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n922), .B(new_n925), .C1(new_n926), .C2(new_n217), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n927), .ZN(G1346gat));
  NOR2_X1   g727(.A1(new_n609), .A2(new_n218), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n898), .A2(new_n608), .A3(new_n899), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n896), .A2(new_n929), .B1(new_n930), .B2(new_n218), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n508), .A2(new_n852), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n845), .A2(new_n851), .A3(new_n670), .A4(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n562), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n508), .A2(new_n467), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n491), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n859), .B2(new_n861), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n746), .A2(new_n330), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  AOI21_X1  g739(.A(new_n331), .B1(new_n938), .B2(new_n662), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n933), .A2(G176gat), .A3(new_n663), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT124), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n942), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n945));
  AOI211_X1 g744(.A(new_n663), .B(new_n937), .C1(new_n859), .C2(new_n861), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n331), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n947), .ZN(G1349gat));
  AOI21_X1  g747(.A(new_n316), .B1(new_n938), .B2(new_n639), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n845), .A2(new_n670), .A3(new_n851), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n317), .A2(new_n319), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n639), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n950), .A2(new_n951), .A3(new_n932), .A4(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT125), .B1(new_n933), .B2(new_n953), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT60), .B1(new_n949), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n955), .A2(new_n956), .ZN(new_n960));
  AOI211_X1 g759(.A(new_n846), .B(new_n937), .C1(new_n859), .C2(new_n861), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n316), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n958), .A2(new_n962), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n934), .A2(new_n320), .A3(new_n608), .ZN(new_n964));
  AOI211_X1 g763(.A(KEYINPUT61), .B(new_n320), .C1(new_n938), .C2(new_n608), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  INV_X1    g765(.A(new_n937), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n862), .A2(new_n608), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n968), .B2(G190gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n964), .B1(new_n965), .B2(new_n969), .ZN(G1351gat));
  INV_X1    g769(.A(new_n950), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n499), .A2(new_n462), .A3(new_n457), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n562), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n499), .A2(new_n936), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n916), .B2(new_n917), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n562), .A2(G197gat), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1352gat));
  INV_X1    g777(.A(G204gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n973), .A2(new_n979), .A3(new_n662), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n973), .A2(new_n982), .A3(new_n979), .A4(new_n662), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n976), .A2(new_n662), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n981), .B(new_n983), .C1(new_n984), .C2(new_n979), .ZN(G1353gat));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT63), .ZN(new_n987));
  AOI211_X1 g786(.A(new_n846), .B(new_n975), .C1(new_n916), .C2(new_n917), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n986), .B(new_n987), .C1(new_n988), .C2(new_n306), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n306), .A3(new_n639), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n306), .B1(new_n976), .B2(new_n639), .ZN(new_n991));
  OAI21_X1  g790(.A(KEYINPUT126), .B1(new_n991), .B2(KEYINPUT63), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n988), .A2(new_n987), .A3(new_n306), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n989), .B(new_n990), .C1(new_n992), .C2(new_n993), .ZN(G1354gat));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n976), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(new_n608), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n976), .A2(new_n995), .ZN(new_n998));
  OAI21_X1  g797(.A(G218gat), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n973), .A2(new_n307), .A3(new_n608), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1355gat));
endmodule


