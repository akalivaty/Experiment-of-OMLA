//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(KEYINPUT75), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(G125), .A3(G140), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(KEYINPUT16), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n191), .B2(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n195), .A2(new_n200), .A3(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT69), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n212), .A3(G119), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n203), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n205), .A2(new_n207), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT23), .B1(new_n215), .B2(new_n209), .ZN(new_n216));
  OAI21_X1  g030(.A(G110), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n213), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT24), .B(G110), .ZN(new_n219));
  OR2_X1    g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n202), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT76), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n202), .A2(new_n217), .A3(KEYINPUT76), .A4(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G125), .B(G140), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n200), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n228));
  INV_X1    g042(.A(G110), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT69), .B(G119), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n203), .B1(new_n230), .B2(G128), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n228), .A2(KEYINPUT77), .A3(new_n229), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n218), .A2(new_n219), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n214), .A2(new_n216), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT77), .B1(new_n235), .B2(new_n229), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n199), .B(new_n227), .C1(new_n234), .C2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G137), .ZN(new_n238));
  INV_X1    g052(.A(G953), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n239), .A2(G221), .A3(G234), .ZN(new_n240));
  XOR2_X1   g054(.A(new_n238), .B(new_n240), .Z(new_n241));
  AND3_X1   g055(.A1(new_n225), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n225), .B2(new_n237), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT25), .B1(new_n244), .B2(new_n188), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n225), .A2(new_n237), .ZN(new_n246));
  INV_X1    g060(.A(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n225), .A2(new_n237), .A3(new_n241), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n189), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n248), .A2(new_n188), .A3(new_n249), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n250), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT78), .A3(new_n189), .ZN(new_n259));
  INV_X1    g073(.A(new_n189), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n188), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT79), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n244), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n254), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n205), .A2(new_n207), .A3(G116), .ZN(new_n265));
  INV_X1    g079(.A(G116), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G119), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G113), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT2), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G113), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n265), .A2(new_n267), .A3(new_n273), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n268), .A2(KEYINPUT70), .A3(new_n274), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G137), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT65), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G137), .ZN(new_n285));
  AND2_X1   g099(.A1(KEYINPUT11), .A2(G134), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(G134), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT11), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT66), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n283), .A2(new_n285), .A3(new_n286), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G134), .ZN(new_n294));
  AOI21_X1  g108(.A(G131), .B1(new_n294), .B2(G137), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n288), .A2(new_n291), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n200), .A2(G143), .ZN(new_n297));
  INV_X1    g111(.A(G143), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G146), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n297), .A2(new_n299), .A3(new_n300), .A4(G128), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT64), .B1(new_n298), .B2(G146), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n200), .A3(G143), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n302), .A2(new_n304), .A3(new_n299), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n210), .A2(new_n212), .B1(new_n297), .B2(KEYINPUT1), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT65), .B(G137), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n289), .B1(new_n308), .B2(G134), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G131), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n296), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n288), .A2(new_n291), .A3(new_n293), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n294), .A2(G137), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n288), .A2(new_n291), .A3(new_n293), .A4(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n312), .A2(new_n295), .B1(new_n314), .B2(G131), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n302), .A2(new_n304), .A3(new_n299), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT0), .A2(G128), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT0), .A2(G128), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n297), .A2(new_n299), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n316), .A2(new_n319), .B1(new_n320), .B2(new_n317), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT30), .B(new_n311), .C1(new_n315), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n311), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT1), .B1(new_n298), .B2(G146), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n211), .A2(G128), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n316), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n330), .A2(new_n301), .B1(new_n309), .B2(G131), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT68), .A3(new_n296), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n314), .A2(G131), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n296), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n325), .A2(new_n332), .B1(new_n334), .B2(new_n321), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n281), .B(new_n323), .C1(new_n335), .C2(KEYINPUT30), .ZN(new_n336));
  INV_X1    g150(.A(G237), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n239), .A3(G210), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n338), .B(KEYINPUT27), .Z(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G101), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n339), .B(new_n340), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n321), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n311), .A3(new_n280), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT31), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n336), .A2(KEYINPUT31), .A3(new_n341), .A4(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n325), .A2(new_n332), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n280), .B1(new_n349), .B2(new_n342), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n322), .B1(new_n333), .B2(new_n296), .ZN(new_n351));
  INV_X1    g165(.A(new_n311), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n281), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(KEYINPUT71), .B(KEYINPUT28), .C1(new_n350), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n341), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n356));
  AND4_X1   g170(.A1(KEYINPUT68), .A2(new_n296), .A3(new_n307), .A4(new_n310), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT68), .B1(new_n331), .B2(new_n296), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n357), .A2(new_n358), .B1(new_n315), .B2(new_n322), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n281), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n356), .B1(new_n360), .B2(new_n343), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n343), .A2(new_n356), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n354), .B(new_n355), .C1(new_n361), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n348), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(KEYINPUT32), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n348), .B2(new_n365), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n281), .B1(new_n351), .B2(new_n352), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n343), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(KEYINPUT74), .B(new_n281), .C1(new_n351), .C2(new_n352), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(KEYINPUT28), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n362), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n341), .A2(KEYINPUT29), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n188), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n336), .A2(new_n343), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(new_n355), .ZN(new_n383));
  AOI211_X1 g197(.A(KEYINPUT73), .B(new_n341), .C1(new_n336), .C2(new_n343), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n354), .B1(new_n361), .B2(new_n364), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT29), .B1(new_n386), .B2(new_n341), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n380), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G472), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n264), .B1(new_n372), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G469), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G101), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n395), .A2(new_n398), .A3(new_n402), .A4(new_n399), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n405), .A3(G101), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n321), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n394), .A2(G107), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n397), .A2(G104), .ZN(new_n409));
  OAI21_X1  g223(.A(G101), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n307), .A2(new_n411), .A3(KEYINPUT10), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  INV_X1    g229(.A(new_n301), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n326), .A2(G128), .B1(new_n297), .B2(new_n299), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n403), .A2(new_n410), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n418), .A2(KEYINPUT80), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n209), .B1(new_n297), .B2(KEYINPUT1), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n301), .B1(new_n320), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n411), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n415), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n414), .A2(new_n425), .A3(new_n315), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n239), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n419), .A2(new_n330), .A3(new_n301), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n420), .B2(new_n424), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n334), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n334), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT12), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n436), .A2(KEYINPUT82), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n433), .A2(new_n440), .A3(new_n334), .A4(new_n435), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n431), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n414), .A2(new_n425), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT80), .B1(new_n418), .B2(new_n419), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n411), .A2(new_n421), .A3(new_n423), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT10), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT83), .B1(new_n447), .B2(new_n413), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n448), .A3(new_n334), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n430), .B1(new_n449), .B2(new_n426), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n393), .B(new_n188), .C1(new_n442), .C2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n430), .A3(new_n426), .ZN(new_n452));
  INV_X1    g266(.A(new_n426), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n439), .B2(new_n441), .ZN(new_n454));
  OAI211_X1 g268(.A(G469), .B(new_n452), .C1(new_n454), .C2(new_n430), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n393), .A2(new_n188), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G221), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT9), .B(G234), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n461), .B2(new_n188), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT84), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n458), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n278), .A2(new_n279), .A3(new_n406), .A4(new_n404), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n411), .A2(new_n277), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT85), .B(KEYINPUT5), .Z(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n265), .A3(new_n267), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n230), .A2(new_n477), .A3(G116), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G113), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT86), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n265), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n269), .B1(new_n481), .B2(new_n477), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n475), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n473), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n470), .B1(new_n472), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n473), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n482), .B2(new_n475), .ZN(new_n488));
  AND4_X1   g302(.A1(new_n483), .A2(new_n475), .A3(G113), .A4(new_n478), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n471), .A3(new_n469), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n486), .A2(KEYINPUT6), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n322), .A2(G125), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n330), .A2(new_n191), .A3(new_n301), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G224), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G953), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n495), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n490), .A2(new_n471), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n469), .A2(KEYINPUT6), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n492), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT7), .B1(new_n496), .B2(G953), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT7), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n493), .A2(new_n494), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n494), .B(new_n508), .C1(new_n191), .C2(new_n321), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n505), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n472), .A2(new_n485), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n469), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n469), .B(KEYINPUT8), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n480), .A2(new_n484), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n411), .B1(new_n516), .B2(new_n277), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n265), .A2(KEYINPUT5), .A3(new_n267), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n473), .B1(new_n482), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(G902), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n504), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G210), .B1(G237), .B2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n504), .A2(new_n521), .A3(new_n523), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G214), .B1(G237), .B2(G902), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n337), .A2(new_n239), .A3(G214), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n298), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT18), .A3(G131), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n192), .A2(G146), .A3(new_n194), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n227), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n530), .B(G143), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT18), .A2(G131), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(G131), .ZN(new_n539));
  INV_X1    g353(.A(G131), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n201), .B(new_n199), .C1(new_n539), .C2(new_n542), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(G113), .B(G122), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(new_n394), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT19), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n226), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n192), .A2(KEYINPUT19), .A3(new_n194), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n200), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT89), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n539), .A2(new_n541), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n199), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n547), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n538), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT20), .ZN(new_n560));
  NOR2_X1   g374(.A1(G475), .A2(G902), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n548), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n545), .A2(new_n547), .B1(new_n556), .B2(new_n558), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n565), .A2(KEYINPUT90), .A3(new_n560), .A4(new_n561), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n548), .A2(new_n559), .A3(new_n561), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT20), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n547), .A2(KEYINPUT91), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n545), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n188), .B1(new_n545), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g386(.A(G475), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G478), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(KEYINPUT15), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n460), .A2(new_n187), .A3(G953), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G122), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G116), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n266), .A2(G122), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G107), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n210), .A2(new_n212), .A3(G143), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n298), .A2(G128), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n298), .A2(KEYINPUT13), .A3(G128), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G134), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n585), .A2(new_n294), .A3(new_n586), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n584), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n581), .A2(KEYINPUT14), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n583), .A2(new_n594), .A3(G107), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n581), .B(new_n582), .C1(KEYINPUT14), .C2(new_n397), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n585), .A2(new_n586), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G134), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n597), .B1(new_n599), .B2(new_n592), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n579), .B1(new_n593), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n584), .A2(new_n591), .A3(new_n592), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n599), .A2(new_n592), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n602), .B(new_n578), .C1(new_n603), .C2(new_n597), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT92), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(KEYINPUT92), .B(new_n579), .C1(new_n593), .C2(new_n600), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n188), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT93), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT93), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n606), .A2(new_n610), .A3(new_n188), .A4(new_n607), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n577), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n576), .B1(new_n608), .B2(KEYINPUT93), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n239), .A2(G952), .ZN(new_n615));
  NAND2_X1  g429(.A1(G234), .A2(G237), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT21), .B(G898), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(G902), .A3(G953), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT94), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n574), .A2(new_n614), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n529), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n392), .A2(new_n468), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  NAND3_X1  g440(.A1(new_n254), .A2(new_n259), .A3(new_n263), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n366), .A2(new_n367), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n348), .B2(new_n365), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n628), .B1(new_n389), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT97), .B(G478), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n608), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT33), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n634), .A2(KEYINPUT96), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(KEYINPUT96), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n606), .A2(new_n607), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(KEYINPUT33), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n188), .A2(G478), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n633), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n569), .A2(new_n573), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n525), .A2(new_n643), .A3(new_n526), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n504), .A2(new_n521), .A3(KEYINPUT95), .A4(new_n523), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n645), .A2(new_n528), .ZN(new_n646));
  AND4_X1   g460(.A1(new_n622), .A2(new_n642), .A3(new_n644), .A4(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n631), .A2(new_n468), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT98), .Z(new_n649));
  XOR2_X1   g463(.A(KEYINPUT34), .B(G104), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NAND2_X1  g465(.A1(new_n568), .A2(new_n562), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n573), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n614), .A2(new_n653), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n622), .A2(new_n644), .A3(new_n654), .A4(new_n646), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n631), .A2(new_n468), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(new_n630), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n246), .B1(KEYINPUT36), .B2(new_n247), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n247), .A2(KEYINPUT36), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n225), .A2(new_n237), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT99), .B1(new_n663), .B2(new_n262), .ZN(new_n664));
  AND4_X1   g478(.A1(KEYINPUT99), .A2(new_n660), .A3(new_n262), .A4(new_n662), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n254), .A2(new_n259), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n458), .A2(new_n466), .A3(new_n463), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n466), .B1(new_n458), .B2(new_n463), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n624), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT37), .B(G110), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT100), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n672), .B(new_n674), .ZN(G12));
  NAND2_X1  g489(.A1(new_n644), .A2(new_n646), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT78), .B1(new_n258), .B2(new_n189), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n253), .B(new_n260), .C1(new_n257), .C2(new_n250), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n676), .B1(new_n679), .B2(new_n666), .ZN(new_n680));
  OAI221_X1 g494(.A(new_n368), .B1(new_n370), .B2(new_n371), .C1(new_n388), .C2(new_n389), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n617), .B(KEYINPUT102), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n683), .A2(KEYINPUT101), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(KEYINPUT101), .ZN(new_n685));
  OR3_X1    g499(.A1(new_n620), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n614), .A2(new_n653), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n468), .A2(new_n680), .A3(new_n681), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XNOR2_X1  g505(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n527), .B(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n612), .ZN(new_n695));
  INV_X1    g509(.A(new_n613), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n695), .A2(new_n696), .B1(new_n569), .B2(new_n573), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n694), .A2(new_n528), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n382), .A2(new_n341), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n188), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n341), .B1(new_n375), .B2(new_n376), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n368), .B(new_n702), .C1(new_n370), .C2(new_n371), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n698), .A2(new_n667), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n687), .B(KEYINPUT39), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n468), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  NAND2_X1  g525(.A1(new_n640), .A2(new_n641), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n688), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n468), .A2(new_n680), .A3(new_n681), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  OAI21_X1  g529(.A(new_n188), .B1(new_n442), .B2(new_n450), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n717), .A2(new_n463), .A3(new_n451), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n681), .A2(new_n264), .A3(new_n647), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n681), .A2(new_n264), .A3(new_n655), .A4(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NAND3_X1  g537(.A1(new_n717), .A2(new_n463), .A3(new_n451), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n623), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n680), .A2(new_n681), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NOR2_X1   g541(.A1(new_n629), .A2(new_n389), .ZN(new_n728));
  XOR2_X1   g542(.A(new_n367), .B(KEYINPUT104), .Z(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n378), .A2(KEYINPUT105), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n377), .A2(new_n732), .A3(new_n362), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n355), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n730), .B1(new_n734), .B2(new_n348), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n644), .A2(new_n646), .A3(new_n697), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n622), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n724), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(new_n264), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NOR2_X1   g556(.A1(new_n676), .A2(new_n724), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n736), .A2(new_n743), .A3(new_n667), .A4(new_n713), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  AND3_X1   g559(.A1(new_n504), .A2(new_n521), .A3(new_n523), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n523), .B1(new_n504), .B2(new_n521), .ZN(new_n747));
  INV_X1    g561(.A(new_n528), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n746), .A2(new_n747), .A3(new_n462), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n458), .A2(KEYINPUT106), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n451), .A2(new_n455), .A3(new_n751), .A4(new_n457), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n681), .A3(new_n264), .A4(new_n713), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n713), .A2(new_n749), .A3(new_n750), .A4(new_n752), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n370), .A2(KEYINPUT32), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n758), .B(new_n368), .C1(new_n389), .C2(new_n388), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n759), .A3(KEYINPUT42), .A4(new_n264), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND4_X1  g576(.A1(new_n753), .A2(new_n681), .A3(new_n264), .A4(new_n689), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT107), .B(G134), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G36));
  NAND2_X1  g579(.A1(new_n574), .A2(new_n640), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT43), .Z(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n630), .A3(new_n667), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT44), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n527), .A2(new_n748), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT108), .Z(new_n771));
  AND2_X1   g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n452), .B1(new_n454), .B2(new_n430), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n393), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n774), .B2(new_n773), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT46), .B1(new_n776), .B2(new_n457), .ZN(new_n777));
  INV_X1    g591(.A(new_n451), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n457), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n462), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n706), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  XNOR2_X1  g598(.A(new_n781), .B(KEYINPUT47), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n372), .A2(new_n390), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n627), .A2(new_n713), .A3(new_n770), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NAND2_X1  g603(.A1(new_n463), .A2(new_n528), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n694), .A2(new_n766), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n717), .A2(new_n451), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT49), .Z(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n264), .A3(new_n704), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  INV_X1    g609(.A(new_n682), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n767), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n627), .A2(new_n728), .A3(new_n735), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n799), .A2(new_n528), .A3(new_n694), .A4(new_n724), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT50), .Z(new_n801));
  NAND2_X1  g615(.A1(new_n718), .A2(new_n770), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n703), .A2(new_n802), .A3(new_n627), .A4(new_n617), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n640), .A2(new_n641), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n797), .A2(new_n718), .A3(new_n770), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n366), .A2(new_n188), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(G472), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n734), .A2(new_n348), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n729), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n667), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n805), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n801), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(KEYINPUT114), .ZN(new_n814));
  INV_X1    g628(.A(new_n799), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n792), .A2(new_n463), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n771), .B(new_n815), .C1(new_n785), .C2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n813), .B2(KEYINPUT114), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n795), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n645), .A2(new_n528), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n746), .A2(new_n747), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n820), .B1(new_n821), .B2(new_n643), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n718), .A3(new_n713), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n811), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n667), .A2(new_n822), .A3(new_n689), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n786), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n826), .B2(new_n468), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n687), .A2(new_n463), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n667), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n750), .A2(new_n752), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n703), .A3(new_n738), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n827), .A2(new_n828), .A3(new_n714), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n690), .A2(new_n714), .A3(new_n744), .A4(new_n832), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n671), .B1(new_n391), .B2(new_n668), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n527), .A2(new_n528), .A3(new_n622), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT109), .B1(new_n612), .B2(new_n613), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n612), .A2(KEYINPUT109), .A3(new_n613), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n574), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n837), .B1(new_n841), .B2(new_n712), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n631), .A2(new_n468), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n836), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n833), .A2(new_n835), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n719), .A2(new_n722), .A3(new_n726), .A4(new_n741), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n725), .A2(new_n822), .A3(new_n667), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n737), .A2(new_n739), .A3(new_n724), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n850), .A2(new_n681), .B1(new_n798), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT113), .A3(new_n719), .A4(new_n722), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n653), .A2(new_n688), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n821), .A2(new_n528), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n840), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n838), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n468), .A2(new_n681), .A3(new_n667), .A4(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n753), .A2(new_n667), .A3(new_n713), .A4(new_n736), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n763), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n849), .A2(new_n853), .A3(new_n761), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n846), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n714), .A2(new_n832), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n828), .B1(new_n865), .B2(new_n827), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n719), .A2(new_n722), .A3(new_n726), .A4(new_n741), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n836), .A2(new_n843), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n761), .A2(new_n869), .A3(new_n861), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT111), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI211_X1 g687(.A(KEYINPUT54), .B(new_n863), .C1(new_n873), .C2(new_n844), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n833), .A2(new_n835), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n761), .A2(new_n869), .A3(new_n861), .A4(new_n870), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n844), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT110), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT110), .B(new_n844), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n871), .A2(new_n872), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT112), .A3(KEYINPUT53), .A4(new_n868), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n868), .A2(KEYINPUT53), .A3(new_n871), .A4(new_n872), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT112), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n874), .B1(new_n887), .B2(KEYINPUT54), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n806), .B1(new_n889), .B2(KEYINPUT48), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n264), .A3(new_n759), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n889), .A2(KEYINPUT48), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n891), .B(new_n892), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n815), .A2(new_n743), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n803), .A2(new_n642), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n615), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n893), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n801), .A2(new_n795), .A3(new_n812), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(new_n817), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n819), .A2(new_n888), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(G952), .A2(G953), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n794), .B1(new_n903), .B2(new_n904), .ZN(G75));
  AOI21_X1  g719(.A(new_n863), .B1(new_n873), .B2(new_n844), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(new_n188), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT56), .B1(new_n907), .B2(G210), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n492), .B1(new_n502), .B2(new_n503), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n498), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT55), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n908), .A2(new_n911), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n239), .A2(G952), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G51));
  XOR2_X1   g729(.A(new_n906), .B(KEYINPUT54), .Z(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n456), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n450), .B2(new_n442), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n906), .A2(new_n188), .A3(new_n776), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(G54));
  INV_X1    g736(.A(KEYINPUT58), .ZN(new_n923));
  INV_X1    g737(.A(G475), .ZN(new_n924));
  OR3_X1    g738(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT118), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT118), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n907), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n565), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n914), .ZN(G60));
  XNOR2_X1  g745(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n638), .B1(new_n888), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n638), .C1(new_n888), .C2(new_n934), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n638), .A2(new_n934), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n914), .B1(new_n916), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n936), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n936), .A2(KEYINPUT121), .A3(new_n938), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT53), .B1(new_n882), .B2(new_n868), .ZN(new_n949));
  OAI211_X1 g763(.A(KEYINPUT122), .B(new_n948), .C1(new_n949), .C2(new_n863), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n906), .B2(new_n947), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n244), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n914), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n953), .A2(KEYINPUT123), .A3(new_n663), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT123), .B1(new_n953), .B2(new_n663), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n955), .B(KEYINPUT61), .C1(new_n957), .C2(new_n956), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G66));
  OAI21_X1  g776(.A(G953), .B1(new_n618), .B2(new_n496), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n847), .A2(new_n843), .A3(new_n836), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(G953), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n909), .B1(G898), .B2(new_n239), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT124), .Z(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  AND2_X1   g782(.A1(new_n827), .A2(new_n714), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n782), .A2(new_n264), .A3(new_n738), .A4(new_n759), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n783), .A2(new_n788), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n761), .A2(new_n763), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(new_n239), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n323), .B1(new_n335), .B2(KEYINPUT30), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n550), .A2(new_n551), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n974), .B(new_n977), .C1(new_n683), .C2(new_n239), .ZN(new_n978));
  INV_X1    g792(.A(new_n707), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n841), .A2(new_n712), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n392), .A2(new_n770), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  AOI22_X1  g796(.A1(new_n772), .A2(new_n782), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(new_n788), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n969), .A2(new_n710), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n984), .A2(KEYINPUT125), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n983), .A2(new_n986), .A3(new_n788), .A4(new_n987), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(G953), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n978), .B1(new_n992), .B2(new_n977), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n978), .B(new_n995), .C1(new_n992), .C2(new_n977), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n239), .B1(G227), .B2(G900), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n994), .A2(new_n998), .A3(new_n996), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(G72));
  NAND3_X1  g816(.A1(new_n988), .A2(new_n991), .A3(new_n964), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  AOI21_X1  g819(.A(new_n699), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1005), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n971), .A2(new_n973), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n964), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n336), .A2(new_n355), .A3(new_n343), .ZN(new_n1010));
  OAI22_X1  g824(.A1(new_n1009), .A2(new_n1010), .B1(G952), .B2(new_n239), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1007), .B1(new_n385), .B2(new_n344), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n1006), .B(new_n1011), .C1(new_n887), .C2(new_n1012), .ZN(G57));
endmodule


