

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n310) );
  XOR2_X1 U325 ( .A(G120GAT), .B(G71GAT), .Z(n417) );
  XNOR2_X1 U326 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U327 ( .A(n426), .B(n425), .ZN(n428) );
  AND2_X1 U328 ( .A1(n522), .A2(n475), .ZN(n476) );
  XNOR2_X1 U329 ( .A(KEYINPUT37), .B(KEYINPUT108), .ZN(n449) );
  XNOR2_X1 U330 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U331 ( .A(KEYINPUT65), .B(n476), .Z(n572) );
  XNOR2_X1 U332 ( .A(n450), .B(n449), .ZN(n520) );
  XNOR2_X1 U333 ( .A(n432), .B(n431), .ZN(n496) );
  XOR2_X1 U334 ( .A(n461), .B(KEYINPUT41), .Z(n539) );
  XNOR2_X1 U335 ( .A(n452), .B(n451), .ZN(n509) );
  XNOR2_X1 U336 ( .A(n481), .B(G176GAT), .ZN(n482) );
  XNOR2_X1 U337 ( .A(n453), .B(G29GAT), .ZN(n454) );
  XNOR2_X1 U338 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  XNOR2_X1 U339 ( .A(n455), .B(n454), .ZN(G1328GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT72), .B(KEYINPUT69), .Z(n293) );
  XOR2_X1 U341 ( .A(G169GAT), .B(G8GAT), .Z(n410) );
  XOR2_X1 U342 ( .A(G15GAT), .B(G1GAT), .Z(n331) );
  XNOR2_X1 U343 ( .A(n410), .B(n331), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U345 ( .A(n294), .B(G113GAT), .Z(n299) );
  XOR2_X1 U346 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n296) );
  XNOR2_X1 U347 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n297), .B(G197GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U351 ( .A(KEYINPUT67), .B(KEYINPUT71), .Z(n301) );
  NAND2_X1 U352 ( .A1(G229GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U354 ( .A(n303), .B(n302), .Z(n309) );
  XNOR2_X1 U355 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n304), .B(G29GAT), .ZN(n305) );
  XOR2_X1 U357 ( .A(n305), .B(KEYINPUT8), .Z(n307) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(G50GAT), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n358) );
  XOR2_X1 U360 ( .A(G141GAT), .B(G22GAT), .Z(n370) );
  XNOR2_X1 U361 ( .A(n358), .B(n370), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n573) );
  XNOR2_X1 U363 ( .A(n573), .B(KEYINPUT73), .ZN(n561) );
  INV_X1 U364 ( .A(n561), .ZN(n468) );
  XNOR2_X1 U365 ( .A(n310), .B(KEYINPUT13), .ZN(n334) );
  XOR2_X1 U366 ( .A(n334), .B(KEYINPUT31), .Z(n312) );
  XNOR2_X1 U367 ( .A(n417), .B(KEYINPUT32), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n318) );
  XNOR2_X1 U369 ( .A(G176GAT), .B(G64GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n313), .B(KEYINPUT79), .ZN(n411) );
  INV_X1 U371 ( .A(KEYINPUT33), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n411), .B(n314), .ZN(n316) );
  NAND2_X1 U373 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U375 ( .A(n318), .B(n317), .Z(n327) );
  XNOR2_X1 U376 ( .A(G148GAT), .B(KEYINPUT75), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n319), .B(KEYINPUT76), .ZN(n320) );
  XOR2_X1 U378 ( .A(n320), .B(G204GAT), .Z(n322) );
  XNOR2_X1 U379 ( .A(G78GAT), .B(G106GAT), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n374) );
  XOR2_X1 U381 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n324) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G92GAT), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U384 ( .A(G85GAT), .B(n325), .Z(n357) );
  XNOR2_X1 U385 ( .A(n374), .B(n357), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n456) );
  INV_X1 U387 ( .A(n456), .ZN(n458) );
  INV_X1 U388 ( .A(n458), .ZN(n578) );
  NOR2_X1 U389 ( .A1(n468), .A2(n578), .ZN(n488) );
  XOR2_X1 U390 ( .A(G155GAT), .B(G78GAT), .Z(n329) );
  XNOR2_X1 U391 ( .A(G127GAT), .B(G71GAT), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U393 ( .A(n330), .B(G211GAT), .Z(n333) );
  XNOR2_X1 U394 ( .A(G22GAT), .B(n331), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n339) );
  BUF_X1 U396 ( .A(n334), .Z(n335) );
  XOR2_X1 U397 ( .A(n335), .B(KEYINPUT12), .Z(n337) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U400 ( .A(n339), .B(n338), .Z(n347) );
  XOR2_X1 U401 ( .A(KEYINPUT84), .B(G64GAT), .Z(n341) );
  XNOR2_X1 U402 ( .A(G8GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U404 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n343) );
  XNOR2_X1 U405 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U408 ( .A(n347), .B(n346), .Z(n583) );
  INV_X1 U409 ( .A(n583), .ZN(n555) );
  XOR2_X1 U410 ( .A(G190GAT), .B(G134GAT), .Z(n418) );
  XOR2_X1 U411 ( .A(KEYINPUT80), .B(G162GAT), .Z(n349) );
  XNOR2_X1 U412 ( .A(G106GAT), .B(G218GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U414 ( .A(n418), .B(n350), .Z(n352) );
  NAND2_X1 U415 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U417 ( .A(KEYINPUT9), .B(KEYINPUT81), .Z(n354) );
  XNOR2_X1 U418 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U420 ( .A(n356), .B(n355), .Z(n360) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U422 ( .A(n360), .B(n359), .Z(n559) );
  XNOR2_X1 U423 ( .A(KEYINPUT36), .B(n559), .ZN(n588) );
  XOR2_X1 U424 ( .A(KEYINPUT92), .B(KEYINPUT23), .Z(n362) );
  XNOR2_X1 U425 ( .A(G50GAT), .B(KEYINPUT93), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U427 ( .A(KEYINPUT91), .B(G162GAT), .Z(n364) );
  XNOR2_X1 U428 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U430 ( .A(KEYINPUT3), .B(n365), .Z(n391) );
  XOR2_X1 U431 ( .A(n366), .B(n391), .Z(n372) );
  XOR2_X1 U432 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n368) );
  NAND2_X1 U433 ( .A1(G228GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U438 ( .A(KEYINPUT21), .B(G218GAT), .Z(n376) );
  XNOR2_X1 U439 ( .A(KEYINPUT90), .B(G211GAT), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U441 ( .A(G197GAT), .B(n377), .Z(n405) );
  XOR2_X1 U442 ( .A(n378), .B(n405), .Z(n477) );
  XOR2_X1 U443 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n379) );
  XOR2_X1 U444 ( .A(n477), .B(n379), .Z(n528) );
  INV_X1 U445 ( .A(n528), .ZN(n533) );
  XOR2_X1 U446 ( .A(G85GAT), .B(G148GAT), .Z(n381) );
  XNOR2_X1 U447 ( .A(G141GAT), .B(G120GAT), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U449 ( .A(G29GAT), .B(G134GAT), .Z(n382) );
  XNOR2_X1 U450 ( .A(n383), .B(n382), .ZN(n397) );
  XOR2_X1 U451 ( .A(KEYINPUT96), .B(KEYINPUT1), .Z(n385) );
  XNOR2_X1 U452 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U454 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n387) );
  XNOR2_X1 U455 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n389), .B(n388), .ZN(n395) );
  XOR2_X1 U458 ( .A(KEYINPUT97), .B(KEYINPUT95), .Z(n393) );
  XNOR2_X1 U459 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n390), .B(G127GAT), .ZN(n427) );
  XNOR2_X1 U461 ( .A(n427), .B(n391), .ZN(n392) );
  XNOR2_X1 U462 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n399) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n398) );
  XOR2_X1 U466 ( .A(n399), .B(n398), .Z(n522) );
  INV_X1 U467 ( .A(n522), .ZN(n490) );
  XOR2_X1 U468 ( .A(KEYINPUT19), .B(G183GAT), .Z(n401) );
  XNOR2_X1 U469 ( .A(KEYINPUT18), .B(KEYINPUT88), .ZN(n400) );
  XNOR2_X1 U470 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U471 ( .A(n402), .B(KEYINPUT17), .Z(n404) );
  XNOR2_X1 U472 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n404), .B(n403), .ZN(n430) );
  INV_X1 U474 ( .A(n405), .ZN(n409) );
  XOR2_X1 U475 ( .A(G92GAT), .B(G204GAT), .Z(n407) );
  XNOR2_X1 U476 ( .A(G36GAT), .B(G190GAT), .ZN(n406) );
  XNOR2_X1 U477 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U478 ( .A(n409), .B(n408), .Z(n415) );
  XOR2_X1 U479 ( .A(n411), .B(n410), .Z(n413) );
  NAND2_X1 U480 ( .A1(G226GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U483 ( .A(n430), .B(n416), .Z(n494) );
  XNOR2_X1 U484 ( .A(KEYINPUT27), .B(n494), .ZN(n441) );
  NAND2_X1 U485 ( .A1(n490), .A2(n441), .ZN(n531) );
  NOR2_X1 U486 ( .A1(n533), .A2(n531), .ZN(n433) );
  XOR2_X1 U487 ( .A(G99GAT), .B(n417), .Z(n420) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n426) );
  XOR2_X1 U490 ( .A(G176GAT), .B(KEYINPUT85), .Z(n422) );
  XNOR2_X1 U491 ( .A(KEYINPUT20), .B(KEYINPUT89), .ZN(n421) );
  XOR2_X1 U492 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U494 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U495 ( .A(G169GAT), .B(G15GAT), .Z(n429) );
  INV_X1 U496 ( .A(n496), .ZN(n534) );
  NAND2_X1 U497 ( .A1(n433), .A2(n534), .ZN(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n437) );
  AND2_X1 U499 ( .A1(n496), .A2(n494), .ZN(n434) );
  XOR2_X1 U500 ( .A(KEYINPUT98), .B(n434), .Z(n435) );
  NAND2_X1 U501 ( .A1(n435), .A2(n477), .ZN(n436) );
  XNOR2_X1 U502 ( .A(n437), .B(n436), .ZN(n439) );
  INV_X1 U503 ( .A(KEYINPUT25), .ZN(n438) );
  XNOR2_X1 U504 ( .A(n439), .B(n438), .ZN(n443) );
  NOR2_X1 U505 ( .A1(n477), .A2(n496), .ZN(n440) );
  XNOR2_X1 U506 ( .A(n440), .B(KEYINPUT26), .ZN(n571) );
  NAND2_X1 U507 ( .A1(n441), .A2(n571), .ZN(n442) );
  NAND2_X1 U508 ( .A1(n443), .A2(n442), .ZN(n444) );
  NAND2_X1 U509 ( .A1(n444), .A2(n522), .ZN(n445) );
  NAND2_X1 U510 ( .A1(n446), .A2(n445), .ZN(n447) );
  XNOR2_X1 U511 ( .A(n447), .B(KEYINPUT101), .ZN(n486) );
  NOR2_X1 U512 ( .A1(n588), .A2(n486), .ZN(n448) );
  NAND2_X1 U513 ( .A1(n555), .A2(n448), .ZN(n450) );
  NAND2_X1 U514 ( .A1(n488), .A2(n520), .ZN(n452) );
  XOR2_X1 U515 ( .A(KEYINPUT109), .B(KEYINPUT38), .Z(n451) );
  NOR2_X1 U516 ( .A1(n509), .A2(n522), .ZN(n455) );
  XNOR2_X1 U517 ( .A(KEYINPUT39), .B(KEYINPUT110), .ZN(n453) );
  INV_X1 U518 ( .A(n494), .ZN(n524) );
  XNOR2_X1 U519 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n456), .A2(KEYINPUT64), .ZN(n460) );
  INV_X1 U521 ( .A(KEYINPUT64), .ZN(n457) );
  NAND2_X1 U522 ( .A1(n458), .A2(n457), .ZN(n459) );
  NAND2_X1 U523 ( .A1(n460), .A2(n459), .ZN(n461) );
  INV_X1 U524 ( .A(n539), .ZN(n551) );
  NOR2_X1 U525 ( .A1(n573), .A2(n551), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n464) );
  INV_X1 U527 ( .A(n559), .ZN(n564) );
  NOR2_X1 U528 ( .A1(n464), .A2(n564), .ZN(n465) );
  NAND2_X1 U529 ( .A1(n555), .A2(n465), .ZN(n466) );
  XNOR2_X1 U530 ( .A(n466), .B(KEYINPUT47), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n588), .A2(n555), .ZN(n467) );
  XNOR2_X1 U532 ( .A(KEYINPUT45), .B(n467), .ZN(n469) );
  NAND2_X1 U533 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U534 ( .A1(n470), .A2(n578), .ZN(n471) );
  NOR2_X1 U535 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n473), .B(KEYINPUT48), .ZN(n532) );
  NOR2_X1 U537 ( .A1(n524), .A2(n532), .ZN(n474) );
  XNOR2_X1 U538 ( .A(KEYINPUT54), .B(n474), .ZN(n475) );
  NAND2_X1 U539 ( .A1(n572), .A2(n477), .ZN(n479) );
  XOR2_X1 U540 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X2 U542 ( .A1(n534), .A2(n480), .ZN(n565) );
  NAND2_X1 U543 ( .A1(n565), .A2(n539), .ZN(n483) );
  XOR2_X1 U544 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n481) );
  XOR2_X1 U545 ( .A(KEYINPUT104), .B(KEYINPUT34), .Z(n492) );
  NOR2_X1 U546 ( .A1(n564), .A2(n555), .ZN(n484) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U548 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT102), .B(n487), .ZN(n511) );
  NAND2_X1 U550 ( .A1(n511), .A2(n488), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(KEYINPUT103), .ZN(n501) );
  NAND2_X1 U552 ( .A1(n501), .A2(n490), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U554 ( .A(G1GAT), .B(n493), .Z(G1324GAT) );
  NAND2_X1 U555 ( .A1(n494), .A2(n501), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G8GAT), .B(n495), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n498) );
  NAND2_X1 U558 ( .A1(n501), .A2(n496), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n500) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT105), .Z(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  XOR2_X1 U562 ( .A(G22GAT), .B(KEYINPUT107), .Z(n503) );
  NAND2_X1 U563 ( .A1(n501), .A2(n533), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1327GAT) );
  NOR2_X1 U565 ( .A1(n509), .A2(n524), .ZN(n504) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT40), .B(KEYINPUT112), .Z(n506) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(KEYINPUT111), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n508) );
  NOR2_X1 U570 ( .A1(n534), .A2(n509), .ZN(n507) );
  XOR2_X1 U571 ( .A(n508), .B(n507), .Z(G1330GAT) );
  NOR2_X1 U572 ( .A1(n509), .A2(n528), .ZN(n510) );
  XOR2_X1 U573 ( .A(G50GAT), .B(n510), .Z(G1331GAT) );
  AND2_X1 U574 ( .A1(n539), .A2(n573), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n521), .A2(n511), .ZN(n517) );
  NOR2_X1 U576 ( .A1(n522), .A2(n517), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n524), .A2(n517), .ZN(n515) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n534), .A2(n517), .ZN(n516) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U584 ( .A1(n528), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U588 ( .A1(n522), .A2(n527), .ZN(n523) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n527), .ZN(n525) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n534), .A2(n527), .ZN(n526) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n529), .Z(n530) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n548) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n548), .A2(n535), .ZN(n536) );
  XNOR2_X1 U600 ( .A(KEYINPUT115), .B(n536), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n561), .A2(n544), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT116), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U605 ( .A1(n544), .A2(n539), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n583), .A2(n544), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U611 ( .A1(n544), .A2(n564), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NAND2_X1 U614 ( .A1(n548), .A2(n571), .ZN(n558) );
  NOR2_X1 U615 ( .A1(n573), .A2(n558), .ZN(n549) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n549), .Z(n550) );
  XNOR2_X1 U617 ( .A(KEYINPUT118), .B(n550), .ZN(G1344GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n558), .ZN(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n558), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NAND2_X1 U627 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n583), .A2(n565), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n568), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n587) );
  NOR2_X1 U639 ( .A1(n573), .A2(n587), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U644 ( .A(n587), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n582), .A2(n578), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U647 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n586) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n590) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U654 ( .A(n590), .B(n589), .Z(G1355GAT) );
endmodule

