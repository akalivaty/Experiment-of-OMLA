

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U323 ( .A(n356), .B(n355), .ZN(n399) );
  XNOR2_X1 U324 ( .A(n343), .B(KEYINPUT75), .ZN(n344) );
  XNOR2_X1 U325 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n405) );
  XNOR2_X1 U326 ( .A(n345), .B(n344), .ZN(n347) );
  XNOR2_X1 U327 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n451) );
  XNOR2_X1 U328 ( .A(n406), .B(n405), .ZN(n533) );
  XNOR2_X1 U329 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U330 ( .A(n374), .B(n373), .Z(n559) );
  XOR2_X1 U331 ( .A(n472), .B(KEYINPUT28), .Z(n537) );
  XNOR2_X1 U332 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1350GAT) );
  XOR2_X1 U334 ( .A(G176GAT), .B(G127GAT), .Z(n291) );
  XNOR2_X1 U335 ( .A(G169GAT), .B(G71GAT), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n291), .B(n290), .ZN(n307) );
  XOR2_X1 U337 ( .A(G120GAT), .B(G99GAT), .Z(n293) );
  XNOR2_X1 U338 ( .A(G15GAT), .B(G190GAT), .ZN(n292) );
  XNOR2_X1 U339 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U340 ( .A(n294), .B(G134GAT), .Z(n296) );
  XOR2_X1 U341 ( .A(G113GAT), .B(KEYINPUT0), .Z(n425) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(n425), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U344 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n298) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U348 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(KEYINPUT19), .B(n303), .Z(n316) );
  XNOR2_X1 U352 ( .A(n316), .B(KEYINPUT81), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n534) );
  XOR2_X1 U355 ( .A(G211GAT), .B(KEYINPUT21), .Z(n309) );
  XNOR2_X1 U356 ( .A(G197GAT), .B(G218GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n439) );
  INV_X1 U358 ( .A(G92GAT), .ZN(n310) );
  NAND2_X1 U359 ( .A1(G64GAT), .A2(n310), .ZN(n313) );
  INV_X1 U360 ( .A(G64GAT), .ZN(n311) );
  NAND2_X1 U361 ( .A1(n311), .A2(G92GAT), .ZN(n312) );
  NAND2_X1 U362 ( .A1(n313), .A2(n312), .ZN(n315) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n342) );
  XNOR2_X1 U365 ( .A(n439), .B(n342), .ZN(n323) );
  XOR2_X1 U366 ( .A(G36GAT), .B(G190GAT), .Z(n326) );
  XOR2_X1 U367 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n318) );
  XOR2_X1 U368 ( .A(G169GAT), .B(G8GAT), .Z(n362) );
  XNOR2_X1 U369 ( .A(n362), .B(n316), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n326), .B(n319), .Z(n321) );
  NAND2_X1 U372 ( .A1(G226GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n523) );
  XOR2_X1 U375 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n325) );
  XNOR2_X1 U376 ( .A(G92GAT), .B(KEYINPUT64), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n340) );
  XOR2_X1 U378 ( .A(G99GAT), .B(G85GAT), .Z(n341) );
  XOR2_X1 U379 ( .A(n326), .B(n341), .Z(n328) );
  XNOR2_X1 U380 ( .A(G162GAT), .B(G218GAT), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n333) );
  XOR2_X1 U382 ( .A(G29GAT), .B(G134GAT), .Z(n421) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n329), .B(KEYINPUT7), .ZN(n370) );
  XOR2_X1 U385 ( .A(n421), .B(n370), .Z(n331) );
  NAND2_X1 U386 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U389 ( .A(G50GAT), .B(KEYINPUT76), .Z(n438) );
  XOR2_X1 U390 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n335) );
  XNOR2_X1 U391 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U393 ( .A(n438), .B(n336), .Z(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n459) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n345) );
  AND2_X1 U397 ( .A1(G230GAT), .A2(G233GAT), .ZN(n343) );
  XOR2_X1 U398 ( .A(G106GAT), .B(G78GAT), .Z(n435) );
  XOR2_X1 U399 ( .A(n435), .B(KEYINPUT32), .Z(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n356) );
  XNOR2_X1 U401 ( .A(G120GAT), .B(G148GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n348), .B(G57GAT), .ZN(n420) );
  XOR2_X1 U403 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n350) );
  XNOR2_X1 U404 ( .A(G71GAT), .B(KEYINPUT72), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n381) );
  XNOR2_X1 U406 ( .A(n420), .B(n381), .ZN(n354) );
  XOR2_X1 U407 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n352) );
  XNOR2_X1 U408 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n351) );
  XOR2_X1 U409 ( .A(n352), .B(n351), .Z(n353) );
  XNOR2_X1 U410 ( .A(n399), .B(KEYINPUT41), .ZN(n551) );
  XOR2_X1 U411 ( .A(KEYINPUT70), .B(G1GAT), .Z(n358) );
  XNOR2_X1 U412 ( .A(G141GAT), .B(G113GAT), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n374) );
  XOR2_X1 U414 ( .A(G197GAT), .B(G50GAT), .Z(n360) );
  XNOR2_X1 U415 ( .A(G29GAT), .B(G36GAT), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n364) );
  AND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U420 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n366) );
  XNOR2_X1 U421 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U423 ( .A(n368), .B(n367), .Z(n372) );
  XNOR2_X1 U424 ( .A(G22GAT), .B(G15GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n369), .B(KEYINPUT69), .ZN(n377) );
  XNOR2_X1 U426 ( .A(n370), .B(n377), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  AND2_X1 U428 ( .A1(n551), .A2(n559), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n375), .B(KEYINPUT46), .ZN(n376) );
  NOR2_X1 U430 ( .A1(n459), .A2(n376), .ZN(n396) );
  XOR2_X1 U431 ( .A(G1GAT), .B(G127GAT), .Z(n418) );
  XOR2_X1 U432 ( .A(n418), .B(n377), .Z(n379) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U435 ( .A(n380), .B(KEYINPUT14), .Z(n383) );
  XNOR2_X1 U436 ( .A(n381), .B(KEYINPUT15), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U438 ( .A(G78GAT), .B(G211GAT), .Z(n385) );
  XNOR2_X1 U439 ( .A(G183GAT), .B(G155GAT), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n395) );
  XOR2_X1 U442 ( .A(KEYINPUT77), .B(KEYINPUT80), .Z(n389) );
  XNOR2_X1 U443 ( .A(KEYINPUT79), .B(KEYINPUT12), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U445 ( .A(KEYINPUT78), .B(G64GAT), .Z(n391) );
  XNOR2_X1 U446 ( .A(G8GAT), .B(G57GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U448 ( .A(n393), .B(n392), .Z(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n577) );
  NAND2_X1 U450 ( .A1(n396), .A2(n577), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n397), .B(KEYINPUT47), .ZN(n404) );
  XOR2_X1 U452 ( .A(KEYINPUT36), .B(n459), .Z(n581) );
  NOR2_X1 U453 ( .A1(n577), .A2(n581), .ZN(n398) );
  XNOR2_X1 U454 ( .A(KEYINPUT45), .B(n398), .ZN(n400) );
  NAND2_X1 U455 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U456 ( .A(KEYINPUT114), .B(n401), .ZN(n402) );
  NOR2_X1 U457 ( .A1(n402), .A2(n559), .ZN(n403) );
  NOR2_X1 U458 ( .A1(n404), .A2(n403), .ZN(n406) );
  NAND2_X1 U459 ( .A1(n523), .A2(n533), .ZN(n407) );
  XNOR2_X1 U460 ( .A(n407), .B(KEYINPUT54), .ZN(n409) );
  INV_X1 U461 ( .A(KEYINPUT120), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n565) );
  XNOR2_X1 U463 ( .A(G155GAT), .B(KEYINPUT86), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n410), .B(KEYINPUT3), .ZN(n411) );
  XOR2_X1 U465 ( .A(n411), .B(KEYINPUT2), .Z(n413) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(G162GAT), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n447) );
  INV_X1 U468 ( .A(n447), .ZN(n431) );
  XOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n415) );
  XNOR2_X1 U470 ( .A(KEYINPUT1), .B(KEYINPUT89), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n429) );
  XOR2_X1 U472 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n417) );
  XNOR2_X1 U473 ( .A(G85GAT), .B(KEYINPUT5), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U475 ( .A(n419), .B(n418), .Z(n427) );
  XOR2_X1 U476 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U481 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n469) );
  XNOR2_X1 U483 ( .A(KEYINPUT92), .B(n469), .ZN(n521) );
  INV_X1 U484 ( .A(n521), .ZN(n564) );
  XOR2_X1 U485 ( .A(G204GAT), .B(KEYINPUT22), .Z(n433) );
  XNOR2_X1 U486 ( .A(KEYINPUT24), .B(KEYINPUT87), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U488 ( .A(n434), .B(G148GAT), .Z(n437) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U491 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n449) );
  XOR2_X1 U495 ( .A(KEYINPUT23), .B(KEYINPUT84), .Z(n445) );
  XNOR2_X1 U496 ( .A(KEYINPUT88), .B(KEYINPUT85), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n472) );
  AND2_X1 U500 ( .A1(n564), .A2(n472), .ZN(n450) );
  NAND2_X1 U501 ( .A1(n565), .A2(n450), .ZN(n452) );
  NOR2_X1 U502 ( .A1(n534), .A2(n453), .ZN(n561) );
  NAND2_X1 U503 ( .A1(n561), .A2(n551), .ZN(n456) );
  XOR2_X1 U504 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n454) );
  XNOR2_X1 U505 ( .A(n454), .B(G176GAT), .ZN(n455) );
  XNOR2_X1 U506 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  INV_X1 U507 ( .A(n577), .ZN(n555) );
  NAND2_X1 U508 ( .A1(n555), .A2(n561), .ZN(n458) );
  XOR2_X1 U509 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n481) );
  NAND2_X1 U510 ( .A1(n559), .A2(n399), .ZN(n494) );
  NOR2_X1 U511 ( .A1(n577), .A2(n459), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT16), .ZN(n478) );
  INV_X1 U513 ( .A(n534), .ZN(n527) );
  NAND2_X1 U514 ( .A1(n523), .A2(n527), .ZN(n461) );
  NAND2_X1 U515 ( .A1(n461), .A2(n472), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n462), .B(KEYINPUT97), .ZN(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(n463), .Z(n467) );
  XOR2_X1 U518 ( .A(n523), .B(KEYINPUT27), .Z(n471) );
  NOR2_X1 U519 ( .A1(n527), .A2(n472), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT26), .B(n464), .Z(n566) );
  NOR2_X1 U521 ( .A1(n471), .A2(n566), .ZN(n465) );
  XNOR2_X1 U522 ( .A(KEYINPUT96), .B(n465), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  XOR2_X1 U525 ( .A(KEYINPUT98), .B(n470), .Z(n477) );
  NOR2_X1 U526 ( .A1(n564), .A2(n471), .ZN(n532) );
  INV_X1 U527 ( .A(n537), .ZN(n473) );
  NAND2_X1 U528 ( .A1(n532), .A2(n473), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n474), .B(KEYINPUT95), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n475), .A2(n534), .ZN(n476) );
  NAND2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n491) );
  NAND2_X1 U532 ( .A1(n478), .A2(n491), .ZN(n507) );
  NOR2_X1 U533 ( .A1(n494), .A2(n507), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT99), .B(n479), .Z(n488) );
  NAND2_X1 U535 ( .A1(n488), .A2(n521), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n482), .Z(G1324GAT) );
  XOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT101), .Z(n484) );
  NAND2_X1 U539 ( .A1(n488), .A2(n523), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U542 ( .A1(n488), .A2(n527), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  XOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT103), .Z(n490) );
  NAND2_X1 U546 ( .A1(n488), .A2(n537), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n490), .B(n489), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n497) );
  NAND2_X1 U549 ( .A1(n577), .A2(n491), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n492), .A2(n581), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n493), .B(KEYINPUT37), .ZN(n520) );
  NOR2_X1 U552 ( .A1(n494), .A2(n520), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT38), .ZN(n505) );
  NAND2_X1 U554 ( .A1(n505), .A2(n521), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(n498), .ZN(G1328GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n500) );
  NAND2_X1 U558 ( .A1(n523), .A2(n505), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n503) );
  NAND2_X1 U562 ( .A1(n527), .A2(n505), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n505), .A2(n537), .ZN(n506) );
  XNOR2_X1 U566 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n509) );
  INV_X1 U568 ( .A(n559), .ZN(n569) );
  NAND2_X1 U569 ( .A1(n569), .A2(n551), .ZN(n519) );
  NOR2_X1 U570 ( .A1(n507), .A2(n519), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n515), .A2(n521), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n510), .Z(G1332GAT) );
  XOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT109), .Z(n512) );
  NAND2_X1 U575 ( .A1(n515), .A2(n523), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n515), .A2(n527), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT110), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n537), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n518), .Z(G1335GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n529) );
  NAND2_X1 U585 ( .A1(n529), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n525) );
  NAND2_X1 U588 ( .A1(n529), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n529), .A2(n527), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n537), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  XOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT117), .Z(n539) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n549) );
  NOR2_X1 U598 ( .A1(n534), .A2(n549), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(n535), .Z(n536) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n546), .A2(n559), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U604 ( .A1(n546), .A2(n551), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n543) );
  NAND2_X1 U608 ( .A1(n546), .A2(n555), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U612 ( .A1(n546), .A2(n459), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n566), .A2(n549), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n559), .A2(n557), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U618 ( .A1(n557), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n557), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n459), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n561), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n459), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G190GAT), .ZN(G1351GAT) );
  AND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n568) );
  INV_X1 U631 ( .A(n566), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n580) );
  NOR2_X1 U633 ( .A1(n569), .A2(n580), .ZN(n574) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT59), .B(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n399), .A2(n580), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n580), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(G218GAT), .B(n584), .Z(G1355GAT) );
endmodule

