//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n562, new_n563, new_n564, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g024(.A(G2106), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT65), .Z(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n450), .B1(new_n458), .B2(new_n455), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT67), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n463), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n462), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n472), .A2(G137), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND3_X1  g052(.A1(new_n472), .A2(G2105), .A3(new_n474), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n473), .A2(G112), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n480), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT68), .Z(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n490), .A2(new_n463), .A3(new_n465), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n472), .A2(G138), .A3(new_n473), .A4(new_n474), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n472), .A2(G126), .A3(G2105), .A4(new_n474), .ZN(new_n496));
  OR3_X1    g071(.A1(new_n473), .A2(KEYINPUT69), .A3(G114), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT69), .B1(new_n473), .B2(G114), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n497), .A2(G2104), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n495), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(G88), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(KEYINPUT71), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n505), .A2(new_n507), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n514), .A2(new_n515), .B1(G651), .B2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n508), .A2(new_n509), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n509), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n523), .A2(new_n525), .A3(new_n527), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n509), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n521), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(new_n522), .A2(G81), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n526), .A2(G43), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n532), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  AOI22_X1  g125(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(KEYINPUT72), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(KEYINPUT72), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n552), .A2(G651), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n526), .A2(new_n555), .A3(G53), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n535), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n556), .A2(new_n558), .B1(G91), .B2(new_n522), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n554), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  NAND2_X1  g136(.A1(new_n519), .A2(G651), .ZN(new_n562));
  INV_X1    g137(.A(new_n515), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT71), .B1(new_n510), .B2(new_n511), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(G303));
  OR2_X1    g140(.A1(new_n508), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(G49), .B2(new_n526), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n568));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n521), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n522), .A2(KEYINPUT73), .A3(G87), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(G288));
  AOI22_X1  g147(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n532), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  INV_X1    g150(.A(G48), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n521), .A2(new_n575), .B1(new_n535), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n532), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n521), .A2(new_n582), .B1(new_n535), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n517), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT10), .B1(new_n521), .B2(new_n592), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n521), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n587), .B1(new_n596), .B2(G868), .ZN(G321));
  XNOR2_X1  g172(.A(G321), .B(KEYINPUT74), .ZN(G284));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G299), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n599), .B2(G168), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(new_n599), .B2(G168), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  NOR2_X1   g179(.A1(new_n595), .A2(G559), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n605), .A2(KEYINPUT75), .A3(new_n599), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT75), .B1(new_n605), .B2(new_n599), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n544), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n479), .A2(G123), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n482), .A2(G135), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n473), .A2(G111), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  NAND3_X1  g190(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2100), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(G2451), .B(G2454), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT76), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(G2443), .B(G2446), .Z(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n631), .A2(new_n633), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n622), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n631), .A2(new_n633), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n638), .A2(new_n621), .A3(new_n634), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n637), .A2(new_n639), .A3(G14), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(G401));
  XNOR2_X1  g216(.A(G2072), .B(G2078), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT17), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n642), .B(KEYINPUT78), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n647), .C1(new_n644), .C2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT79), .ZN(new_n650));
  OR3_X1    g225(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n644), .A3(new_n642), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT77), .B(KEYINPUT18), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n650), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT80), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XOR2_X1   g234(.A(KEYINPUT81), .B(KEYINPUT19), .Z(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT82), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(KEYINPUT82), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n664), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n668), .B(new_n670), .C1(new_n661), .C2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  INV_X1    g251(.A(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G25), .ZN(new_n682));
  AOI22_X1  g257(.A1(G119), .A2(new_n479), .B1(new_n482), .B2(G131), .ZN(new_n683));
  OR2_X1    g258(.A1(G95), .A2(G2105), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n684), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT83), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n682), .B1(new_n688), .B2(new_n681), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT35), .B(G1991), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G24), .ZN(new_n692));
  OAI21_X1  g267(.A(KEYINPUT84), .B1(new_n692), .B2(G16), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n692), .A2(KEYINPUT84), .A3(G16), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n693), .B(new_n694), .C1(new_n585), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1986), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G23), .ZN(new_n699));
  AND3_X1   g274(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT33), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n695), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G6), .A2(G16), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n578), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n703), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(KEYINPUT34), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n714), .A2(new_n713), .A3(KEYINPUT34), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n713), .B2(KEYINPUT34), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n698), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT86), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n714), .B(new_n719), .Z(new_n720));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n720), .A2(new_n721), .A3(new_n698), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n718), .A2(new_n722), .A3(KEYINPUT36), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n717), .A2(KEYINPUT86), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n479), .A2(G128), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n482), .A2(G140), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n473), .A2(G116), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n681), .A2(G26), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2067), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n695), .A2(G4), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n596), .B2(new_n695), .ZN(new_n741));
  INV_X1    g316(.A(G1348), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n544), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G16), .B2(G19), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT87), .B(G1341), .Z(new_n748));
  XOR2_X1   g323(.A(new_n747), .B(new_n748), .Z(new_n749));
  OAI21_X1  g324(.A(new_n727), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n743), .A2(new_n744), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n747), .B(new_n748), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n751), .A2(KEYINPUT89), .A3(new_n739), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n479), .A2(G129), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT92), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n482), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n469), .A2(G105), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n756), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n755), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  OR2_X1    g338(.A1(G29), .A2(G32), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT27), .B(G1996), .Z(new_n765));
  NAND3_X1  g340(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  NOR2_X1   g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n767), .A2(new_n768), .A3(G29), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n476), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G171), .A2(G16), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G5), .B2(G16), .ZN(new_n774));
  INV_X1    g349(.A(G1961), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n766), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n766), .A2(KEYINPUT97), .A3(new_n772), .A4(new_n776), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n750), .A2(new_n753), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n463), .A2(new_n465), .A3(G127), .ZN(new_n782));
  INV_X1    g357(.A(G115), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n462), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT90), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G2105), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n482), .A2(G139), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n469), .A2(G103), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G2072), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n695), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n695), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT94), .B(G1966), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT31), .B(G11), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n614), .A2(new_n681), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT30), .B(G28), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n799), .B(new_n800), .C1(new_n681), .C2(new_n801), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n797), .B(new_n802), .C1(new_n775), .C2(new_n774), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n763), .A2(new_n764), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(new_n765), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n781), .A2(new_n792), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G27), .A2(G29), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G164), .B2(G29), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT98), .B(G2078), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n681), .A2(G35), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n681), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(G2090), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n808), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n695), .A2(G20), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT99), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT23), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G299), .B2(G16), .ZN(new_n821));
  INV_X1    g396(.A(G1956), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n815), .B2(G2090), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT100), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n770), .A2(new_n771), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT91), .Z(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n817), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n808), .A2(new_n827), .A3(new_n812), .A4(new_n816), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n831), .A2(new_n832), .A3(new_n825), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n726), .B1(new_n830), .B2(new_n833), .ZN(G311));
  INV_X1    g409(.A(new_n726), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n831), .A2(new_n832), .A3(new_n825), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n832), .B1(new_n831), .B2(new_n825), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(G150));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  INV_X1    g414(.A(G80), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n517), .A2(new_n839), .B1(new_n840), .B2(new_n504), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  OAI221_X1 g418(.A(new_n843), .B1(new_n840), .B2(new_n504), .C1(new_n517), .C2(new_n839), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(G651), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n522), .A2(G93), .B1(new_n526), .B2(G55), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  OAI211_X1 g424(.A(new_n539), .B(new_n540), .C1(new_n532), .C2(new_n542), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n850), .A3(new_n846), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n845), .B2(new_n846), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT39), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n595), .A2(new_n603), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n855), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n849), .B1(new_n859), .B2(G860), .ZN(G145));
  NAND2_X1  g435(.A1(new_n479), .A2(G130), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n482), .A2(G142), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n473), .A2(G118), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n732), .B(new_n865), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n688), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n790), .A2(new_n617), .ZN(new_n868));
  INV_X1    g443(.A(new_n617), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n786), .A2(new_n869), .A3(new_n787), .A4(new_n789), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n762), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n762), .B1(new_n868), .B2(new_n870), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n492), .ZN(new_n876));
  INV_X1    g451(.A(new_n501), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n495), .A2(new_n501), .A3(KEYINPUT104), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n872), .A2(new_n873), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n868), .A2(new_n870), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n755), .A2(new_n761), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n885), .B2(new_n871), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n867), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n880), .B1(new_n872), .B2(new_n873), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n866), .B(new_n687), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n882), .A3(new_n871), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n614), .B(G160), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n487), .B(new_n893), .Z(new_n894));
  AOI21_X1  g469(.A(G37), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n887), .A2(new_n896), .A3(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT105), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n887), .A2(new_n899), .A3(new_n896), .A4(new_n891), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n895), .A2(new_n898), .A3(KEYINPUT106), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g481(.A1(new_n847), .A2(G868), .ZN(new_n907));
  XNOR2_X1  g482(.A(G290), .B(G288), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT109), .ZN(new_n909));
  XNOR2_X1  g484(.A(G303), .B(new_n578), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n908), .B(KEYINPUT109), .Z(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(new_n910), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n554), .A2(KEYINPUT107), .A3(new_n559), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n596), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT107), .B1(new_n554), .B2(new_n559), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NAND2_X1  g495(.A1(G299), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(new_n596), .A3(new_n916), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT41), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n919), .A2(new_n922), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n854), .B(new_n605), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n923), .B2(new_n929), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n914), .B(new_n915), .C1(new_n932), .C2(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(KEYINPUT110), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n933), .B(new_n934), .Z(new_n935));
  AOI21_X1  g510(.A(new_n907), .B1(new_n935), .B2(G868), .ZN(G295));
  AOI21_X1  g511(.A(new_n907), .B1(new_n935), .B2(G868), .ZN(G331));
  OAI211_X1 g512(.A(KEYINPUT111), .B(G171), .C1(new_n852), .C2(new_n853), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n939));
  AOI21_X1  g514(.A(G168), .B1(new_n939), .B2(G301), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n847), .A2(new_n544), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n941), .B(new_n851), .C1(new_n939), .C2(G301), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n938), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n940), .B1(new_n938), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n928), .A3(new_n930), .ZN(new_n946));
  INV_X1    g521(.A(new_n923), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n943), .B2(new_n944), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n913), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G37), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n913), .B1(new_n946), .B2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n924), .A2(new_n955), .A3(new_n927), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n947), .A2(KEYINPUT113), .A3(new_n926), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n945), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT114), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n945), .A2(new_n956), .A3(new_n960), .A4(new_n957), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n948), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n913), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  INV_X1    g540(.A(new_n951), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(KEYINPUT43), .C1(new_n951), .C2(new_n952), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n954), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n966), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n951), .A2(new_n952), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT44), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(G397));
  XOR2_X1   g552(.A(G171), .B(KEYINPUT54), .Z(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n495), .B2(new_n501), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT50), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n468), .A2(G2105), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n469), .A2(G101), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(G40), .A3(new_n475), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT115), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n470), .A2(new_n986), .A3(G40), .A4(new_n475), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n989), .B(new_n979), .C1(new_n495), .C2(new_n501), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n981), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n775), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT45), .B(new_n979), .C1(new_n878), .C2(new_n879), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n876), .A2(new_n874), .A3(new_n877), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT104), .B1(new_n495), .B2(new_n501), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(KEYINPUT117), .A3(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G2078), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1003), .A2(new_n980), .B1(new_n985), .B2(new_n987), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n993), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n984), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1006), .A2(G2078), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1003), .B1(new_n880), .B2(G1384), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1001), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n978), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n876), .B2(new_n877), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n988), .B1(KEYINPUT45), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n996), .B2(new_n1000), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT53), .B1(new_n1015), .B2(new_n1002), .ZN(new_n1016));
  INV_X1    g591(.A(new_n978), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT45), .B(new_n979), .C1(new_n495), .C2(new_n501), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1004), .A2(new_n1018), .A3(new_n1009), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR4_X1   g595(.A1(new_n1016), .A2(new_n1017), .A3(new_n993), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(G166), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(G303), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n991), .A2(G2090), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n994), .A2(new_n995), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT117), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1004), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1032), .B1(new_n1035), .B2(new_n706), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1031), .B1(new_n1036), .B2(new_n1027), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1032), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n1015), .B2(G1971), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1030), .A2(KEYINPUT119), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1025), .A2(new_n1028), .A3(new_n1041), .A4(new_n1029), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1043), .A3(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n578), .A2(new_n677), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT120), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n578), .A2(new_n677), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OR3_X1    g623(.A1(new_n578), .A2(KEYINPUT120), .A3(new_n677), .ZN(new_n1049));
  NAND2_X1  g624(.A1(KEYINPUT121), .A2(KEYINPUT49), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n1048), .A2(new_n1051), .B1(KEYINPUT121), .B2(KEYINPUT49), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1027), .B1(new_n988), .B2(new_n1013), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1047), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(KEYINPUT120), .A3(new_n1045), .ZN(new_n1055));
  NOR2_X1   g630(.A1(KEYINPUT121), .A2(KEYINPUT49), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n1050), .A4(new_n1049), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1053), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n700), .A2(G1976), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1053), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1060), .B(new_n1061), .C1(G1976), .C2(new_n700), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1058), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1037), .A2(new_n1044), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1018), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n796), .B1(new_n1014), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n981), .A2(new_n988), .A3(new_n771), .A4(new_n990), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(G168), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1066), .B1(new_n1070), .B2(G8), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n795), .B1(new_n1004), .B2(new_n1018), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1069), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1072), .A2(new_n1073), .A3(G286), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n1027), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT51), .B1(new_n1076), .B2(G168), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1071), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1022), .A2(new_n1065), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1004), .B(new_n1081), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT122), .B1(new_n556), .B2(new_n558), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(KEYINPUT57), .ZN(new_n1084));
  XOR2_X1   g659(.A(G299), .B(new_n1084), .Z(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n991), .A2(new_n822), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1082), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1080), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1085), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1082), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n991), .A2(new_n742), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n988), .A2(new_n738), .A3(new_n1013), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1096), .A2(KEYINPUT123), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT123), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1098), .A2(new_n1099), .A3(KEYINPUT60), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT60), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n596), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT60), .B(new_n595), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  INV_X1    g680(.A(G1996), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n1004), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT58), .B(G1341), .Z(new_n1108));
  INV_X1    g683(.A(new_n988), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(new_n980), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1105), .B1(new_n1111), .B2(new_n544), .ZN(new_n1112));
  AOI211_X1 g687(.A(KEYINPUT59), .B(new_n850), .C1(new_n1107), .C2(new_n1110), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1095), .A2(new_n1104), .A3(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1098), .A2(new_n1099), .A3(new_n595), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1089), .B1(KEYINPUT124), .B2(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1116), .A2(KEYINPUT124), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1088), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1079), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n1121));
  AOI21_X1  g696(.A(G301), .B1(new_n1078), .B2(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1039), .A2(G8), .A3(new_n1043), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1030), .B1(new_n1039), .B2(G8), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1058), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1007), .A2(new_n1019), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1122), .A2(new_n1126), .A3(KEYINPUT125), .A4(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1078), .A2(new_n1121), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1127), .A2(new_n1037), .A3(new_n1044), .A4(new_n1064), .ZN(new_n1131));
  AOI21_X1  g706(.A(G168), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1132));
  OAI211_X1 g707(.A(G8), .B(new_n1070), .C1(new_n1132), .C2(new_n1066), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT51), .B1(new_n1074), .B2(new_n1027), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n1121), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G171), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1130), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1128), .A2(new_n1129), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1076), .A2(new_n1027), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1126), .A2(KEYINPUT63), .A3(G168), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1037), .A2(new_n1064), .A3(G168), .A4(new_n1044), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1139), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G1976), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1058), .A2(new_n1146), .A3(new_n700), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1045), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1053), .A2(new_n1148), .B1(new_n1123), .B2(new_n1064), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1120), .A2(new_n1138), .A3(new_n1145), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1010), .A2(new_n1109), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n687), .B(new_n690), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT116), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n732), .B(new_n738), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n762), .A2(G1996), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n884), .A2(new_n1106), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n585), .B(G1986), .Z(new_n1160));
  OAI21_X1  g735(.A(new_n1151), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1150), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1151), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1163), .B1(new_n762), .B2(new_n1154), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1151), .A2(KEYINPUT46), .A3(new_n1106), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT46), .B1(new_n1151), .B2(new_n1106), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT47), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1163), .A2(G1986), .A3(G290), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT48), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1151), .B2(new_n1159), .ZN(new_n1171));
  OR3_X1    g746(.A1(new_n1157), .A2(new_n690), .A3(new_n687), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n732), .A2(G2067), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1163), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1168), .A2(new_n1171), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1162), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n1178));
  NOR2_X1   g752(.A1(G227), .A2(new_n460), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n640), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g756(.A(G229), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n640), .A2(KEYINPUT126), .A3(new_n1179), .ZN(new_n1184));
  AND4_X1   g758(.A1(new_n1178), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1185), .B1(new_n903), .B2(new_n904), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1187), .A2(KEYINPUT127), .ZN(new_n1188));
  AND3_X1   g762(.A1(new_n1186), .A2(new_n970), .A3(new_n1188), .ZN(G308));
  NAND3_X1  g763(.A1(new_n1186), .A2(new_n970), .A3(new_n1188), .ZN(G225));
endmodule


