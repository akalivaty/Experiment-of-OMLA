//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT67), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT68), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT69), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT70), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  INV_X1    g040(.A(G113), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(new_n461), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n469), .A2(new_n471), .A3(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n463), .B1(new_n461), .B2(KEYINPUT72), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n461), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n474), .A2(new_n478), .B1(G101), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT73), .ZN(G160));
  XNOR2_X1  g057(.A(KEYINPUT71), .B(G2105), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n483), .C2(G112), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n478), .A2(new_n472), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n478), .A2(new_n468), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(G136), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT74), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n462), .A2(new_n464), .A3(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(new_n472), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n478), .A2(new_n483), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n479), .A2(G102), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT3), .B1(new_n476), .B2(G2104), .ZN(new_n501));
  OAI21_X1  g076(.A(G126), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n468), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT75), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT76), .B(G51), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n520), .A2(new_n522), .A3(G543), .A4(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT77), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n508), .A2(new_n521), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n525), .B1(new_n524), .B2(new_n526), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n537), .A2(KEYINPUT78), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(KEYINPUT78), .ZN(new_n539));
  NOR3_X1   g114(.A1(new_n538), .A2(new_n539), .A3(new_n510), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n520), .A2(new_n522), .A3(G543), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n530), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n540), .A2(new_n544), .ZN(G171));
  AND3_X1   g120(.A1(new_n520), .A2(new_n522), .A3(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G43), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n510), .ZN(new_n549));
  INV_X1    g124(.A(new_n530), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND3_X1  g133(.A1(new_n546), .A2(KEYINPUT9), .A3(G53), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n541), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n508), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n510), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(G91), .B2(new_n550), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(new_n535), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n570), .A2(new_n527), .A3(new_n533), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  AND2_X1   g147(.A1(new_n546), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n530), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n573), .A2(new_n576), .ZN(G288));
  AOI22_X1  g152(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n510), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n530), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  AND2_X1   g159(.A1(new_n508), .A2(G60), .ZN(new_n585));
  AND2_X1   g160(.A1(G72), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(KEYINPUT79), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G85), .B2(new_n550), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(KEYINPUT79), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n546), .A2(G47), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  INV_X1    g168(.A(G54), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n541), .A2(new_n594), .B1(new_n510), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT80), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n550), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(G168), .A2(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n608), .ZN(G297));
  OAI211_X1 g184(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n608), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n601), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT82), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g192(.A1(new_n462), .A2(new_n464), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n479), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  INV_X1    g197(.A(new_n486), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n483), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n489), .A2(KEYINPUT83), .A3(G135), .ZN(new_n627));
  AOI21_X1  g202(.A(KEYINPUT83), .B1(new_n489), .B2(G135), .ZN(new_n628));
  OAI221_X1 g203(.A(new_n624), .B1(new_n625), .B2(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n622), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT86), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT15), .B(G2435), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n644), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G14), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n640), .A2(new_n648), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT17), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  OR3_X1    g233(.A1(new_n655), .A2(new_n653), .A3(new_n656), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n655), .A2(new_n653), .A3(new_n656), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n630), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G1986), .Z(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  INV_X1    g255(.A(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n682), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(G229));
  MUX2_X1   g260(.A(G23), .B(G288), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT91), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT33), .B(G1976), .Z(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(KEYINPUT92), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n687), .B(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n693));
  NOR2_X1   g268(.A1(G6), .A2(G16), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n583), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT32), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1981), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT89), .B(G16), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1971), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n691), .A2(new_n693), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  MUX2_X1   g282(.A(G24), .B(G290), .S(new_n699), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1986), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT87), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n489), .A2(G131), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n623), .A2(G119), .ZN(new_n714));
  OAI221_X1 g289(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n483), .C2(G107), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n712), .B1(new_n716), .B2(G29), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT88), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n709), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n706), .A2(new_n707), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n710), .B1(KEYINPUT24), .B2(G34), .ZN(new_n726));
  OAI22_X1  g301(.A1(G160), .A2(new_n710), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2084), .ZN(new_n728));
  NOR2_X1   g303(.A1(G27), .A2(G29), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G164), .B2(G29), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G2078), .ZN(new_n731));
  INV_X1    g306(.A(G28), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(KEYINPUT30), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n732), .B2(KEYINPUT30), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT31), .A2(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n629), .B2(new_n710), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G2078), .B2(new_n730), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n710), .A2(G33), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT93), .Z(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT25), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n618), .A2(G127), .ZN(new_n746));
  INV_X1    g321(.A(G115), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n461), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n748), .A2(new_n472), .B1(G139), .B2(new_n489), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n744), .A2(new_n745), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n741), .B1(new_n750), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(G2072), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n710), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  OAI221_X1 g330(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n483), .C2(G116), .ZN(new_n756));
  INV_X1    g331(.A(G140), .ZN(new_n757));
  INV_X1    g332(.A(G128), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n756), .B1(new_n488), .B2(new_n757), .C1(new_n758), .C2(new_n486), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n755), .B1(new_n759), .B2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G2067), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n728), .A2(new_n740), .A3(new_n753), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n699), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n553), .B2(new_n699), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1341), .ZN(new_n766));
  INV_X1    g341(.A(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G5), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G171), .B2(new_n767), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1961), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n766), .B(new_n770), .C1(G2072), .C2(new_n752), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT26), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n774), .A2(new_n775), .B1(G105), .B2(new_n479), .ZN(new_n776));
  INV_X1    g351(.A(G141), .ZN(new_n777));
  INV_X1    g352(.A(G129), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n776), .B1(new_n488), .B2(new_n777), .C1(new_n778), .C2(new_n486), .ZN(new_n779));
  MUX2_X1   g354(.A(G32), .B(new_n779), .S(G29), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT27), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1996), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n767), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n767), .ZN(new_n784));
  INV_X1    g359(.A(G1966), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n763), .A2(new_n771), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G29), .A2(G35), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G162), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2090), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n698), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT95), .B(KEYINPUT23), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n608), .B2(new_n767), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1956), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n767), .A2(G4), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n601), .B2(new_n767), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n797), .B1(G1348), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n792), .B(new_n800), .C1(G1348), .C2(new_n799), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n724), .A2(new_n787), .A3(new_n801), .ZN(G311));
  OR3_X1    g377(.A1(new_n724), .A2(new_n787), .A3(new_n801), .ZN(G150));
  NAND2_X1  g378(.A1(new_n550), .A2(G93), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n805));
  INV_X1    g380(.A(G55), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n804), .B1(new_n510), .B2(new_n805), .C1(new_n806), .C2(new_n541), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G860), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT37), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n601), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n552), .B(new_n807), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT97), .ZN(new_n817));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n815), .B2(KEYINPUT39), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n809), .B1(new_n817), .B2(new_n819), .ZN(G145));
  AOI22_X1  g395(.A1(G130), .A2(new_n623), .B1(new_n489), .B2(G142), .ZN(new_n821));
  INV_X1    g396(.A(G118), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n472), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n620), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n716), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT99), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n506), .B(new_n759), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n779), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n750), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n830), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(G160), .B(new_n629), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G162), .ZN(new_n836));
  AOI21_X1  g411(.A(G37), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n836), .B(KEYINPUT100), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n833), .A2(new_n829), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n838), .B(new_n839), .C1(new_n830), .C2(new_n833), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g417(.A1(new_n807), .A2(new_n604), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n613), .B(new_n811), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n600), .A2(new_n608), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT41), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n600), .B2(new_n608), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n597), .A2(KEYINPUT101), .A3(G299), .A4(new_n599), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n852), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT41), .B1(new_n856), .B2(new_n846), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n846), .B1(new_n853), .B2(new_n854), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n844), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n845), .A2(new_n859), .B1(new_n861), .B2(KEYINPUT103), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(KEYINPUT103), .B2(new_n861), .ZN(new_n863));
  XNOR2_X1  g438(.A(G290), .B(new_n583), .ZN(new_n864));
  XNOR2_X1  g439(.A(G288), .B(G166), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n863), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n843), .B1(new_n868), .B2(new_n604), .ZN(G295));
  OAI21_X1  g444(.A(new_n843), .B1(new_n868), .B2(new_n604), .ZN(G331));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n872));
  AOI21_X1  g447(.A(G286), .B1(G171), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(G171), .ZN(new_n874));
  NAND3_X1  g449(.A1(G301), .A2(KEYINPUT104), .A3(G286), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n811), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(KEYINPUT105), .A3(new_n811), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n876), .A2(new_n811), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n885), .B2(new_n846), .ZN(new_n886));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n877), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n881), .A2(new_n886), .B1(new_n859), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g464(.A(KEYINPUT106), .B(new_n871), .C1(new_n889), .C2(new_n866), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n847), .B1(new_n883), .B2(new_n884), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n892), .B2(new_n857), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n860), .A2(new_n887), .A3(new_n880), .A4(new_n879), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n866), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n895), .B2(G37), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n866), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n890), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n881), .A2(new_n887), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n848), .A2(new_n856), .ZN(new_n901));
  INV_X1    g476(.A(new_n846), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n883), .B2(new_n884), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n903), .B2(KEYINPUT41), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n900), .A2(new_n904), .B1(new_n877), .B2(new_n886), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(new_n866), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n897), .A2(new_n871), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n906), .A2(KEYINPUT107), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n871), .B(new_n897), .C1(new_n905), .C2(new_n866), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(KEYINPUT43), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n899), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n898), .A2(new_n907), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n911), .A2(new_n907), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(G397));
  INV_X1    g494(.A(G1384), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n504), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n473), .A2(new_n480), .A3(G40), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n927), .A2(G290), .A3(G1986), .ZN(new_n928));
  AND3_X1   g503(.A1(G290), .A2(G1986), .A3(new_n926), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n930), .B(KEYINPUT108), .Z(new_n931));
  XNOR2_X1  g506(.A(new_n759), .B(new_n761), .ZN(new_n932));
  INV_X1    g507(.A(G1996), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n779), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n716), .B(new_n719), .Z(new_n936));
  OAI21_X1  g511(.A(new_n926), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n922), .ZN(new_n939));
  INV_X1    g514(.A(new_n925), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1976), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n941), .B(G8), .C1(G288), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT52), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT111), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n583), .B(new_n681), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT49), .ZN(new_n948));
  INV_X1    g523(.A(new_n941), .ZN(new_n949));
  INV_X1    g524(.A(G8), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n943), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT52), .B1(G288), .B2(new_n942), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n499), .B2(new_n505), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n960), .A2(new_n961), .B1(new_n922), .B2(KEYINPUT50), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n921), .B2(new_n504), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n925), .B1(new_n963), .B2(KEYINPUT109), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT110), .B(G2090), .Z(new_n966));
  NAND3_X1  g541(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n920), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n940), .A3(new_n924), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n965), .A2(new_n966), .B1(new_n969), .B2(G1971), .ZN(new_n970));
  NAND2_X1  g545(.A1(G303), .A2(G8), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT55), .Z(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(G8), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n969), .A2(G1971), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n922), .A2(KEYINPUT50), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n940), .A3(new_n963), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(new_n966), .ZN(new_n977));
  OAI21_X1  g552(.A(G8), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n972), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n946), .A2(new_n957), .A3(new_n973), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n968), .A2(G2078), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n982), .A2(KEYINPUT53), .ZN(new_n983));
  INV_X1    g558(.A(G1961), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n965), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(KEYINPUT53), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(G301), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G2084), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n961), .B(new_n958), .C1(new_n921), .C2(new_n504), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n964), .A2(new_n993), .A3(new_n994), .A4(new_n975), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n962), .A2(KEYINPUT113), .A3(new_n993), .A4(new_n964), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n968), .A2(new_n785), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT120), .B1(G168), .B2(new_n950), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G286), .A2(new_n1002), .A3(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT122), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1001), .A2(new_n1008), .A3(new_n1003), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT121), .B1(new_n1000), .B2(G8), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT123), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1000), .A2(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1004), .A2(KEYINPUT51), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1014), .A2(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT124), .B(new_n1006), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT124), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1019), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1021), .B1(new_n1024), .B2(new_n1005), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n992), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT125), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT125), .B(new_n992), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1029));
  XOR2_X1   g604(.A(G299), .B(KEYINPUT117), .Z(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n563), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1030), .B(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT115), .B(G1956), .Z(new_n1034));
  NAND2_X1  g609(.A1(new_n976), .A2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT56), .B(G2072), .Z(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n968), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n962), .A2(new_n964), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1040), .A2(G1348), .B1(G2067), .B2(new_n941), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(new_n601), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(new_n1038), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1041), .A2(new_n601), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT60), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  OR3_X1    g623(.A1(new_n1041), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1039), .A2(KEYINPUT61), .A3(new_n1038), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT58), .B(G1341), .ZN(new_n1052));
  OAI22_X1  g627(.A1(G1996), .A2(new_n968), .B1(new_n949), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT118), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n552), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1038), .B(new_n1043), .C1(new_n1051), .C2(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1028), .A2(new_n1029), .A3(new_n1059), .ZN(new_n1060));
  AOI211_X1 g635(.A(G1976), .B(G288), .C1(new_n948), .C2(new_n951), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n583), .A2(new_n681), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n951), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n945), .A2(new_n956), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT112), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(new_n973), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n972), .B1(new_n970), .B2(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n973), .A2(KEYINPUT63), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1016), .A2(G286), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1071), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n981), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1070), .A2(new_n1071), .B1(KEYINPUT114), .B2(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1074), .A2(KEYINPUT114), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1067), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT62), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n987), .A2(G171), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n981), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1020), .A2(new_n1025), .A3(KEYINPUT62), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1077), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n938), .B1(new_n1060), .B2(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n928), .A2(KEYINPUT48), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n928), .A2(KEYINPUT48), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n937), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n713), .A2(new_n714), .A3(new_n719), .A4(new_n715), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n935), .A2(new_n1088), .B1(G2067), .B2(new_n759), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n926), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT47), .ZN(new_n1091));
  INV_X1    g666(.A(new_n932), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n926), .B1(new_n1092), .B2(new_n779), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n926), .A2(KEYINPUT46), .A3(new_n933), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT46), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n927), .B2(G1996), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1087), .B(new_n1090), .C1(new_n1091), .C2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1084), .A2(new_n1099), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g675(.A(KEYINPUT127), .ZN(new_n1102));
  OAI21_X1  g676(.A(G319), .B1(new_n650), .B2(new_n651), .ZN(new_n1103));
  NOR2_X1   g677(.A1(new_n1103), .A2(G227), .ZN(new_n1104));
  OAI21_X1  g678(.A(new_n1104), .B1(new_n683), .B2(new_n684), .ZN(new_n1105));
  XOR2_X1   g679(.A(new_n1105), .B(KEYINPUT126), .Z(new_n1106));
  NOR2_X1   g680(.A1(new_n1106), .A2(new_n841), .ZN(new_n1107));
  AND3_X1   g681(.A1(new_n913), .A2(new_n1102), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g682(.A(new_n1102), .B1(new_n913), .B2(new_n1107), .ZN(new_n1109));
  NOR2_X1   g683(.A1(new_n1108), .A2(new_n1109), .ZN(G308));
  NAND2_X1  g684(.A1(new_n913), .A2(new_n1107), .ZN(G225));
endmodule


