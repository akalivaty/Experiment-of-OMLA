

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U551 ( .A1(n541), .A2(G2104), .ZN(n886) );
  NOR2_X1 U552 ( .A1(n762), .A2(KEYINPUT33), .ZN(n764) );
  XNOR2_X1 U553 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U554 ( .A(KEYINPUT98), .B(n748), .ZN(n519) );
  AND2_X1 U555 ( .A1(G8), .A2(n750), .ZN(n520) );
  XOR2_X1 U556 ( .A(n708), .B(KEYINPUT31), .Z(n521) );
  XNOR2_X1 U557 ( .A(n749), .B(KEYINPUT93), .ZN(n697) );
  INV_X1 U558 ( .A(KEYINPUT101), .ZN(n763) );
  NAND2_X1 U559 ( .A1(n778), .A2(n776), .ZN(n739) );
  XNOR2_X1 U560 ( .A(n690), .B(KEYINPUT85), .ZN(n776) );
  NOR2_X1 U561 ( .A1(n545), .A2(n544), .ZN(G160) );
  XNOR2_X1 U562 ( .A(KEYINPUT7), .B(KEYINPUT74), .ZN(n536) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U564 ( .A1(n645), .A2(G89), .ZN(n522) );
  XNOR2_X1 U565 ( .A(n522), .B(KEYINPUT4), .ZN(n524) );
  XOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .Z(n638) );
  XNOR2_X1 U567 ( .A(G651), .B(KEYINPUT65), .ZN(n526) );
  NOR2_X1 U568 ( .A1(n638), .A2(n526), .ZN(n644) );
  NAND2_X1 U569 ( .A1(G76), .A2(n644), .ZN(n523) );
  NAND2_X1 U570 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U571 ( .A(KEYINPUT5), .B(n525), .ZN(n534) );
  NOR2_X1 U572 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n527), .Z(n652) );
  NAND2_X1 U574 ( .A1(n652), .A2(G63), .ZN(n528) );
  XOR2_X1 U575 ( .A(KEYINPUT73), .B(n528), .Z(n531) );
  NOR2_X1 U576 ( .A1(G651), .A2(n638), .ZN(n529) );
  XNOR2_X1 U577 ( .A(KEYINPUT64), .B(n529), .ZN(n648) );
  NAND2_X1 U578 ( .A1(G51), .A2(n648), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U580 ( .A(KEYINPUT6), .B(n532), .Z(n533) );
  NAND2_X1 U581 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U582 ( .A(n536), .B(n535), .ZN(G168) );
  XOR2_X1 U583 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  XOR2_X2 U585 ( .A(KEYINPUT17), .B(n537), .Z(n885) );
  NAND2_X1 U586 ( .A1(n885), .A2(G137), .ZN(n540) );
  INV_X1 U587 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U588 ( .A1(G101), .A2(n886), .ZN(n538) );
  XOR2_X1 U589 ( .A(n538), .B(KEYINPUT23), .Z(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n545) );
  AND2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U592 ( .A1(G113), .A2(n889), .ZN(n543) );
  NOR2_X1 U593 ( .A1(G2104), .A2(n541), .ZN(n890) );
  NAND2_X1 U594 ( .A1(G125), .A2(n890), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U596 ( .A(G2451), .B(G2427), .ZN(n555) );
  XOR2_X1 U597 ( .A(KEYINPUT103), .B(G2443), .Z(n547) );
  XNOR2_X1 U598 ( .A(G2435), .B(G2438), .ZN(n546) );
  XNOR2_X1 U599 ( .A(n547), .B(n546), .ZN(n551) );
  XOR2_X1 U600 ( .A(G2454), .B(G2430), .Z(n549) );
  XNOR2_X1 U601 ( .A(G1341), .B(G1348), .ZN(n548) );
  XNOR2_X1 U602 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U603 ( .A(n551), .B(n550), .Z(n553) );
  XNOR2_X1 U604 ( .A(G2446), .B(KEYINPUT104), .ZN(n552) );
  XNOR2_X1 U605 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U606 ( .A(n555), .B(n554), .ZN(n556) );
  AND2_X1 U607 ( .A1(n556), .A2(G14), .ZN(G401) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U609 ( .A(G108), .ZN(G238) );
  INV_X1 U610 ( .A(G120), .ZN(G236) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  XOR2_X1 U612 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n558) );
  NAND2_X1 U613 ( .A1(G7), .A2(G661), .ZN(n557) );
  XOR2_X1 U614 ( .A(n558), .B(n557), .Z(n827) );
  INV_X1 U615 ( .A(n827), .ZN(G223) );
  INV_X1 U616 ( .A(G567), .ZN(n679) );
  NOR2_X1 U617 ( .A1(n679), .A2(G223), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n559), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U619 ( .A1(n652), .A2(G56), .ZN(n560) );
  XOR2_X1 U620 ( .A(KEYINPUT14), .B(n560), .Z(n566) );
  NAND2_X1 U621 ( .A1(n645), .A2(G81), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G68), .A2(n644), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT13), .B(n564), .Z(n565) );
  NOR2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G43), .A2(n648), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n992) );
  INV_X1 U629 ( .A(G860), .ZN(n598) );
  OR2_X1 U630 ( .A1(n992), .A2(n598), .ZN(G153) );
  NAND2_X1 U631 ( .A1(n645), .A2(G90), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT68), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G77), .A2(n644), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT9), .ZN(n574) );
  NAND2_X1 U636 ( .A1(G64), .A2(n652), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G52), .A2(n648), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT67), .B(n575), .ZN(n576) );
  NOR2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT69), .B(n578), .ZN(G301) );
  NAND2_X1 U642 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U643 ( .A1(G54), .A2(n648), .ZN(n585) );
  NAND2_X1 U644 ( .A1(G79), .A2(n644), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G66), .A2(n652), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n645), .A2(G92), .ZN(n581) );
  XOR2_X1 U648 ( .A(KEYINPUT72), .B(n581), .Z(n582) );
  NOR2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(KEYINPUT15), .B(n586), .ZN(n1003) );
  INV_X1 U652 ( .A(n1003), .ZN(n726) );
  INV_X1 U653 ( .A(G868), .ZN(n665) );
  NAND2_X1 U654 ( .A1(n726), .A2(n665), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G65), .A2(n652), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G53), .A2(n648), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G91), .A2(n645), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G78), .A2(n644), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n990) );
  XOR2_X1 U663 ( .A(n990), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U664 ( .A1(G286), .A2(n665), .ZN(n595) );
  XOR2_X1 U665 ( .A(KEYINPUT75), .B(n595), .Z(n597) );
  NOR2_X1 U666 ( .A1(G299), .A2(G868), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U668 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n599), .A2(n1003), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U671 ( .A1(n1003), .A2(G868), .ZN(n601) );
  NOR2_X1 U672 ( .A1(G559), .A2(n601), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT76), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n992), .A2(G868), .ZN(n603) );
  NOR2_X1 U675 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G123), .A2(n890), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n889), .A2(G111), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G135), .A2(n885), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G99), .A2(n886), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n945) );
  XNOR2_X1 U684 ( .A(G2096), .B(n945), .ZN(n612) );
  INV_X1 U685 ( .A(G2100), .ZN(n852) );
  NAND2_X1 U686 ( .A1(n612), .A2(n852), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G93), .A2(n645), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G80), .A2(n644), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U690 ( .A(KEYINPUT78), .B(n615), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G55), .A2(n648), .ZN(n616) );
  XOR2_X1 U692 ( .A(KEYINPUT79), .B(n616), .Z(n618) );
  NAND2_X1 U693 ( .A1(n652), .A2(G67), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U695 ( .A(KEYINPUT80), .B(n619), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n664) );
  NAND2_X1 U697 ( .A1(n1003), .A2(G559), .ZN(n662) );
  XOR2_X1 U698 ( .A(KEYINPUT77), .B(n992), .Z(n622) );
  XNOR2_X1 U699 ( .A(n662), .B(n622), .ZN(n623) );
  NOR2_X1 U700 ( .A1(G860), .A2(n623), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n664), .B(n624), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G88), .A2(n645), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G75), .A2(n644), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G62), .A2(n652), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G50), .A2(n648), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(G166) );
  INV_X1 U709 ( .A(G166), .ZN(G303) );
  NAND2_X1 U710 ( .A1(G86), .A2(n645), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G61), .A2(n652), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n644), .A2(G73), .ZN(n633) );
  XOR2_X1 U714 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G48), .A2(n648), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G87), .A2(n638), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U721 ( .A1(n652), .A2(n641), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G49), .A2(n648), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U724 ( .A1(n644), .A2(G72), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n645), .A2(G85), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n648), .A2(G47), .ZN(n649) );
  XOR2_X1 U728 ( .A(KEYINPUT66), .B(n649), .Z(n650) );
  NOR2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n652), .A2(G60), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(G290) );
  XOR2_X1 U732 ( .A(G303), .B(G305), .Z(n657) );
  XOR2_X1 U733 ( .A(KEYINPUT19), .B(G290), .Z(n655) );
  XNOR2_X1 U734 ( .A(G288), .B(n655), .ZN(n656) );
  XNOR2_X1 U735 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U736 ( .A(G299), .B(n658), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n992), .B(n664), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n660), .B(n659), .ZN(n834) );
  XOR2_X1 U739 ( .A(n834), .B(KEYINPUT81), .Z(n661) );
  XNOR2_X1 U740 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X1 U741 ( .A1(n663), .A2(n665), .ZN(n667) );
  AND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U743 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U750 ( .A1(G132), .A2(G82), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(KEYINPUT22), .ZN(n673) );
  XNOR2_X1 U752 ( .A(n673), .B(KEYINPUT82), .ZN(n674) );
  NOR2_X1 U753 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G96), .A2(n675), .ZN(n832) );
  NAND2_X1 U755 ( .A1(G2106), .A2(n832), .ZN(n676) );
  XNOR2_X1 U756 ( .A(n676), .B(KEYINPUT83), .ZN(n681) );
  NOR2_X1 U757 ( .A1(G236), .A2(G238), .ZN(n677) );
  NAND2_X1 U758 ( .A1(G69), .A2(n677), .ZN(n678) );
  NOR2_X1 U759 ( .A1(G237), .A2(n678), .ZN(n831) );
  NOR2_X1 U760 ( .A1(n679), .A2(n831), .ZN(n680) );
  NOR2_X1 U761 ( .A1(n681), .A2(n680), .ZN(G319) );
  INV_X1 U762 ( .A(G319), .ZN(n904) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U764 ( .A1(n904), .A2(n682), .ZN(n830) );
  NAND2_X1 U765 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U766 ( .A1(n889), .A2(G114), .ZN(n683) );
  XNOR2_X1 U767 ( .A(n683), .B(KEYINPUT84), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G138), .A2(n885), .ZN(n684) );
  NAND2_X1 U769 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U770 ( .A1(G102), .A2(n886), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G126), .A2(n890), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U773 ( .A1(n689), .A2(n688), .ZN(G164) );
  INV_X1 U774 ( .A(G301), .ZN(G171) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n778) );
  NAND2_X1 U776 ( .A1(G40), .A2(G160), .ZN(n690) );
  NAND2_X1 U777 ( .A1(G8), .A2(n739), .ZN(n772) );
  NOR2_X1 U778 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XOR2_X1 U779 ( .A(n691), .B(KEYINPUT24), .Z(n692) );
  XNOR2_X1 U780 ( .A(KEYINPUT92), .B(n692), .ZN(n693) );
  NOR2_X1 U781 ( .A1(n772), .A2(n693), .ZN(n768) );
  XOR2_X1 U782 ( .A(G1981), .B(G305), .Z(n987) );
  NOR2_X1 U783 ( .A1(G1976), .A2(G288), .ZN(n998) );
  NAND2_X1 U784 ( .A1(n998), .A2(KEYINPUT33), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n772), .A2(n694), .ZN(n695) );
  XOR2_X1 U786 ( .A(KEYINPUT102), .B(n695), .Z(n696) );
  NAND2_X1 U787 ( .A1(n987), .A2(n696), .ZN(n766) );
  XOR2_X1 U788 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n747) );
  NOR2_X1 U789 ( .A1(n739), .A2(G2084), .ZN(n749) );
  NAND2_X1 U790 ( .A1(G8), .A2(n697), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n772), .A2(G1966), .ZN(n698) );
  XNOR2_X1 U792 ( .A(n698), .B(KEYINPUT94), .ZN(n751) );
  NOR2_X1 U793 ( .A1(n699), .A2(n751), .ZN(n700) );
  XOR2_X1 U794 ( .A(KEYINPUT30), .B(n700), .Z(n701) );
  NOR2_X1 U795 ( .A1(G168), .A2(n701), .ZN(n707) );
  XNOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .ZN(n702) );
  XNOR2_X1 U797 ( .A(n702), .B(KEYINPUT95), .ZN(n911) );
  NOR2_X1 U798 ( .A1(n911), .A2(n739), .ZN(n703) );
  XOR2_X1 U799 ( .A(KEYINPUT96), .B(n703), .Z(n705) );
  INV_X1 U800 ( .A(G1961), .ZN(n838) );
  NAND2_X1 U801 ( .A1(n739), .A2(n838), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n735) );
  NOR2_X1 U803 ( .A1(G171), .A2(n735), .ZN(n706) );
  NOR2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n708) );
  INV_X1 U805 ( .A(KEYINPUT29), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n739), .A2(G1956), .ZN(n711) );
  INV_X1 U807 ( .A(n739), .ZN(n720) );
  NAND2_X1 U808 ( .A1(n720), .A2(G2072), .ZN(n709) );
  XOR2_X1 U809 ( .A(KEYINPUT27), .B(n709), .Z(n710) );
  NAND2_X1 U810 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U811 ( .A(n712), .B(KEYINPUT97), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n990), .A2(n715), .ZN(n714) );
  INV_X1 U813 ( .A(KEYINPUT28), .ZN(n713) );
  XNOR2_X1 U814 ( .A(n714), .B(n713), .ZN(n732) );
  NAND2_X1 U815 ( .A1(n990), .A2(n715), .ZN(n730) );
  AND2_X1 U816 ( .A1(n720), .A2(G1996), .ZN(n716) );
  XOR2_X1 U817 ( .A(n716), .B(KEYINPUT26), .Z(n718) );
  NAND2_X1 U818 ( .A1(n739), .A2(G1341), .ZN(n717) );
  NAND2_X1 U819 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U820 ( .A1(n992), .A2(n719), .ZN(n724) );
  NAND2_X1 U821 ( .A1(G1348), .A2(n739), .ZN(n722) );
  NAND2_X1 U822 ( .A1(G2067), .A2(n720), .ZN(n721) );
  NAND2_X1 U823 ( .A1(n722), .A2(n721), .ZN(n725) );
  NOR2_X1 U824 ( .A1(n726), .A2(n725), .ZN(n723) );
  OR2_X1 U825 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U826 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U827 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U828 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U829 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U830 ( .A(n734), .B(n733), .ZN(n737) );
  NAND2_X1 U831 ( .A1(G171), .A2(n735), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U833 ( .A1(n521), .A2(n738), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n748), .A2(G286), .ZN(n744) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n772), .ZN(n741) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U837 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U838 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U840 ( .A1(G8), .A2(n745), .ZN(n746) );
  XNOR2_X1 U841 ( .A(n747), .B(n746), .ZN(n754) );
  XOR2_X1 U842 ( .A(KEYINPUT93), .B(n749), .Z(n750) );
  NOR2_X1 U843 ( .A1(n751), .A2(n520), .ZN(n752) );
  NAND2_X1 U844 ( .A1(n519), .A2(n752), .ZN(n753) );
  NAND2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n771) );
  INV_X1 U846 ( .A(n998), .ZN(n757) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n755) );
  XOR2_X1 U848 ( .A(n755), .B(KEYINPUT100), .Z(n756) );
  AND2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n771), .A2(n758), .ZN(n761) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n995) );
  INV_X1 U852 ( .A(n995), .ZN(n759) );
  NOR2_X1 U853 ( .A1(n759), .A2(n772), .ZN(n760) );
  AND2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n811) );
  INV_X1 U862 ( .A(n776), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n822) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(KEYINPUT91), .Z(n780) );
  NAND2_X1 U865 ( .A1(G105), .A2(n886), .ZN(n779) );
  XNOR2_X1 U866 ( .A(n780), .B(n779), .ZN(n787) );
  NAND2_X1 U867 ( .A1(G117), .A2(n889), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G141), .A2(n885), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n890), .A2(G129), .ZN(n783) );
  XOR2_X1 U871 ( .A(KEYINPUT90), .B(n783), .Z(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n869) );
  AND2_X1 U874 ( .A1(n869), .A2(G1996), .ZN(n946) );
  NAND2_X1 U875 ( .A1(G131), .A2(n885), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G119), .A2(n890), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G107), .A2(n889), .ZN(n790) );
  XNOR2_X1 U879 ( .A(KEYINPUT89), .B(n790), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n886), .A2(G95), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n868) );
  AND2_X1 U883 ( .A1(n868), .A2(G1991), .ZN(n938) );
  OR2_X1 U884 ( .A1(n946), .A2(n938), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n822), .A2(n795), .ZN(n812) );
  NAND2_X1 U886 ( .A1(G140), .A2(n885), .ZN(n797) );
  NAND2_X1 U887 ( .A1(G104), .A2(n886), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n798), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n889), .A2(G116), .ZN(n799) );
  XNOR2_X1 U891 ( .A(n799), .B(KEYINPUT86), .ZN(n801) );
  NAND2_X1 U892 ( .A1(G128), .A2(n890), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U894 ( .A(KEYINPUT35), .B(n802), .Z(n803) );
  NOR2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT36), .B(n805), .Z(n898) );
  XOR2_X1 U897 ( .A(KEYINPUT37), .B(G2067), .Z(n820) );
  NAND2_X1 U898 ( .A1(n898), .A2(n820), .ZN(n806) );
  XNOR2_X1 U899 ( .A(KEYINPUT87), .B(n806), .ZN(n936) );
  NAND2_X1 U900 ( .A1(n936), .A2(n822), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n807), .B(KEYINPUT88), .ZN(n818) );
  NAND2_X1 U902 ( .A1(n812), .A2(n818), .ZN(n809) );
  XNOR2_X1 U903 ( .A(G1986), .B(G290), .ZN(n1000) );
  AND2_X1 U904 ( .A1(n1000), .A2(n822), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n825) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n869), .ZN(n942) );
  INV_X1 U908 ( .A(n812), .ZN(n815) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n868), .ZN(n937) );
  NOR2_X1 U911 ( .A1(n813), .A2(n937), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U913 ( .A1(n942), .A2(n816), .ZN(n817) );
  XNOR2_X1 U914 ( .A(KEYINPUT39), .B(n817), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n821) );
  OR2_X1 U916 ( .A1(n898), .A2(n820), .ZN(n933) );
  NAND2_X1 U917 ( .A1(n821), .A2(n933), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U923 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U927 ( .A(G132), .ZN(G219) );
  INV_X1 U928 ( .A(G82), .ZN(G220) );
  INV_X1 U929 ( .A(n831), .ZN(n833) );
  NOR2_X1 U930 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XOR2_X1 U932 ( .A(n834), .B(n1003), .Z(n835) );
  XNOR2_X1 U933 ( .A(n835), .B(G286), .ZN(n836) );
  XOR2_X1 U934 ( .A(n836), .B(G301), .Z(n837) );
  NOR2_X1 U935 ( .A1(G37), .A2(n837), .ZN(G397) );
  XNOR2_X1 U936 ( .A(G1991), .B(G2474), .ZN(n848) );
  XNOR2_X1 U937 ( .A(G1956), .B(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1966), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(G1976), .B(G1981), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1971), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G229) );
  XNOR2_X1 U947 ( .A(G2072), .B(G2090), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n849), .B(KEYINPUT43), .ZN(n860) );
  XOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .Z(n851) );
  XNOR2_X1 U950 ( .A(KEYINPUT106), .B(G2096), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n856) );
  XNOR2_X1 U952 ( .A(n852), .B(G2084), .ZN(n854) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2078), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U955 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U956 ( .A(KEYINPUT105), .B(KEYINPUT107), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(G227) );
  NAND2_X1 U959 ( .A1(G124), .A2(n890), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n889), .A2(G112), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U963 ( .A1(G136), .A2(n885), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G100), .A2(n886), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(G162) );
  XNOR2_X1 U967 ( .A(n945), .B(n868), .ZN(n871) );
  XOR2_X1 U968 ( .A(G164), .B(n869), .Z(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n884) );
  XOR2_X1 U970 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n882) );
  NAND2_X1 U971 ( .A1(G118), .A2(n889), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G130), .A2(n890), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G142), .A2(n885), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G106), .A2(n886), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(KEYINPUT45), .B(n876), .ZN(n877) );
  XNOR2_X1 U978 ( .A(KEYINPUT109), .B(n877), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U980 ( .A(G162), .B(n880), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n884), .B(n883), .Z(n897) );
  NAND2_X1 U983 ( .A1(G139), .A2(n885), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U986 ( .A1(G115), .A2(n889), .ZN(n892) );
  NAND2_X1 U987 ( .A1(G127), .A2(n890), .ZN(n891) );
  NAND2_X1 U988 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U990 ( .A1(n895), .A2(n894), .ZN(n929) );
  XNOR2_X1 U991 ( .A(G160), .B(n929), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G37), .A2(n900), .ZN(G395) );
  NOR2_X1 U995 ( .A1(G229), .A2(G227), .ZN(n901) );
  XOR2_X1 U996 ( .A(KEYINPUT49), .B(n901), .Z(n902) );
  XNOR2_X1 U997 ( .A(n902), .B(KEYINPUT111), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G397), .A2(n903), .ZN(n908) );
  NOR2_X1 U999 ( .A1(n904), .A2(G401), .ZN(n905) );
  XOR2_X1 U1000 ( .A(KEYINPUT110), .B(n905), .Z(n906) );
  NOR2_X1 U1001 ( .A1(G395), .A2(n906), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(G69), .ZN(G235) );
  INV_X1 U1005 ( .A(G96), .ZN(G221) );
  INV_X1 U1006 ( .A(KEYINPUT55), .ZN(n955) );
  XNOR2_X1 U1007 ( .A(G2067), .B(G26), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(G32), .B(G1996), .ZN(n909) );
  NOR2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(n911), .B(G27), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(G2072), .B(G33), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(G1991), .B(G25), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(KEYINPUT115), .ZN(n917) );
  NAND2_X1 U1016 ( .A1(G28), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(KEYINPUT116), .B(n918), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1019 ( .A(KEYINPUT53), .B(n921), .Z(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT54), .B(G34), .Z(n922) );
  XNOR2_X1 U1021 ( .A(G2084), .B(n922), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(G35), .B(G2090), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n955), .B(n927), .ZN(n928) );
  NOR2_X1 U1026 ( .A1(G29), .A2(n928), .ZN(n960) );
  XOR2_X1 U1027 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(n932), .B(KEYINPUT50), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n952) );
  XNOR2_X1 U1033 ( .A(G160), .B(G2084), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n950) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1038 ( .A(KEYINPUT112), .B(n943), .Z(n944) );
  XNOR2_X1 U1039 ( .A(KEYINPUT51), .B(n944), .ZN(n948) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(KEYINPUT113), .B(n953), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(n954), .ZN(n956) );
  NAND2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1047 ( .A1(n957), .A2(G29), .ZN(n958) );
  XOR2_X1 U1048 ( .A(KEYINPUT114), .B(n958), .Z(n959) );
  NOR2_X1 U1049 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1050 ( .A1(G11), .A2(n961), .ZN(n1019) );
  XOR2_X1 U1051 ( .A(G1971), .B(G22), .Z(n964) );
  XOR2_X1 U1052 ( .A(G23), .B(KEYINPUT124), .Z(n962) );
  XNOR2_X1 U1053 ( .A(n962), .B(G1976), .ZN(n963) );
  NAND2_X1 U1054 ( .A1(n964), .A2(n963), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(G24), .B(G1986), .ZN(n965) );
  NOR2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1057 ( .A(KEYINPUT58), .B(n967), .Z(n984) );
  XOR2_X1 U1058 ( .A(G1966), .B(G21), .Z(n969) );
  XOR2_X1 U1059 ( .A(G1961), .B(G5), .Z(n968) );
  NAND2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n981) );
  XNOR2_X1 U1061 ( .A(KEYINPUT59), .B(G1348), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n970), .B(G4), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(G1956), .B(G20), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G6), .B(G1981), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT121), .B(n973), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT60), .B(n978), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(KEYINPUT122), .B(n979), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT123), .B(n982), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1075 ( .A(KEYINPUT61), .B(n985), .Z(n986) );
  NOR2_X1 U1076 ( .A1(G16), .A2(n986), .ZN(n1016) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n989), .Z(n1010) );
  XOR2_X1 U1080 ( .A(n990), .B(G1956), .Z(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT118), .B(n991), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n1007) );
  XOR2_X1 U1086 ( .A(G301), .B(G1961), .Z(n1002) );
  XOR2_X1 U1087 ( .A(G1971), .B(G166), .Z(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1090 ( .A(G1348), .B(n1003), .Z(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1093 ( .A(KEYINPUT119), .B(n1008), .Z(n1009) );
  NOR2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(G16), .B(KEYINPUT117), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(KEYINPUT56), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(n1014), .B(KEYINPUT120), .ZN(n1015) );
  NOR2_X1 U1099 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(n1017), .B(KEYINPUT125), .ZN(n1018) );
  NOR2_X1 U1101 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1020), .ZN(G311) );
  XOR2_X1 U1103 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

