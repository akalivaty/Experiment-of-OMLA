

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U325 ( .A(n337), .B(n336), .ZN(n342) );
  XNOR2_X1 U326 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U327 ( .A(n421), .B(n396), .Z(n293) );
  NOR2_X1 U328 ( .A1(n570), .A2(n569), .ZN(n294) );
  XOR2_X1 U329 ( .A(G71GAT), .B(G78GAT), .Z(n295) );
  NOR2_X1 U330 ( .A1(n567), .A2(n494), .ZN(n344) );
  XNOR2_X1 U331 ( .A(n349), .B(n295), .ZN(n316) );
  XNOR2_X1 U332 ( .A(n316), .B(n315), .ZN(n318) );
  XNOR2_X1 U333 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U334 ( .A(n329), .B(n328), .ZN(n481) );
  XNOR2_X1 U335 ( .A(n343), .B(n293), .ZN(n383) );
  XNOR2_X1 U336 ( .A(n462), .B(KEYINPUT123), .ZN(n584) );
  XNOR2_X1 U337 ( .A(n456), .B(G176GAT), .ZN(n457) );
  XNOR2_X1 U338 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U339 ( .A(G176GAT), .B(G64GAT), .Z(n348) );
  XOR2_X1 U340 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n297) );
  XNOR2_X1 U341 ( .A(G204GAT), .B(G92GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U343 ( .A(n348), .B(n298), .Z(n300) );
  NAND2_X1 U344 ( .A1(G226GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U346 ( .A(G8GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n301), .B(KEYINPUT79), .ZN(n317) );
  XOR2_X1 U348 ( .A(n302), .B(n317), .Z(n308) );
  XOR2_X1 U349 ( .A(KEYINPUT21), .B(KEYINPUT92), .Z(n304) );
  XNOR2_X1 U350 ( .A(KEYINPUT91), .B(G211GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U352 ( .A(G197GAT), .B(n305), .ZN(n433) );
  XNOR2_X1 U353 ( .A(G36GAT), .B(G190GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n306), .B(G218GAT), .ZN(n340) );
  XOR2_X1 U355 ( .A(n433), .B(n340), .Z(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U357 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n310) );
  XNOR2_X1 U358 ( .A(KEYINPUT17), .B(KEYINPUT87), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(n311), .ZN(n451) );
  XOR2_X1 U361 ( .A(n312), .B(n451), .Z(n526) );
  INV_X1 U362 ( .A(n526), .ZN(n514) );
  XOR2_X1 U363 ( .A(G57GAT), .B(KEYINPUT13), .Z(n349) );
  XOR2_X1 U364 ( .A(KEYINPUT80), .B(G64GAT), .Z(n314) );
  XNOR2_X1 U365 ( .A(G211GAT), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U367 ( .A(n318), .B(n317), .Z(n320) );
  XOR2_X1 U368 ( .A(G22GAT), .B(G1GAT), .Z(n365) );
  XOR2_X1 U369 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XNOR2_X1 U370 ( .A(n365), .B(n442), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n329) );
  XOR2_X1 U372 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n322) );
  XNOR2_X1 U373 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n323), .B(KEYINPUT15), .ZN(n327) );
  XOR2_X1 U376 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n325) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  INV_X1 U379 ( .A(n481), .ZN(n567) );
  XOR2_X1 U380 ( .A(G29GAT), .B(G43GAT), .Z(n331) );
  XNOR2_X1 U381 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n366) );
  XNOR2_X1 U383 ( .A(KEYINPUT76), .B(n366), .ZN(n337) );
  XOR2_X1 U384 ( .A(KEYINPUT11), .B(KEYINPUT67), .Z(n333) );
  XNOR2_X1 U385 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n332) );
  XOR2_X1 U386 ( .A(n333), .B(n332), .Z(n335) );
  AND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n334) );
  XOR2_X1 U388 ( .A(G92GAT), .B(G85GAT), .Z(n339) );
  XNOR2_X1 U389 ( .A(G99GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n347) );
  XNOR2_X1 U391 ( .A(n340), .B(n347), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U393 ( .A(G50GAT), .B(G162GAT), .Z(n421) );
  XOR2_X1 U394 ( .A(G134GAT), .B(KEYINPUT77), .Z(n396) );
  XOR2_X1 U395 ( .A(n383), .B(KEYINPUT78), .Z(n570) );
  XNOR2_X1 U396 ( .A(KEYINPUT36), .B(n570), .ZN(n494) );
  XNOR2_X1 U397 ( .A(n344), .B(KEYINPUT45), .ZN(n363) );
  XOR2_X1 U398 ( .A(G78GAT), .B(G148GAT), .Z(n346) );
  XNOR2_X1 U399 ( .A(KEYINPUT72), .B(G204GAT), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n428) );
  XNOR2_X1 U401 ( .A(n428), .B(n347), .ZN(n362) );
  XOR2_X1 U402 ( .A(n349), .B(n348), .Z(n351) );
  NAND2_X1 U403 ( .A1(G230GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(KEYINPUT74), .Z(n353) );
  XNOR2_X1 U406 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U408 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U409 ( .A(G120GAT), .B(G71GAT), .Z(n450) );
  XOR2_X1 U410 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n357) );
  XNOR2_X1 U411 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n450), .B(n358), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U415 ( .A(n362), .B(n361), .Z(n579) );
  AND2_X1 U416 ( .A1(n363), .A2(n579), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n364), .B(KEYINPUT116), .ZN(n381) );
  XOR2_X1 U418 ( .A(n366), .B(n365), .Z(n368) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U421 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n370) );
  XNOR2_X1 U422 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U424 ( .A(n372), .B(n371), .Z(n380) );
  XOR2_X1 U425 ( .A(G15GAT), .B(G113GAT), .Z(n374) );
  XNOR2_X1 U426 ( .A(G50GAT), .B(G36GAT), .ZN(n373) );
  XNOR2_X1 U427 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U428 ( .A(G8GAT), .B(G141GAT), .Z(n376) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(G197GAT), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U432 ( .A(n380), .B(n379), .Z(n509) );
  INV_X1 U433 ( .A(n509), .ZN(n575) );
  NAND2_X1 U434 ( .A1(n381), .A2(n575), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n382), .B(KEYINPUT117), .ZN(n391) );
  XOR2_X1 U436 ( .A(KEYINPUT47), .B(KEYINPUT115), .Z(n389) );
  BUF_X1 U437 ( .A(n383), .Z(n560) );
  XNOR2_X1 U438 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n384) );
  XOR2_X1 U439 ( .A(n579), .B(n384), .Z(n556) );
  NOR2_X1 U440 ( .A1(n575), .A2(n556), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n385), .B(KEYINPUT46), .ZN(n386) );
  NOR2_X1 U442 ( .A1(n560), .A2(n386), .ZN(n387) );
  NAND2_X1 U443 ( .A1(n387), .A2(n567), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  NOR2_X1 U445 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n392), .B(KEYINPUT48), .ZN(n536) );
  NOR2_X1 U447 ( .A1(n514), .A2(n536), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n393), .B(KEYINPUT54), .ZN(n416) );
  XOR2_X1 U449 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n395) );
  XNOR2_X1 U450 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n400) );
  XOR2_X1 U452 ( .A(G85GAT), .B(n396), .Z(n398) );
  XOR2_X1 U453 ( .A(G113GAT), .B(KEYINPUT0), .Z(n445) );
  XNOR2_X1 U454 ( .A(G29GAT), .B(n445), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U456 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U459 ( .A(n403), .B(KEYINPUT6), .Z(n407) );
  XOR2_X1 U460 ( .A(G155GAT), .B(KEYINPUT2), .Z(n405) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n427) );
  XNOR2_X1 U463 ( .A(n427), .B(KEYINPUT97), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n415) );
  XOR2_X1 U465 ( .A(KEYINPUT1), .B(G57GAT), .Z(n409) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U468 ( .A(G162GAT), .B(G148GAT), .Z(n411) );
  XNOR2_X1 U469 ( .A(G120GAT), .B(G127GAT), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U471 ( .A(n413), .B(n412), .Z(n414) );
  XOR2_X1 U472 ( .A(n415), .B(n414), .Z(n524) );
  INV_X1 U473 ( .A(n524), .ZN(n511) );
  NAND2_X1 U474 ( .A1(n416), .A2(n511), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n417), .B(KEYINPUT65), .ZN(n461) );
  XOR2_X1 U476 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n419) );
  XNOR2_X1 U477 ( .A(G218GAT), .B(G106GAT), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U479 ( .A(n420), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U480 ( .A(G22GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n432) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n425) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U485 ( .A(n426), .B(KEYINPUT90), .Z(n430) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n435) );
  INV_X1 U489 ( .A(n433), .ZN(n434) );
  XOR2_X1 U490 ( .A(n435), .B(n434), .Z(n475) );
  NAND2_X1 U491 ( .A1(n461), .A2(n475), .ZN(n436) );
  XNOR2_X1 U492 ( .A(KEYINPUT55), .B(n436), .ZN(n571) );
  XOR2_X1 U493 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n438) );
  XNOR2_X1 U494 ( .A(G176GAT), .B(KEYINPUT66), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n455) );
  XOR2_X1 U496 ( .A(KEYINPUT20), .B(G183GAT), .Z(n440) );
  XNOR2_X1 U497 ( .A(G134GAT), .B(G190GAT), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U499 ( .A(n441), .B(G99GAT), .Z(n444) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n449) );
  XOR2_X1 U502 ( .A(n445), .B(KEYINPUT85), .Z(n447) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U505 ( .A(n449), .B(n448), .Z(n453) );
  XOR2_X1 U506 ( .A(n451), .B(n450), .Z(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n569) );
  INV_X1 U509 ( .A(n569), .ZN(n540) );
  NAND2_X1 U510 ( .A1(n571), .A2(n540), .ZN(n566) );
  XNOR2_X1 U511 ( .A(n556), .B(KEYINPUT110), .ZN(n542) );
  NOR2_X1 U512 ( .A1(n566), .A2(n542), .ZN(n458) );
  XNOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n456) );
  NOR2_X1 U514 ( .A1(n540), .A2(n475), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT101), .B(n459), .Z(n460) );
  XNOR2_X1 U516 ( .A(KEYINPUT26), .B(n460), .ZN(n551) );
  AND2_X1 U517 ( .A1(n551), .A2(n461), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n567), .A2(n584), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT126), .ZN(n465) );
  INV_X1 U520 ( .A(G211GAT), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(G1354GAT) );
  INV_X1 U522 ( .A(n579), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n575), .A2(n466), .ZN(n498) );
  NAND2_X1 U524 ( .A1(n526), .A2(n540), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n467), .A2(n475), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT102), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n469), .Z(n471) );
  XNOR2_X1 U528 ( .A(n526), .B(KEYINPUT27), .ZN(n474) );
  NAND2_X1 U529 ( .A1(n474), .A2(n551), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n511), .A2(n472), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT103), .ZN(n479) );
  NAND2_X1 U533 ( .A1(n524), .A2(n474), .ZN(n535) );
  XNOR2_X1 U534 ( .A(KEYINPUT28), .B(n475), .ZN(n538) );
  INV_X1 U535 ( .A(n538), .ZN(n531) );
  NOR2_X1 U536 ( .A1(n535), .A2(n531), .ZN(n476) );
  XOR2_X1 U537 ( .A(KEYINPUT100), .B(n476), .Z(n477) );
  NOR2_X1 U538 ( .A1(n477), .A2(n540), .ZN(n478) );
  NOR2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U540 ( .A(KEYINPUT104), .B(n480), .ZN(n495) );
  NAND2_X1 U541 ( .A1(n481), .A2(n570), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT16), .B(n482), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n495), .A2(n483), .ZN(n510) );
  NAND2_X1 U544 ( .A1(n498), .A2(n510), .ZN(n492) );
  NOR2_X1 U545 ( .A1(n511), .A2(n492), .ZN(n485) );
  XNOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT105), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n514), .A2(n492), .ZN(n487) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n487), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n492), .A2(n569), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n489) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n538), .A2(n492), .ZN(n493) );
  XOR2_X1 U557 ( .A(G22GAT), .B(n493), .Z(G1327GAT) );
  BUF_X1 U558 ( .A(n494), .Z(n585) );
  NOR2_X1 U559 ( .A1(n585), .A2(n495), .ZN(n496) );
  NAND2_X1 U560 ( .A1(n496), .A2(n567), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(KEYINPUT37), .ZN(n521) );
  NAND2_X1 U562 ( .A1(n498), .A2(n521), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT38), .ZN(n505) );
  NOR2_X1 U564 ( .A1(n505), .A2(n511), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n514), .A2(n505), .ZN(n502) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U569 ( .A1(n505), .A2(n569), .ZN(n503) );
  XOR2_X1 U570 ( .A(KEYINPUT40), .B(n503), .Z(n504) );
  XNOR2_X1 U571 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  XNOR2_X1 U572 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n507) );
  NOR2_X1 U573 ( .A1(n538), .A2(n505), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  NOR2_X1 U576 ( .A1(n509), .A2(n542), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n522), .A2(n510), .ZN(n518) );
  NOR2_X1 U578 ( .A1(n511), .A2(n518), .ZN(n512) );
  XOR2_X1 U579 ( .A(G57GAT), .B(n512), .Z(n513) );
  XNOR2_X1 U580 ( .A(KEYINPUT42), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n518), .ZN(n515) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n569), .A2(n518), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  NOR2_X1 U586 ( .A1(n538), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U590 ( .A(KEYINPUT112), .B(n523), .Z(n532) );
  NAND2_X1 U591 ( .A1(n532), .A2(n524), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U593 ( .A(G92GAT), .B(KEYINPUT113), .Z(n528) );
  NAND2_X1 U594 ( .A1(n532), .A2(n526), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n540), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n529), .B(KEYINPUT114), .ZN(n530) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  NAND2_X1 U599 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n533), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT118), .B(n537), .ZN(n550) );
  AND2_X1 U604 ( .A1(n550), .A2(n538), .ZN(n539) );
  NAND2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n547) );
  NOR2_X1 U606 ( .A1(n575), .A2(n547), .ZN(n541) );
  XOR2_X1 U607 ( .A(G113GAT), .B(n541), .Z(G1340GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n547), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  NOR2_X1 U611 ( .A1(n567), .A2(n547), .ZN(n545) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(n545), .Z(n546) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  NOR2_X1 U614 ( .A1(n570), .A2(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n575), .A2(n561), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n556), .A2(n561), .ZN(n557) );
  XOR2_X1 U625 ( .A(n558), .B(n557), .Z(G1345GAT) );
  NOR2_X1 U626 ( .A1(n567), .A2(n561), .ZN(n559) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  INV_X1 U628 ( .A(n560), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NOR2_X1 U631 ( .A1(n575), .A2(n566), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  AND2_X1 U636 ( .A1(n571), .A2(n294), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(n574), .B(G190GAT), .Z(G1351GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n584), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n584), .A2(n579), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  INV_X1 U650 ( .A(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G218GAT), .ZN(G1355GAT) );
endmodule

