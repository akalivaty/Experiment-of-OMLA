

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749;

  NAND2_X1 U382 ( .A1(n547), .A2(n658), .ZN(n374) );
  XNOR2_X1 U383 ( .A(n480), .B(KEYINPUT10), .ZN(n733) );
  NAND2_X2 U384 ( .A1(n749), .A2(n746), .ZN(n606) );
  INV_X1 U385 ( .A(n608), .ZN(n393) );
  NOR2_X2 U386 ( .A1(n576), .A2(n654), .ZN(n582) );
  XNOR2_X2 U387 ( .A(n734), .B(n471), .ZN(n631) );
  XNOR2_X2 U388 ( .A(n530), .B(n531), .ZN(n571) );
  XNOR2_X2 U389 ( .A(n463), .B(G119), .ZN(n510) );
  XNOR2_X2 U390 ( .A(n539), .B(n538), .ZN(n570) );
  XNOR2_X2 U391 ( .A(n432), .B(KEYINPUT35), .ZN(n743) );
  XNOR2_X1 U392 ( .A(n496), .B(n495), .ZN(n672) );
  XNOR2_X1 U393 ( .A(G146), .B(G125), .ZN(n480) );
  AND2_X1 U394 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U395 ( .A(n431), .B(KEYINPUT67), .ZN(n604) );
  XNOR2_X1 U396 ( .A(n397), .B(n383), .ZN(n382) );
  NOR2_X2 U397 ( .A1(n672), .A2(n671), .ZN(n677) );
  NOR2_X2 U398 ( .A1(n542), .A2(n571), .ZN(n568) );
  XNOR2_X1 U399 ( .A(n537), .B(n385), .ZN(n707) );
  XNOR2_X1 U400 ( .A(n430), .B(G101), .ZN(n508) );
  NOR2_X2 U401 ( .A1(G902), .A2(n631), .ZN(n473) );
  XNOR2_X2 U402 ( .A(n396), .B(n395), .ZN(n734) );
  INV_X1 U403 ( .A(G134), .ZN(n454) );
  XNOR2_X1 U404 ( .A(KEYINPUT73), .B(G128), .ZN(n461) );
  XNOR2_X1 U405 ( .A(n508), .B(n429), .ZN(n466) );
  INV_X1 U406 ( .A(G110), .ZN(n429) );
  XNOR2_X1 U407 ( .A(n464), .B(KEYINPUT85), .ZN(n447) );
  NAND2_X1 U408 ( .A1(n627), .A2(n623), .ZN(n375) );
  XNOR2_X1 U409 ( .A(n414), .B(n511), .ZN(n514) );
  XOR2_X1 U410 ( .A(KEYINPUT65), .B(n625), .Z(n626) );
  AND2_X1 U411 ( .A1(n392), .A2(n381), .ZN(n380) );
  INV_X1 U412 ( .A(n365), .ZN(n381) );
  NAND2_X1 U413 ( .A1(n393), .A2(n363), .ZN(n392) );
  INV_X1 U414 ( .A(n671), .ZN(n398) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n534) );
  NOR2_X1 U416 ( .A1(n735), .A2(n623), .ZN(n449) );
  XOR2_X1 U417 ( .A(KEYINPUT84), .B(KEYINPUT18), .Z(n459) );
  XNOR2_X1 U418 ( .A(n480), .B(n428), .ZN(n427) );
  XNOR2_X1 U419 ( .A(KEYINPUT72), .B(KEYINPUT17), .ZN(n428) );
  INV_X1 U420 ( .A(KEYINPUT4), .ZN(n462) );
  OR2_X2 U421 ( .A1(n743), .A2(KEYINPUT44), .ZN(n431) );
  AND2_X1 U422 ( .A1(n442), .A2(n438), .ZN(n619) );
  XNOR2_X1 U423 ( .A(n419), .B(KEYINPUT46), .ZN(n418) );
  NOR2_X1 U424 ( .A1(n748), .A2(n747), .ZN(n419) );
  XNOR2_X1 U425 ( .A(G953), .B(KEYINPUT64), .ZN(n502) );
  XNOR2_X1 U426 ( .A(n404), .B(n402), .ZN(n721) );
  XNOR2_X1 U427 ( .A(n521), .B(n403), .ZN(n402) );
  XNOR2_X1 U428 ( .A(n510), .B(n535), .ZN(n404) );
  INV_X1 U429 ( .A(KEYINPUT16), .ZN(n403) );
  XNOR2_X1 U430 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U431 ( .A(n573), .B(n371), .ZN(n693) );
  INV_X1 U432 ( .A(n693), .ZN(n389) );
  XNOR2_X1 U433 ( .A(n413), .B(n412), .ZN(n567) );
  INV_X1 U434 ( .A(KEYINPUT39), .ZN(n412) );
  NOR2_X1 U435 ( .A1(n540), .A2(n572), .ZN(n413) );
  INV_X1 U436 ( .A(KEYINPUT34), .ZN(n409) );
  AND2_X1 U437 ( .A1(n382), .A2(n608), .ZN(n591) );
  INV_X1 U438 ( .A(KEYINPUT98), .ZN(n425) );
  INV_X1 U439 ( .A(KEYINPUT0), .ZN(n384) );
  NAND2_X1 U440 ( .A1(n713), .A2(n373), .ZN(n445) );
  NOR2_X1 U441 ( .A1(n444), .A2(n720), .ZN(n443) );
  NOR2_X1 U442 ( .A1(n372), .A2(G472), .ZN(n444) );
  INV_X1 U443 ( .A(n502), .ZN(n736) );
  XNOR2_X1 U444 ( .A(n423), .B(n422), .ZN(n537) );
  XNOR2_X1 U445 ( .A(n536), .B(n387), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U447 ( .A1(n405), .A2(n367), .ZN(n441) );
  INV_X1 U448 ( .A(KEYINPUT79), .ZN(n406) );
  INV_X1 U449 ( .A(KEYINPUT66), .ZN(n430) );
  INV_X1 U450 ( .A(KEYINPUT102), .ZN(n439) );
  NAND2_X1 U451 ( .A1(n441), .A2(n369), .ZN(n440) );
  XOR2_X1 U452 ( .A(G113), .B(KEYINPUT5), .Z(n507) );
  XNOR2_X1 U453 ( .A(n388), .B(G122), .ZN(n521) );
  INV_X1 U454 ( .A(G107), .ZN(n388) );
  XNOR2_X1 U455 ( .A(G146), .B(G104), .ZN(n468) );
  INV_X1 U456 ( .A(n485), .ZN(n395) );
  NAND2_X1 U457 ( .A1(n659), .A2(n658), .ZN(n663) );
  XNOR2_X1 U458 ( .A(n547), .B(n426), .ZN(n659) );
  INV_X1 U459 ( .A(KEYINPUT38), .ZN(n426) );
  XNOR2_X1 U460 ( .A(n379), .B(n378), .ZN(n668) );
  INV_X1 U461 ( .A(KEYINPUT33), .ZN(n378) );
  NAND2_X1 U462 ( .A1(n380), .A2(n394), .ZN(n379) );
  XNOR2_X1 U463 ( .A(n401), .B(G472), .ZN(n611) );
  INV_X1 U464 ( .A(KEYINPUT22), .ZN(n383) );
  XNOR2_X1 U465 ( .A(G128), .B(G110), .ZN(n486) );
  XNOR2_X1 U466 ( .A(n733), .B(n437), .ZN(n481) );
  XNOR2_X1 U467 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n437) );
  XOR2_X1 U468 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n479) );
  XOR2_X1 U469 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n484) );
  XNOR2_X1 U470 ( .A(KEYINPUT69), .B(G131), .ZN(n536) );
  XNOR2_X1 U471 ( .A(G143), .B(G140), .ZN(n387) );
  XNOR2_X1 U472 ( .A(n733), .B(n424), .ZN(n423) );
  XNOR2_X1 U473 ( .A(n532), .B(KEYINPUT96), .ZN(n424) );
  XNOR2_X1 U474 ( .A(G122), .B(KEYINPUT97), .ZN(n532) );
  XNOR2_X1 U475 ( .A(n533), .B(n455), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n377), .B(n376), .ZN(n627) );
  XNOR2_X1 U477 ( .A(n460), .B(n465), .ZN(n376) );
  XNOR2_X1 U478 ( .A(n721), .B(n364), .ZN(n377) );
  XNOR2_X1 U479 ( .A(n417), .B(KEYINPUT48), .ZN(n576) );
  XNOR2_X1 U480 ( .A(n494), .B(n456), .ZN(n495) );
  INV_X1 U481 ( .A(KEYINPUT103), .ZN(n416) );
  INV_X1 U482 ( .A(n611), .ZN(n592) );
  INV_X1 U483 ( .A(KEYINPUT1), .ZN(n557) );
  INV_X1 U484 ( .A(G953), .ZN(n583) );
  NAND2_X1 U485 ( .A1(n389), .A2(n574), .ZN(n575) );
  XNOR2_X1 U486 ( .A(n569), .B(n411), .ZN(n748) );
  INV_X1 U487 ( .A(KEYINPUT40), .ZN(n411) );
  XNOR2_X1 U488 ( .A(n560), .B(KEYINPUT108), .ZN(n744) );
  INV_X1 U489 ( .A(n603), .ZN(n407) );
  NAND2_X1 U490 ( .A1(n362), .A2(n366), .ZN(n400) );
  XNOR2_X1 U491 ( .A(n719), .B(n718), .ZN(n399) );
  XNOR2_X1 U492 ( .A(n717), .B(KEYINPUT126), .ZN(n718) );
  XNOR2_X1 U493 ( .A(n714), .B(n715), .ZN(n410) );
  NOR2_X1 U494 ( .A1(n710), .A2(n720), .ZN(n711) );
  XNOR2_X1 U495 ( .A(n633), .B(n632), .ZN(n634) );
  INV_X1 U496 ( .A(KEYINPUT56), .ZN(n433) );
  INV_X1 U497 ( .A(n441), .ZN(n636) );
  OR2_X1 U498 ( .A1(n713), .A2(n372), .ZN(n362) );
  AND2_X1 U499 ( .A1(n677), .A2(KEYINPUT105), .ZN(n363) );
  XOR2_X1 U500 ( .A(n466), .B(n427), .Z(n364) );
  XNOR2_X1 U501 ( .A(KEYINPUT6), .B(n592), .ZN(n365) );
  AND2_X1 U502 ( .A1(n445), .A2(n443), .ZN(n366) );
  AND2_X1 U503 ( .A1(n608), .A2(n607), .ZN(n367) );
  XOR2_X1 U504 ( .A(n536), .B(n454), .Z(n368) );
  OR2_X1 U505 ( .A1(n616), .A2(n615), .ZN(n369) );
  AND2_X1 U506 ( .A1(n590), .A2(n398), .ZN(n370) );
  XOR2_X1 U507 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n371) );
  XOR2_X1 U508 ( .A(n635), .B(KEYINPUT62), .Z(n372) );
  AND2_X1 U509 ( .A1(n372), .A2(G472), .ZN(n373) );
  NOR2_X1 U510 ( .A1(n736), .A2(G952), .ZN(n720) );
  INV_X1 U511 ( .A(n720), .ZN(n446) );
  XNOR2_X2 U512 ( .A(n374), .B(KEYINPUT19), .ZN(n587) );
  NOR2_X1 U513 ( .A1(n577), .A2(n374), .ZN(n556) );
  XNOR2_X2 U514 ( .A(n375), .B(n447), .ZN(n547) );
  INV_X1 U515 ( .A(n668), .ZN(n601) );
  AND2_X1 U516 ( .A1(n382), .A2(n365), .ZN(n609) );
  NAND2_X1 U517 ( .A1(n600), .A2(n370), .ZN(n397) );
  XNOR2_X2 U518 ( .A(n589), .B(n384), .ZN(n600) );
  XNOR2_X1 U519 ( .A(n535), .B(n386), .ZN(n385) );
  NAND2_X1 U520 ( .A1(n686), .A2(n389), .ZN(n687) );
  NAND2_X1 U521 ( .A1(n554), .A2(n649), .ZN(n577) );
  XNOR2_X2 U522 ( .A(n568), .B(KEYINPUT106), .ZN(n649) );
  XNOR2_X1 U523 ( .A(n570), .B(n425), .ZN(n542) );
  NAND2_X1 U524 ( .A1(n390), .A2(n599), .ZN(n394) );
  NAND2_X1 U525 ( .A1(n391), .A2(n677), .ZN(n390) );
  INV_X1 U526 ( .A(n608), .ZN(n391) );
  NAND2_X1 U527 ( .A1(n393), .A2(n677), .ZN(n610) );
  XNOR2_X1 U528 ( .A(n514), .B(n396), .ZN(n635) );
  XNOR2_X2 U529 ( .A(n465), .B(n368), .ZN(n396) );
  NOR2_X1 U530 ( .A1(n399), .A2(n720), .ZN(G66) );
  NAND2_X1 U531 ( .A1(n448), .A2(n626), .ZN(n704) );
  NAND2_X1 U532 ( .A1(n713), .A2(G210), .ZN(n436) );
  XNOR2_X1 U533 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U534 ( .A(n400), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U535 ( .A(n436), .B(n630), .ZN(n435) );
  NAND2_X1 U536 ( .A1(n435), .A2(n446), .ZN(n434) );
  NOR2_X1 U537 ( .A1(n614), .A2(n592), .ZN(n638) );
  NOR2_X1 U538 ( .A1(n635), .A2(G902), .ZN(n401) );
  XNOR2_X1 U539 ( .A(n512), .B(n513), .ZN(n414) );
  NAND2_X1 U540 ( .A1(n606), .A2(KEYINPUT44), .ZN(n442) );
  XNOR2_X1 U541 ( .A(n440), .B(n439), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n609), .B(n406), .ZN(n405) );
  XNOR2_X1 U543 ( .A(n602), .B(n409), .ZN(n408) );
  NAND2_X1 U544 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U545 ( .A1(n604), .A2(n605), .ZN(n621) );
  NAND2_X1 U546 ( .A1(n408), .A2(n407), .ZN(n432) );
  NAND2_X1 U547 ( .A1(n587), .A2(n588), .ZN(n589) );
  NOR2_X1 U548 ( .A1(n410), .A2(n720), .ZN(G63) );
  NAND2_X1 U549 ( .A1(n452), .A2(n446), .ZN(n451) );
  XNOR2_X2 U550 ( .A(n415), .B(n622), .ZN(n727) );
  NAND2_X1 U551 ( .A1(n620), .A2(n621), .ZN(n415) );
  XNOR2_X1 U552 ( .A(n453), .B(n634), .ZN(n452) );
  XNOR2_X1 U553 ( .A(n591), .B(n416), .ZN(n594) );
  NAND2_X1 U554 ( .A1(KEYINPUT2), .A2(n698), .ZN(n703) );
  NAND2_X1 U555 ( .A1(n420), .A2(n418), .ZN(n417) );
  AND2_X1 U556 ( .A1(n565), .A2(n421), .ZN(n420) );
  AND2_X1 U557 ( .A1(n457), .A2(n566), .ZN(n421) );
  INV_X1 U558 ( .A(n547), .ZN(n580) );
  INV_X1 U559 ( .A(n659), .ZN(n572) );
  XNOR2_X1 U560 ( .A(n434), .B(n433), .ZN(G51) );
  NOR2_X2 U561 ( .A1(n727), .A2(n735), .ZN(n698) );
  XNOR2_X2 U562 ( .A(n595), .B(KEYINPUT104), .ZN(n749) );
  AND2_X2 U563 ( .A1(n704), .A2(n703), .ZN(n713) );
  INV_X1 U564 ( .A(n727), .ZN(n450) );
  NAND2_X1 U565 ( .A1(n450), .A2(n449), .ZN(n448) );
  XNOR2_X1 U566 ( .A(n451), .B(KEYINPUT123), .ZN(G54) );
  NAND2_X1 U567 ( .A1(n713), .A2(G469), .ZN(n453) );
  XNOR2_X2 U568 ( .A(n522), .B(n462), .ZN(n465) );
  BUF_X1 U569 ( .A(n713), .Z(n716) );
  XNOR2_X2 U570 ( .A(G116), .B(KEYINPUT3), .ZN(n463) );
  AND2_X1 U571 ( .A1(G214), .A2(n534), .ZN(n455) );
  XOR2_X1 U572 ( .A(n493), .B(n492), .Z(n456) );
  OR2_X1 U573 ( .A1(KEYINPUT47), .A2(n564), .ZN(n457) );
  XNOR2_X1 U574 ( .A(n467), .B(n466), .ZN(n470) );
  NOR2_X1 U575 ( .A1(n553), .A2(n365), .ZN(n554) );
  XNOR2_X1 U576 ( .A(n490), .B(n489), .ZN(n717) );
  NOR2_X1 U577 ( .A1(n607), .A2(n592), .ZN(n593) );
  OR2_X1 U578 ( .A1(G237), .A2(G902), .ZN(n515) );
  NAND2_X1 U579 ( .A1(n515), .A2(G210), .ZN(n464) );
  NAND2_X1 U580 ( .A1(G224), .A2(n736), .ZN(n458) );
  XNOR2_X1 U581 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X2 U582 ( .A(n461), .B(G143), .ZN(n522) );
  XOR2_X1 U583 ( .A(G113), .B(G104), .Z(n535) );
  XNOR2_X1 U584 ( .A(G902), .B(KEYINPUT15), .ZN(n623) );
  XNOR2_X1 U585 ( .A(G137), .B(G140), .ZN(n485) );
  NAND2_X1 U586 ( .A1(G227), .A2(n736), .ZN(n467) );
  XOR2_X1 U587 ( .A(n468), .B(G107), .Z(n469) );
  XOR2_X1 U588 ( .A(KEYINPUT70), .B(G469), .Z(n472) );
  XNOR2_X2 U589 ( .A(n473), .B(n472), .ZN(n558) );
  XOR2_X1 U590 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n475) );
  NAND2_X1 U591 ( .A1(G234), .A2(n623), .ZN(n474) );
  XNOR2_X1 U592 ( .A(n475), .B(n474), .ZN(n491) );
  NAND2_X1 U593 ( .A1(n491), .A2(G221), .ZN(n476) );
  XNOR2_X1 U594 ( .A(n476), .B(KEYINPUT21), .ZN(n477) );
  XOR2_X1 U595 ( .A(KEYINPUT95), .B(n477), .Z(n671) );
  XNOR2_X1 U596 ( .A(G119), .B(KEYINPUT89), .ZN(n478) );
  XNOR2_X1 U597 ( .A(n479), .B(n478), .ZN(n482) );
  XOR2_X1 U598 ( .A(n482), .B(n481), .Z(n490) );
  NAND2_X1 U599 ( .A1(G234), .A2(n736), .ZN(n483) );
  XNOR2_X1 U600 ( .A(n484), .B(n483), .ZN(n527) );
  NAND2_X1 U601 ( .A1(n527), .A2(G221), .ZN(n488) );
  XNOR2_X1 U602 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U603 ( .A(n488), .B(n487), .ZN(n489) );
  NOR2_X1 U604 ( .A1(G902), .A2(n717), .ZN(n496) );
  NAND2_X1 U605 ( .A1(G217), .A2(n491), .ZN(n494) );
  XOR2_X1 U606 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n493) );
  XNOR2_X1 U607 ( .A(KEYINPUT71), .B(KEYINPUT25), .ZN(n492) );
  AND2_X1 U608 ( .A1(n558), .A2(n677), .ZN(n613) );
  NAND2_X1 U609 ( .A1(G234), .A2(G237), .ZN(n497) );
  XNOR2_X1 U610 ( .A(n497), .B(KEYINPUT86), .ZN(n498) );
  XNOR2_X1 U611 ( .A(KEYINPUT14), .B(n498), .ZN(n500) );
  NAND2_X1 U612 ( .A1(G952), .A2(n500), .ZN(n692) );
  NOR2_X1 U613 ( .A1(G953), .A2(n692), .ZN(n499) );
  XNOR2_X1 U614 ( .A(KEYINPUT87), .B(n499), .ZN(n585) );
  INV_X1 U615 ( .A(n585), .ZN(n505) );
  NAND2_X1 U616 ( .A1(n500), .A2(G902), .ZN(n501) );
  XOR2_X1 U617 ( .A(KEYINPUT88), .B(n501), .Z(n584) );
  NAND2_X1 U618 ( .A1(n584), .A2(n502), .ZN(n503) );
  NOR2_X1 U619 ( .A1(G900), .A2(n503), .ZN(n504) );
  NOR2_X1 U620 ( .A1(n505), .A2(n504), .ZN(n543) );
  NAND2_X1 U621 ( .A1(n534), .A2(G210), .ZN(n506) );
  XNOR2_X1 U622 ( .A(n507), .B(n506), .ZN(n513) );
  INV_X1 U623 ( .A(n508), .ZN(n509) );
  XNOR2_X1 U624 ( .A(n509), .B(G146), .ZN(n512) );
  XNOR2_X1 U625 ( .A(n510), .B(G137), .ZN(n511) );
  NAND2_X1 U626 ( .A1(G214), .A2(n515), .ZN(n658) );
  NAND2_X1 U627 ( .A1(n592), .A2(n658), .ZN(n516) );
  XNOR2_X1 U628 ( .A(KEYINPUT30), .B(n516), .ZN(n517) );
  NOR2_X1 U629 ( .A1(n543), .A2(n517), .ZN(n518) );
  NAND2_X1 U630 ( .A1(n613), .A2(n518), .ZN(n540) );
  XNOR2_X1 U631 ( .A(KEYINPUT101), .B(G478), .ZN(n531) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n520) );
  XNOR2_X1 U633 ( .A(KEYINPUT7), .B(KEYINPUT100), .ZN(n519) );
  XNOR2_X1 U634 ( .A(n520), .B(n519), .ZN(n526) );
  XOR2_X1 U635 ( .A(n521), .B(G116), .Z(n524) );
  XNOR2_X1 U636 ( .A(n522), .B(G134), .ZN(n523) );
  XNOR2_X1 U637 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U638 ( .A(n526), .B(n525), .Z(n529) );
  NAND2_X1 U639 ( .A1(G217), .A2(n527), .ZN(n528) );
  XNOR2_X1 U640 ( .A(n529), .B(n528), .ZN(n712) );
  NOR2_X1 U641 ( .A1(G902), .A2(n712), .ZN(n530) );
  XNOR2_X1 U642 ( .A(KEYINPUT13), .B(G475), .ZN(n539) );
  XOR2_X1 U643 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n533) );
  NOR2_X1 U644 ( .A1(G902), .A2(n707), .ZN(n538) );
  AND2_X1 U645 ( .A1(n571), .A2(n542), .ZN(n651) );
  AND2_X1 U646 ( .A1(n567), .A2(n651), .ZN(n654) );
  NAND2_X1 U647 ( .A1(n571), .A2(n570), .ZN(n603) );
  OR2_X1 U648 ( .A1(n580), .A2(n540), .ZN(n541) );
  NOR2_X1 U649 ( .A1(n603), .A2(n541), .ZN(n645) );
  NOR2_X1 U650 ( .A1(n568), .A2(n651), .ZN(n664) );
  INV_X1 U651 ( .A(n664), .ZN(n561) );
  OR2_X1 U652 ( .A1(KEYINPUT75), .A2(n561), .ZN(n548) );
  NOR2_X1 U653 ( .A1(n671), .A2(n543), .ZN(n544) );
  NAND2_X1 U654 ( .A1(n672), .A2(n544), .ZN(n553) );
  NOR2_X1 U655 ( .A1(n553), .A2(n611), .ZN(n545) );
  XNOR2_X1 U656 ( .A(n545), .B(KEYINPUT28), .ZN(n546) );
  AND2_X1 U657 ( .A1(n546), .A2(n558), .ZN(n574) );
  NAND2_X1 U658 ( .A1(n574), .A2(n587), .ZN(n562) );
  INV_X1 U659 ( .A(n562), .ZN(n646) );
  NAND2_X1 U660 ( .A1(n548), .A2(n646), .ZN(n549) );
  NAND2_X1 U661 ( .A1(n549), .A2(KEYINPUT47), .ZN(n551) );
  NAND2_X1 U662 ( .A1(n561), .A2(KEYINPUT75), .ZN(n550) );
  NAND2_X1 U663 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U664 ( .A1(n645), .A2(n552), .ZN(n566) );
  XNOR2_X1 U665 ( .A(KEYINPUT36), .B(KEYINPUT82), .ZN(n555) );
  XNOR2_X1 U666 ( .A(n556), .B(n555), .ZN(n559) );
  XNOR2_X2 U667 ( .A(n558), .B(n557), .ZN(n608) );
  XOR2_X1 U668 ( .A(n391), .B(KEYINPUT83), .Z(n596) );
  NAND2_X1 U669 ( .A1(n559), .A2(n596), .ZN(n560) );
  XNOR2_X1 U670 ( .A(n744), .B(KEYINPUT78), .ZN(n565) );
  XOR2_X1 U671 ( .A(n561), .B(KEYINPUT76), .Z(n616) );
  NOR2_X1 U672 ( .A1(n616), .A2(n562), .ZN(n563) );
  NOR2_X1 U673 ( .A1(KEYINPUT75), .A2(n563), .ZN(n564) );
  NAND2_X1 U674 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U675 ( .A1(n571), .A2(n570), .ZN(n590) );
  INV_X1 U676 ( .A(n590), .ZN(n661) );
  NOR2_X1 U677 ( .A1(n661), .A2(n663), .ZN(n573) );
  XOR2_X1 U678 ( .A(KEYINPUT42), .B(n575), .Z(n747) );
  NOR2_X1 U679 ( .A1(n393), .A2(n577), .ZN(n578) );
  NAND2_X1 U680 ( .A1(n578), .A2(n658), .ZN(n579) );
  XNOR2_X1 U681 ( .A(n579), .B(KEYINPUT43), .ZN(n581) );
  NAND2_X1 U682 ( .A1(n581), .A2(n580), .ZN(n656) );
  NAND2_X1 U683 ( .A1(n582), .A2(n656), .ZN(n735) );
  NOR2_X1 U684 ( .A1(G898), .A2(n583), .ZN(n723) );
  NAND2_X1 U685 ( .A1(n584), .A2(n723), .ZN(n586) );
  NAND2_X1 U686 ( .A1(n586), .A2(n585), .ZN(n588) );
  INV_X1 U687 ( .A(n672), .ZN(n607) );
  AND2_X1 U688 ( .A1(n672), .A2(n596), .ZN(n597) );
  NAND2_X1 U689 ( .A1(n609), .A2(n597), .ZN(n598) );
  XNOR2_X1 U690 ( .A(KEYINPUT32), .B(n598), .ZN(n746) );
  XNOR2_X1 U691 ( .A(n606), .B(KEYINPUT81), .ZN(n605) );
  INV_X1 U692 ( .A(KEYINPUT105), .ZN(n599) );
  NAND2_X1 U693 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n684) );
  NAND2_X1 U695 ( .A1(n600), .A2(n684), .ZN(n612) );
  XNOR2_X1 U696 ( .A(n612), .B(KEYINPUT31), .ZN(n652) );
  NAND2_X1 U697 ( .A1(n613), .A2(n600), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n652), .A2(n638), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n743), .A2(KEYINPUT44), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT80), .ZN(n618) );
  XNOR2_X1 U701 ( .A(KEYINPUT77), .B(KEYINPUT45), .ZN(n622) );
  INV_X1 U702 ( .A(n623), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n624), .A2(KEYINPUT2), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n629) );
  XNOR2_X1 U705 ( .A(n627), .B(KEYINPUT74), .ZN(n628) );
  XNOR2_X1 U706 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT57), .ZN(n632) );
  XOR2_X1 U708 ( .A(G101), .B(n636), .Z(G3) );
  NAND2_X1 U709 ( .A1(n649), .A2(n638), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n637), .B(G104), .ZN(G6) );
  XOR2_X1 U711 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n640) );
  NAND2_X1 U712 ( .A1(n638), .A2(n651), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U714 ( .A(G107), .B(n641), .ZN(G9) );
  XOR2_X1 U715 ( .A(KEYINPUT29), .B(KEYINPUT109), .Z(n643) );
  NAND2_X1 U716 ( .A1(n646), .A2(n651), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(n644) );
  XOR2_X1 U718 ( .A(G128), .B(n644), .Z(G30) );
  XOR2_X1 U719 ( .A(G143), .B(n645), .Z(G45) );
  NAND2_X1 U720 ( .A1(n649), .A2(n646), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT110), .ZN(n648) );
  XNOR2_X1 U722 ( .A(G146), .B(n648), .ZN(G48) );
  NAND2_X1 U723 ( .A1(n649), .A2(n652), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n650), .B(G113), .ZN(G15) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(G116), .ZN(G18) );
  XNOR2_X1 U727 ( .A(G134), .B(n654), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(KEYINPUT111), .ZN(G36) );
  XNOR2_X1 U729 ( .A(G140), .B(KEYINPUT112), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(G42) );
  NOR2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U733 ( .A(KEYINPUT117), .B(n662), .Z(n667) );
  NOR2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U735 ( .A(KEYINPUT118), .B(n665), .ZN(n666) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n669) );
  BUF_X1 U737 ( .A(n668), .Z(n694) );
  NOR2_X1 U738 ( .A1(n669), .A2(n694), .ZN(n670) );
  XNOR2_X1 U739 ( .A(KEYINPUT119), .B(n670), .ZN(n688) );
  XOR2_X1 U740 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n674) );
  NAND2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n592), .A2(n675), .ZN(n676) );
  XOR2_X1 U744 ( .A(KEYINPUT114), .B(n676), .Z(n682) );
  XOR2_X1 U745 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n679) );
  OR2_X1 U746 ( .A1(n677), .A2(n391), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n680) );
  XOR2_X1 U748 ( .A(KEYINPUT115), .B(n680), .Z(n681) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(KEYINPUT51), .B(n685), .ZN(n686) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U753 ( .A(n689), .B(KEYINPUT120), .ZN(n690) );
  XOR2_X1 U754 ( .A(KEYINPUT52), .B(n690), .Z(n691) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U756 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U758 ( .A(KEYINPUT121), .B(n697), .Z(n700) );
  XNOR2_X1 U759 ( .A(n698), .B(KEYINPUT2), .ZN(n699) );
  NAND2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U761 ( .A1(n701), .A2(G953), .ZN(n702) );
  XNOR2_X1 U762 ( .A(n702), .B(KEYINPUT53), .ZN(G75) );
  AND2_X1 U763 ( .A1(n703), .A2(G475), .ZN(n705) );
  NAND2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n709) );
  XOR2_X1 U765 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n706) );
  XNOR2_X1 U766 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U768 ( .A(n712), .B(KEYINPUT125), .Z(n715) );
  NAND2_X1 U769 ( .A1(n716), .A2(G478), .ZN(n714) );
  NAND2_X1 U770 ( .A1(n716), .A2(G217), .ZN(n719) );
  XOR2_X1 U771 ( .A(n721), .B(G101), .Z(n722) );
  XNOR2_X1 U772 ( .A(G110), .B(n722), .ZN(n724) );
  NOR2_X1 U773 ( .A1(n724), .A2(n723), .ZN(n731) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n725) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n725), .ZN(n726) );
  AND2_X1 U776 ( .A1(n726), .A2(G898), .ZN(n729) );
  NOR2_X1 U777 ( .A1(G953), .A2(n727), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U779 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(KEYINPUT127), .B(n732), .ZN(G69) );
  XOR2_X1 U781 ( .A(n734), .B(n733), .Z(n738) );
  XNOR2_X1 U782 ( .A(n735), .B(n738), .ZN(n737) );
  NAND2_X1 U783 ( .A1(n737), .A2(n736), .ZN(n742) );
  XNOR2_X1 U784 ( .A(G227), .B(n738), .ZN(n739) );
  NAND2_X1 U785 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n740), .A2(G953), .ZN(n741) );
  NAND2_X1 U787 ( .A1(n742), .A2(n741), .ZN(G72) );
  XOR2_X1 U788 ( .A(n743), .B(G122), .Z(G24) );
  XOR2_X1 U789 ( .A(n744), .B(G125), .Z(n745) );
  XNOR2_X1 U790 ( .A(KEYINPUT37), .B(n745), .ZN(G27) );
  XNOR2_X1 U791 ( .A(G119), .B(n746), .ZN(G21) );
  XOR2_X1 U792 ( .A(G137), .B(n747), .Z(G39) );
  XOR2_X1 U793 ( .A(G131), .B(n748), .Z(G33) );
  XNOR2_X1 U794 ( .A(n749), .B(G110), .ZN(G12) );
endmodule

