//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G169gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G197gat), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n204), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G197gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n206), .A2(new_n210), .A3(KEYINPUT12), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT12), .B1(new_n206), .B2(new_n210), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n214));
  OR2_X1    g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT14), .ZN(new_n216));
  XOR2_X1   g015(.A(G43gat), .B(G50gat), .Z(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G29gat), .A2(G36gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n217), .A2(new_n218), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n221), .A2(new_n222), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n214), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n225), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT17), .A3(new_n223), .ZN(new_n228));
  XNOR2_X1  g027(.A(G15gat), .B(G22gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(G1gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G1gat), .B2(new_n229), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(G8gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n226), .A2(new_n228), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n224), .B2(new_n225), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT18), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n224), .A2(new_n225), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n236), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n237), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n235), .A2(new_n237), .A3(new_n236), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n239), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n213), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n249), .A2(new_n213), .A3(new_n246), .A4(new_n241), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n255));
  OR2_X1    g054(.A1(G113gat), .A2(G120gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n257));
  NAND2_X1  g056(.A1(G113gat), .A2(G120gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G134gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G127gat), .ZN(new_n261));
  INV_X1    g060(.A(G127gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G134gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n255), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(G113gat), .A2(G120gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(G113gat), .A2(G120gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT70), .A4(new_n257), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n272), .A3(new_n258), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n266), .B2(new_n267), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n257), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n276), .A2(new_n262), .A3(G134gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n277), .B1(new_n276), .B2(new_n269), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n271), .A2(new_n279), .A3(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT24), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(G183gat), .A3(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n207), .A2(new_n294), .A3(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(KEYINPUT64), .ZN(new_n302));
  OR3_X1    g101(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n289), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AND4_X1   g103(.A1(KEYINPUT25), .A2(new_n295), .A3(new_n297), .A4(new_n298), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n300), .A2(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n290), .A2(KEYINPUT27), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n291), .B1(new_n308), .B2(KEYINPUT65), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT27), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G183gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n290), .A2(KEYINPUT27), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n307), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n307), .A2(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT26), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT66), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n327), .A2(new_n298), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n326), .A2(new_n328), .B1(G183gat), .B2(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n306), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n319), .A2(new_n329), .A3(KEYINPUT67), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n284), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n316), .A2(new_n317), .ZN(new_n335));
  AOI21_X1  g134(.A(G190gat), .B1(new_n312), .B2(new_n310), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n310), .B2(new_n316), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n337), .B2(new_n307), .ZN(new_n338));
  INV_X1    g137(.A(new_n325), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n324), .B1(new_n320), .B2(new_n321), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n328), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n285), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n331), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n300), .A2(new_n301), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n305), .A2(new_n304), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n333), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n271), .A2(new_n279), .A3(KEYINPUT71), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT71), .B1(new_n271), .B2(new_n279), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G227gat), .ZN(new_n352));
  INV_X1    g151(.A(G233gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT32), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n359));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n355), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n358), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n355), .B(KEYINPUT32), .C1(new_n363), .C2(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT34), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n347), .B(new_n284), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(new_n354), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n334), .A2(new_n351), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n371), .B(KEYINPUT34), .C1(new_n352), .C2(new_n353), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT73), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n365), .A2(new_n373), .A3(new_n366), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n377), .A2(KEYINPUT36), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n365), .B2(new_n366), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT36), .B1(new_n375), .B2(new_n377), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  INV_X1    g187(.A(G148gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G141gat), .ZN(new_n390));
  INV_X1    g189(.A(G141gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G148gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n390), .A2(new_n392), .B1(KEYINPUT2), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G155gat), .ZN(new_n395));
  INV_X1    g194(.A(G162gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT77), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(G155gat), .B2(G162gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n393), .A2(KEYINPUT76), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(G155gat), .A3(G162gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n394), .B1(new_n405), .B2(KEYINPUT78), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n399), .A2(new_n397), .B1(new_n401), .B2(new_n403), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n389), .A2(KEYINPUT80), .A3(G141gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(G141gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n411), .B(new_n412), .C1(new_n414), .C2(new_n389), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n393), .A2(KEYINPUT2), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(KEYINPUT81), .ZN(new_n417));
  INV_X1    g216(.A(new_n393), .ZN(new_n418));
  NOR2_X1   g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT81), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n393), .B2(KEYINPUT2), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n417), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n406), .A2(new_n409), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n350), .A2(new_n387), .A3(new_n388), .A4(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n282), .A2(new_n388), .A3(new_n424), .A4(new_n283), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT82), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n409), .ZN(new_n428));
  INV_X1    g227(.A(new_n417), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n420), .A2(new_n422), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n413), .A2(G148gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n412), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n429), .B(new_n430), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n428), .A2(new_n433), .A3(new_n279), .A4(new_n271), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT4), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n425), .A2(new_n427), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(KEYINPUT5), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n428), .A2(new_n440), .A3(new_n433), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n280), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n424), .A2(new_n440), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n439), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n394), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n407), .B2(new_n408), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n405), .A2(KEYINPUT78), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n433), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT3), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(new_n280), .A3(new_n441), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n434), .B1(new_n388), .B2(new_n438), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n282), .A2(KEYINPUT4), .A3(new_n424), .A4(new_n283), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n449), .A2(new_n280), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n434), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n457), .B2(new_n438), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n436), .A2(new_n445), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT0), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(G57gat), .ZN(new_n462));
  INV_X1    g261(.A(G85gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n386), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT6), .B1(new_n459), .B2(new_n464), .ZN(new_n466));
  INV_X1    g265(.A(new_n464), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n454), .A2(new_n458), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n426), .A2(KEYINPUT82), .B1(KEYINPUT4), .B2(new_n434), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n444), .B1(new_n469), .B2(new_n425), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT83), .B(new_n467), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT6), .B(new_n467), .C1(new_n468), .C2(new_n470), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(KEYINPUT29), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n347), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n330), .A2(new_n346), .A3(new_n475), .ZN(new_n478));
  XNOR2_X1  g277(.A(G197gat), .B(G204gat), .ZN(new_n479));
  INV_X1    g278(.A(G211gat), .ZN(new_n480));
  INV_X1    g279(.A(G218gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(KEYINPUT22), .B2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(G211gat), .B(G218gat), .Z(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n477), .A2(new_n478), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n343), .A2(new_n333), .A3(new_n475), .A4(new_n346), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n338), .A2(new_n342), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n476), .B1(new_n489), .B2(new_n306), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n485), .ZN(new_n492));
  XNOR2_X1  g291(.A(G64gat), .B(G92gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G36gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT74), .B(G8gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n487), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT75), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT30), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n487), .A2(new_n492), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n501), .A2(new_n496), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n497), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n474), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n485), .B1(new_n441), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT3), .B1(new_n485), .B2(new_n508), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(new_n424), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT84), .B1(new_n510), .B2(new_n424), .ZN(new_n513));
  AND2_X1   g312(.A1(G228gat), .A2(G233gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n513), .B(new_n514), .C1(new_n509), .C2(new_n511), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G22gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n517), .A3(G22gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT31), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(G50gat), .Z(new_n525));
  AOI21_X1  g324(.A(G22gat), .B1(new_n516), .B2(new_n517), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(KEYINPUT85), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n520), .A2(KEYINPUT85), .A3(new_n521), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n507), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT86), .B1(new_n459), .B2(new_n464), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(new_n467), .C1(new_n468), .C2(new_n470), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n466), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT37), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n487), .A2(new_n492), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n477), .A2(new_n478), .A3(new_n485), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n491), .A2(new_n486), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT37), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT38), .ZN(new_n541));
  INV_X1    g340(.A(new_n496), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n537), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n473), .A2(new_n543), .A3(new_n497), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n535), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n535), .B2(new_n544), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n501), .A2(new_n536), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n537), .A2(new_n542), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n532), .A2(new_n534), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT40), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n437), .B1(new_n436), .B2(new_n451), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n456), .A2(new_n434), .A3(new_n437), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT39), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n464), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n451), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n469), .B2(new_n425), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n559), .A2(KEYINPUT39), .A3(new_n437), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n553), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT39), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT39), .B(new_n555), .C1(new_n559), .C2(new_n437), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT40), .A4(new_n464), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n552), .A2(new_n561), .A3(new_n565), .A4(new_n505), .ZN(new_n566));
  INV_X1    g365(.A(new_n530), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n385), .B(new_n531), .C1(new_n551), .C2(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n375), .A2(new_n377), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n535), .A2(new_n473), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n570), .A2(new_n567), .A3(new_n506), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT35), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n379), .A2(new_n380), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n528), .A2(new_n377), .A3(new_n529), .ZN(new_n575));
  AOI211_X1 g374(.A(KEYINPUT73), .B(new_n373), .C1(new_n365), .C2(new_n366), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI211_X1 g376(.A(new_n573), .B(new_n505), .C1(new_n473), .C2(new_n472), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n572), .A2(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n254), .B1(new_n569), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G57gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G64gat), .ZN(new_n582));
  INV_X1    g381(.A(G64gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G57gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT90), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n582), .B2(new_n584), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n586), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n585), .A2(new_n588), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n596));
  INV_X1    g395(.A(new_n586), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT89), .B1(new_n591), .B2(new_n586), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT92), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n233), .B1(KEYINPUT21), .B2(new_n601), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT93), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT20), .ZN(new_n610));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT94), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n608), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n242), .ZN(new_n617));
  NAND2_X1  g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(KEYINPUT95), .A2(G99gat), .A3(G106gat), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(KEYINPUT8), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT7), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n625), .A2(new_n463), .A3(G92gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n622), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G99gat), .B(G106gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n630), .B(new_n622), .C1(new_n624), .C2(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n617), .A2(new_n633), .B1(KEYINPUT41), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n226), .A2(new_n228), .A3(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n637), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n634), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(G190gat), .B(G218gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n640), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n591), .A2(KEYINPUT89), .A3(new_n586), .ZN(new_n647));
  AND4_X1   g446(.A1(new_n592), .A2(new_n585), .A3(new_n586), .A4(new_n588), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n592), .B1(new_n591), .B2(new_n586), .ZN(new_n649));
  OAI22_X1  g448(.A1(new_n646), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n632), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n594), .A2(new_n600), .A3(new_n629), .A4(new_n631), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(KEYINPUT96), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n601), .A2(new_n633), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT97), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n652), .A2(KEYINPUT10), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n653), .A2(new_n659), .A3(new_n656), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  INV_X1    g464(.A(G204gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT98), .B(G176gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n664), .A2(new_n669), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n580), .A2(new_n616), .A3(new_n645), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT99), .ZN(new_n675));
  INV_X1    g474(.A(new_n474), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT100), .B(G1gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1324gat));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  NAND3_X1  g479(.A1(new_n675), .A2(new_n505), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n675), .A2(new_n505), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n681), .A2(new_n682), .B1(new_n683), .B2(G8gat), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n685), .A2(KEYINPUT101), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(KEYINPUT101), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(G1325gat));
  INV_X1    g487(.A(G15gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n675), .A2(new_n689), .A3(new_n570), .ZN(new_n690));
  INV_X1    g489(.A(new_n385), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n675), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n692), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g492(.A1(new_n675), .A2(new_n530), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT102), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n694), .B(new_n696), .ZN(G1327gat));
  INV_X1    g496(.A(new_n616), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n673), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n645), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n580), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(G29gat), .A3(new_n474), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n699), .A2(new_n254), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n569), .A2(new_n579), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n644), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT44), .B(new_n645), .C1(new_n569), .C2(new_n579), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710), .B2(new_n474), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n704), .A2(new_n711), .ZN(G1328gat));
  OAI21_X1  g511(.A(G36gat), .B1(new_n710), .B2(new_n506), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n701), .A2(G36gat), .A3(new_n506), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n716), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT105), .B1(new_n716), .B2(KEYINPUT46), .ZN(new_n718));
  OAI221_X1 g517(.A(new_n713), .B1(KEYINPUT46), .B2(new_n716), .C1(new_n717), .C2(new_n718), .ZN(G1329gat));
  NAND2_X1  g518(.A1(new_n375), .A2(new_n377), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n701), .A2(G43gat), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT107), .ZN(new_n722));
  OAI21_X1  g521(.A(G43gat), .B1(new_n710), .B2(new_n385), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT106), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g524(.A(G50gat), .B1(new_n710), .B2(new_n567), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n567), .A2(G50gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n701), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g528(.A1(new_n616), .A2(new_n645), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n253), .A3(new_n673), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n707), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n676), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT108), .B(G57gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1332gat));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n505), .B1(new_n736), .B2(new_n583), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT109), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n583), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  NAND2_X1  g540(.A1(new_n732), .A2(new_n691), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n720), .A2(G71gat), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n742), .A2(G71gat), .B1(new_n732), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n732), .A2(new_n530), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g546(.A1(new_n616), .A2(new_n253), .A3(new_n673), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n708), .B2(new_n709), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT110), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n748), .C1(new_n708), .C2(new_n709), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n676), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G85gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n616), .A2(new_n253), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n547), .A2(new_n550), .ZN(new_n756));
  INV_X1    g555(.A(new_n546), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n568), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n377), .A2(KEYINPUT36), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n574), .A2(new_n576), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n531), .B1(new_n760), .B2(new_n383), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n572), .A2(new_n573), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n577), .A2(new_n578), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n644), .B(new_n755), .C1(new_n762), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT51), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n707), .A2(new_n768), .A3(new_n644), .A4(new_n755), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n767), .A2(new_n672), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n463), .A3(new_n676), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT111), .ZN(G1336gat));
  OAI21_X1  g572(.A(G92gat), .B1(new_n749), .B2(new_n506), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n506), .A2(G92gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n767), .A2(new_n672), .A3(new_n769), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n750), .A2(new_n505), .A3(new_n752), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n777), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n779), .B1(new_n784), .B2(KEYINPUT52), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT113), .B(new_n775), .C1(new_n781), .C2(new_n783), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n778), .B1(new_n785), .B2(new_n786), .ZN(G1337gat));
  AOI21_X1  g586(.A(G99gat), .B1(new_n770), .B2(new_n570), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n750), .A2(new_n752), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n691), .A2(G99gat), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(G1338gat));
  NOR2_X1   g590(.A1(new_n567), .A2(G106gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n770), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  OAI21_X1  g593(.A(G106gat), .B1(new_n749), .B2(new_n567), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT114), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n789), .A2(new_n530), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n798), .A2(G106gat), .B1(new_n770), .B2(new_n792), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n794), .B2(new_n799), .ZN(G1339gat));
  NOR3_X1   g599(.A1(new_n730), .A2(new_n253), .A3(new_n672), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n662), .A2(KEYINPUT54), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n669), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n657), .A2(new_n661), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n659), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(KEYINPUT54), .A3(new_n662), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n805), .B2(new_n659), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n808), .A2(KEYINPUT116), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811));
  AOI211_X1 g610(.A(KEYINPUT115), .B(new_n660), .C1(new_n657), .C2(new_n661), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n662), .A2(KEYINPUT54), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n809), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n804), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(KEYINPUT117), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT116), .B1(new_n808), .B2(new_n809), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n814), .A2(new_n811), .A3(new_n815), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n803), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n823), .B2(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n822), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n803), .A2(new_n818), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n206), .A2(new_n210), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n244), .A2(new_n245), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n237), .B1(new_n235), .B2(new_n236), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n252), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n835), .A2(new_n644), .A3(new_n670), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n825), .A2(new_n828), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n673), .A2(new_n833), .ZN(new_n838));
  INV_X1    g637(.A(new_n252), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n670), .B1(new_n250), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n826), .B2(new_n827), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n838), .B1(new_n825), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n837), .B1(new_n842), .B2(new_n644), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n801), .B1(new_n843), .B2(new_n698), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n474), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n577), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(KEYINPUT119), .A3(new_n577), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n505), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n253), .ZN(new_n851));
  INV_X1    g650(.A(new_n844), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n676), .A2(new_n506), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n530), .A3(new_n720), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n253), .A2(G113gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(G1340gat));
  AOI21_X1  g656(.A(G120gat), .B1(new_n850), .B2(new_n672), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(G120gat), .A3(new_n672), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n505), .B(new_n673), .C1(new_n848), .C2(new_n849), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n862), .B(new_n859), .C1(new_n863), .C2(G120gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(G1341gat));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n262), .A3(new_n616), .ZN(new_n866));
  INV_X1    g665(.A(new_n855), .ZN(new_n867));
  OAI21_X1  g666(.A(G127gat), .B1(new_n867), .B2(new_n698), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(G1342gat));
  NAND2_X1  g668(.A1(new_n848), .A2(new_n849), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n644), .A2(new_n506), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT121), .Z(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n260), .A3(new_n873), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n867), .B2(new_n645), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n567), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n838), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n828), .A2(new_n253), .A3(new_n670), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n823), .A2(KEYINPUT55), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n817), .A2(new_n818), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n838), .B1(new_n887), .B2(new_n841), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT122), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n886), .A2(new_n645), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n616), .B1(new_n890), .B2(new_n837), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n880), .B1(new_n891), .B2(new_n801), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n882), .B1(new_n824), .B2(new_n819), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n645), .B1(new_n894), .B2(new_n838), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n616), .B1(new_n895), .B2(new_n837), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n530), .B1(new_n896), .B2(new_n801), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n892), .A2(new_n893), .B1(new_n897), .B2(new_n879), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT123), .B(new_n880), .C1(new_n891), .C2(new_n801), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n691), .A2(new_n853), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n253), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n414), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n845), .A2(new_n530), .A3(new_n385), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(new_n505), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n391), .A3(new_n253), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n901), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n898), .B2(new_n899), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n413), .B1(new_n910), .B2(new_n253), .ZN(new_n911));
  INV_X1    g710(.A(new_n907), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT58), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n906), .A2(new_n389), .A3(new_n672), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n844), .B2(new_n567), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n645), .B1(new_n888), .B2(KEYINPUT122), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n885), .B(new_n838), .C1(new_n887), .C2(new_n841), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n837), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n616), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n890), .A2(KEYINPUT124), .A3(new_n837), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n801), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n530), .A2(new_n879), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n926), .A2(new_n673), .A3(new_n909), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n916), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT59), .B(new_n389), .C1(new_n910), .C2(new_n672), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n915), .B1(new_n928), .B2(new_n929), .ZN(G1345gat));
  AOI21_X1  g729(.A(new_n395), .B1(new_n910), .B2(new_n616), .ZN(new_n931));
  NOR4_X1   g730(.A1(new_n905), .A2(G155gat), .A3(new_n505), .A4(new_n698), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n931), .A2(new_n932), .ZN(G1346gat));
  AOI21_X1  g732(.A(new_n396), .B1(new_n910), .B2(new_n644), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n905), .A2(G162gat), .A3(new_n872), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(G1347gat));
  NOR3_X1   g735(.A1(new_n844), .A2(new_n676), .A3(new_n506), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n720), .A2(new_n530), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n207), .A3(new_n254), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n937), .A2(new_n577), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n253), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n940), .B1(new_n207), .B2(new_n943), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n939), .B2(new_n673), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n672), .A2(new_n294), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT125), .ZN(G1349gat));
  OAI21_X1  g747(.A(G183gat), .B1(new_n939), .B2(new_n698), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n616), .A2(new_n316), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n941), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n942), .A2(new_n291), .A3(new_n644), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n644), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n955), .A3(G190gat), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n955), .B1(new_n954), .B2(G190gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  OR2_X1    g758(.A1(new_n926), .A2(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n926), .A2(KEYINPUT126), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n676), .A2(new_n506), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n385), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(new_n209), .A3(new_n254), .ZN(new_n965));
  INV_X1    g764(.A(new_n897), .ZN(new_n966));
  INV_X1    g765(.A(new_n964), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n253), .A3(new_n967), .ZN(new_n968));
  AOI22_X1  g767(.A1(new_n962), .A2(new_n965), .B1(new_n209), .B2(new_n968), .ZN(G1352gat));
  NOR2_X1   g768(.A1(new_n964), .A2(new_n673), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n960), .A2(new_n961), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G204gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n966), .A2(new_n666), .A3(new_n970), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1353gat));
  NOR2_X1   g774(.A1(new_n964), .A2(new_n698), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n966), .A2(new_n480), .A3(new_n976), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n917), .B(new_n976), .C1(new_n924), .C2(new_n925), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n983), .B(new_n977), .C1(new_n979), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1354gat));
  NOR3_X1   g784(.A1(new_n964), .A2(new_n481), .A3(new_n645), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n966), .A2(new_n644), .A3(new_n967), .ZN(new_n987));
  AOI22_X1  g786(.A1(new_n962), .A2(new_n986), .B1(new_n481), .B2(new_n987), .ZN(G1355gat));
endmodule


