//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n458), .B1(new_n448), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n468), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n465), .A2(new_n472), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G124), .B1(G136), .B2(new_n471), .ZN(new_n477));
  INV_X1    g052(.A(G100), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n478), .A2(new_n472), .A3(KEYINPUT66), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT66), .B1(new_n478), .B2(new_n472), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G112), .B2(new_n472), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n469), .A2(new_n470), .ZN(new_n489));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(KEYINPUT68), .B(new_n490), .C1(new_n463), .C2(new_n464), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n472), .C1(new_n463), .C2(new_n464), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n489), .A2(new_n498), .A3(G138), .A4(new_n472), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n494), .A2(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n490), .B1(new_n463), .B2(new_n464), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI211_X1 g078(.A(new_n495), .B(new_n487), .C1(new_n503), .C2(new_n492), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT71), .Z(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n512), .A2(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(KEYINPUT70), .A3(G50), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT5), .B(G543), .Z(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n517), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n521), .A2(new_n524), .B1(G88), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n512), .A2(KEYINPUT72), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n513), .A2(new_n527), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n523), .A2(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n518), .A2(new_n508), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G89), .Z(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n534), .A2(new_n538), .ZN(G168));
  NAND2_X1  g114(.A1(new_n523), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n532), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G651), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(new_n523), .A2(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n532), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n544), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n525), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n526), .B2(G91), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI211_X1 g138(.A(KEYINPUT74), .B(new_n562), .C1(new_n519), .C2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n565), .B2(KEYINPUT9), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n523), .B(new_n566), .C1(new_n565), .C2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n561), .A2(new_n564), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  NAND2_X1  g145(.A1(new_n526), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n523), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n525), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n523), .B2(G48), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(new_n532), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n526), .A2(new_n581), .A3(G86), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n544), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n523), .A2(G47), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT76), .B(G85), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n532), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n586), .B(new_n590), .C1(new_n532), .C2(new_n587), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n585), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n532), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n525), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(new_n523), .B2(G54), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G171), .ZN(G284));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G171), .ZN(G321));
  NAND2_X1  g182(.A1(G299), .A2(new_n604), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n604), .B2(G168), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(new_n604), .B2(G168), .ZN(G280));
  AND2_X1   g185(.A1(new_n598), .A2(new_n602), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n489), .A2(new_n473), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n471), .A2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n472), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n489), .A2(G2105), .ZN(new_n628));
  OAI221_X1 g203(.A(new_n624), .B1(new_n625), .B2(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n622), .A2(new_n623), .A3(new_n630), .ZN(G156));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n641), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n643), .B1(new_n642), .B2(new_n644), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n632), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g225(.A(KEYINPUT78), .B(new_n648), .C1(new_n645), .C2(new_n646), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G14), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n647), .B2(new_n649), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT79), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n656), .A2(new_n657), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n664), .B(new_n668), .Z(G227));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT81), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(KEYINPUT20), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n671), .A2(new_n672), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n680), .A3(new_n676), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n671), .A2(new_n672), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(new_n677), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n676), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n683), .ZN(new_n686));
  AOI21_X1  g261(.A(KEYINPUT82), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n686), .A3(KEYINPUT82), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(new_n689), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n687), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  INV_X1    g273(.A(new_n696), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n691), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  AND3_X1   g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n698), .B1(new_n697), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(G229));
  MUX2_X1   g278(.A(G6), .B(G305), .S(G16), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT84), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(G166), .A2(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G16), .B2(G22), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  INV_X1    g289(.A(G288), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT85), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  AND4_X1   g294(.A1(new_n707), .A2(new_n711), .A3(new_n712), .A4(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n471), .A2(G131), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n472), .A2(G107), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  INV_X1    g300(.A(G119), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n723), .B1(new_n724), .B2(new_n725), .C1(new_n726), .C2(new_n628), .ZN(new_n727));
  MUX2_X1   g302(.A(G25), .B(new_n727), .S(G29), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n713), .A2(G24), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT83), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n592), .B2(new_n713), .ZN(new_n733));
  INV_X1    g308(.A(G1986), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n722), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n720), .A2(new_n721), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT36), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G26), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT88), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n471), .A2(G140), .ZN(new_n747));
  INV_X1    g322(.A(G128), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n628), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n746), .A2(new_n749), .A3(KEYINPUT89), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT89), .B1(new_n746), .B2(new_n749), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n741), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n743), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(G162), .A2(G29), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G29), .B2(G35), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT29), .B(G2090), .Z(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR2_X1   g338(.A1(G4), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n611), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT86), .B(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n762), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G19), .ZN(new_n770));
  OR3_X1    g345(.A1(new_n770), .A2(KEYINPUT87), .A3(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(KEYINPUT87), .B1(new_n770), .B2(G16), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n771), .B(new_n772), .C1(new_n552), .C2(new_n713), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G1341), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT30), .B(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n775), .A2(new_n741), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n629), .B2(new_n741), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(new_n472), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n782));
  NAND2_X1  g357(.A1(G103), .A2(G2104), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G2105), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n471), .A2(G139), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n741), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n741), .B2(G33), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT92), .B(G2072), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n779), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n713), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT95), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT23), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT96), .B(G1956), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n774), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G171), .A2(new_n713), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G5), .B2(new_n713), .ZN(new_n801));
  INV_X1    g376(.A(G1961), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(G160), .A2(G29), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G34), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n804), .B1(G29), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G2084), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n803), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n790), .A2(new_n791), .B1(new_n801), .B2(new_n802), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n713), .A2(G21), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G168), .B2(new_n713), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1966), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n799), .A2(new_n811), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n741), .A2(G32), .ZN(new_n817));
  NAND3_X1  g392(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT94), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT26), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n471), .A2(G141), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n473), .A2(G105), .ZN(new_n823));
  INV_X1    g398(.A(G129), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n822), .B(new_n823), .C1(new_n824), .C2(new_n628), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n817), .B1(new_n826), .B2(new_n741), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT27), .ZN(new_n828));
  INV_X1    g403(.A(G1996), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n741), .A2(G27), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G164), .B2(new_n741), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G2078), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n758), .A2(new_n769), .A3(new_n816), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n739), .A2(new_n835), .ZN(G311));
  OR2_X1    g411(.A1(new_n739), .A2(new_n835), .ZN(G150));
  XNOR2_X1  g412(.A(KEYINPUT97), .B(G55), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n526), .A2(G93), .B1(new_n523), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n544), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT99), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n839), .B(new_n843), .C1(new_n544), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n611), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n842), .B(new_n844), .C1(new_n551), .C2(new_n549), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n552), .A2(new_n841), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n552), .A2(new_n841), .A3(KEYINPUT98), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n849), .B(new_n855), .Z(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  INV_X1    g433(.A(G860), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n857), .B2(KEYINPUT39), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n847), .B1(new_n858), .B2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n727), .B(new_n619), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n821), .A2(new_n825), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n787), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n788), .A2(new_n826), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n727), .B(new_n619), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n787), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n788), .A2(new_n826), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n750), .A2(new_n751), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n498), .B1(new_n471), .B2(G138), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT100), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n487), .B1(new_n503), .B2(new_n492), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n497), .A2(new_n499), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(new_n497), .B2(new_n499), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(new_n494), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n750), .A2(new_n751), .A3(new_n878), .A4(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  INV_X1    g459(.A(G118), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(G2105), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n476), .B2(G130), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n471), .A2(KEYINPUT101), .A3(G142), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT101), .B1(new_n471), .B2(G142), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n880), .A2(new_n883), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n880), .B2(new_n883), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n871), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n866), .A2(new_n870), .ZN(new_n895));
  INV_X1    g470(.A(new_n891), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G160), .B(new_n629), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n899), .A2(new_n483), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n483), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n900), .A2(new_n902), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n894), .A2(new_n897), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT102), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n894), .A2(new_n897), .A3(new_n912), .A4(new_n909), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n908), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(G395));
  NAND2_X1  g491(.A1(new_n845), .A2(new_n604), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n855), .B(new_n614), .Z(new_n919));
  INV_X1    g494(.A(G299), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n603), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT105), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n920), .A2(new_n603), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n920), .A2(new_n603), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n927), .A2(new_n928), .B1(new_n921), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n919), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n921), .ZN(new_n932));
  AOI211_X1 g507(.A(new_n918), .B(new_n931), .C1(new_n919), .C2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n918), .B2(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  XNOR2_X1  g510(.A(G305), .B(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(G303), .ZN(new_n937));
  NAND2_X1  g512(.A1(G290), .A2(KEYINPUT107), .ZN(new_n938));
  AOI211_X1 g513(.A(KEYINPUT107), .B(new_n585), .C1(new_n589), .C2(new_n591), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n940), .A3(new_n715), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n592), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(G288), .B1(new_n943), .B2(new_n939), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n937), .A2(KEYINPUT109), .A3(new_n941), .A4(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(KEYINPUT109), .A3(new_n944), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n936), .B(G166), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT109), .B1(new_n941), .B2(new_n944), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT42), .Z(new_n951));
  XNOR2_X1  g526(.A(new_n934), .B(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n917), .B1(new_n952), .B2(new_n604), .ZN(G295));
  OAI21_X1  g528(.A(new_n917), .B1(new_n952), .B2(new_n604), .ZN(G331));
  XNOR2_X1  g529(.A(G168), .B(G171), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n855), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n855), .A2(new_n956), .A3(KEYINPUT110), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n955), .A2(new_n850), .A3(new_n854), .A4(new_n853), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n932), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n957), .A2(new_n962), .ZN(new_n964));
  OAI22_X1  g539(.A1(new_n961), .A2(new_n963), .B1(new_n964), .B2(new_n930), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n907), .B1(new_n965), .B2(new_n950), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n964), .A2(new_n930), .ZN(new_n967));
  INV_X1    g542(.A(new_n963), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n959), .A3(new_n960), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n941), .A2(new_n944), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(new_n946), .A3(new_n947), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n967), .A2(new_n969), .B1(new_n973), .B2(new_n945), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n966), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n968), .A2(new_n957), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n855), .A2(new_n956), .A3(KEYINPUT110), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT110), .B1(new_n855), .B2(new_n956), .ZN(new_n978));
  INV_X1    g553(.A(new_n962), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n922), .A2(new_n926), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n981), .A2(new_n929), .B1(new_n928), .B2(new_n932), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n976), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n950), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n967), .A2(new_n973), .A3(new_n945), .A4(new_n969), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n907), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n975), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(KEYINPUT44), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n966), .B1(new_n950), .B2(new_n983), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n991));
  OR3_X1    g566(.A1(new_n990), .A2(new_n991), .A3(new_n986), .ZN(new_n992));
  OR3_X1    g567(.A1(new_n966), .A2(new_n974), .A3(KEYINPUT43), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n990), .B2(new_n986), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n989), .B1(new_n995), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n497), .A2(new_n499), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n876), .B2(KEYINPUT69), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n999), .B2(new_n504), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n879), .A2(new_n997), .A3(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1001), .A2(new_n808), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT45), .B1(new_n879), .B2(new_n997), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G1384), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n500), .B2(new_n505), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1007), .A2(new_n1011), .A3(new_n1002), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1006), .B1(new_n1012), .B2(G1966), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1013), .A2(G8), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1014), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n882), .B2(new_n878), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1003), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n715), .A2(G1976), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(G8), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT52), .ZN(new_n1020));
  INV_X1    g595(.A(G48), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n519), .A2(new_n1021), .B1(new_n1022), .B2(new_n544), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n532), .A2(new_n579), .ZN(new_n1024));
  OAI21_X1  g599(.A(G1981), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(G305), .B2(G1981), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1025), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(G8), .A3(new_n1017), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1017), .A2(G8), .A3(new_n1018), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1020), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1002), .B1(new_n879), .B2(new_n1009), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1384), .B1(new_n500), .B2(new_n505), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(KEYINPUT45), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n710), .ZN(new_n1042));
  INV_X1    g617(.A(G2090), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1001), .A2(new_n1043), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1038), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1034), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(KEYINPUT113), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1037), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1045), .B2(KEYINPUT113), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1015), .B(new_n1046), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1014), .A2(G168), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1045), .A2(new_n1037), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1020), .A2(new_n1033), .A3(new_n1030), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1055), .B(new_n997), .C1(new_n999), .C2(new_n504), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(new_n1003), .C1(new_n1016), .C2(new_n1004), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1042), .B1(G2090), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1037), .B1(new_n1058), .B2(G8), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1051), .A2(new_n1054), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1050), .B1(new_n1060), .B2(KEYINPUT63), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n879), .A2(new_n997), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n1002), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1030), .A2(new_n1031), .A3(new_n715), .ZN(new_n1064));
  OR2_X1    g639(.A1(G305), .A2(G1981), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1038), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1052), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(new_n1053), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1061), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1006), .B(G168), .C1(new_n1012), .C2(G1966), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1070), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(new_n1070), .B2(G8), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1014), .A2(G286), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT62), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1041), .B2(G2078), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n802), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1007), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1011), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1083), .A2(G2078), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1003), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1084), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1082), .B1(new_n1091), .B2(G171), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n1082), .A3(G171), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1058), .A2(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1048), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1046), .A2(KEYINPUT123), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1069), .B1(new_n1081), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1091), .A2(new_n1082), .A3(G171), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n1009), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT53), .B1(KEYINPUT122), .B2(G2078), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(KEYINPUT122), .B2(G2078), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1087), .A2(new_n1003), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1084), .A2(new_n1086), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(G171), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1107), .A2(new_n1092), .A3(new_n1113), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1114), .A2(KEYINPUT54), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(G171), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1116), .B(KEYINPUT54), .C1(G171), .C2(new_n1091), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1097), .A2(new_n1100), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1106), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1097), .A2(new_n1100), .A3(new_n1117), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1095), .B2(new_n1113), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(new_n1080), .A3(new_n1122), .A4(KEYINPUT124), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1039), .B(new_n1124), .C1(new_n1040), .C2(KEYINPUT45), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1956), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1057), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT114), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n920), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(KEYINPUT114), .A2(KEYINPUT57), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1134));
  NAND3_X1  g709(.A1(G299), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1000), .A2(new_n1008), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1138), .A2(KEYINPUT115), .A3(new_n1039), .A4(new_n1124), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1127), .A2(new_n1129), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1348), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1085), .A2(new_n1142), .B1(new_n757), .B2(new_n1063), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1143), .A2(new_n603), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1127), .A2(new_n1129), .A3(new_n1139), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1136), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT116), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1146), .A2(new_n1148), .A3(new_n1140), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1136), .A3(KEYINPUT116), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT117), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1146), .A2(new_n1148), .A3(new_n1140), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(new_n1151), .A4(new_n1150), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1146), .A2(KEYINPUT61), .A3(new_n1140), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT58), .B(G1341), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1041), .A2(G1996), .B1(new_n1063), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n552), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT59), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1160), .A2(new_n1163), .A3(new_n552), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g741(.A(KEYINPUT118), .B(new_n611), .C1(new_n1143), .C2(KEYINPUT60), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1085), .A2(new_n1142), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1063), .A2(new_n757), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n603), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n1167), .A2(new_n1172), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1166), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1147), .B1(new_n1157), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1119), .B(new_n1123), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g753(.A(KEYINPUT119), .B(new_n1147), .C1(new_n1157), .C2(new_n1175), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1105), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1087), .A2(new_n1002), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n872), .B(new_n757), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n826), .B(G1996), .ZN(new_n1183));
  INV_X1    g758(.A(new_n729), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n727), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n727), .A2(new_n1184), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n592), .B(new_n734), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1181), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1180), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1182), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1181), .B1(new_n1191), .B2(new_n863), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT46), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(new_n1181), .B2(new_n829), .ZN(new_n1194));
  NOR4_X1   g769(.A1(new_n1087), .A2(KEYINPUT46), .A3(G1996), .A4(new_n1002), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1192), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT47), .Z(new_n1197));
  NAND2_X1  g772(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1198));
  OAI22_X1  g773(.A1(new_n1198), .A2(new_n1185), .B1(G2067), .B2(new_n872), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1181), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT125), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1181), .A2(new_n734), .A3(new_n592), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT48), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1205));
  AOI211_X1 g780(.A(new_n1204), .B(new_n1205), .C1(new_n1181), .C2(new_n1187), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n1197), .A2(new_n1201), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1190), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n1210));
  OR2_X1    g784(.A1(new_n460), .A2(G227), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1211), .B1(new_n652), .B2(new_n654), .ZN(new_n1212));
  OAI21_X1  g786(.A(new_n1212), .B1(new_n701), .B2(new_n702), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n914), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n1215));
  AND3_X1   g789(.A1(new_n988), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n988), .B2(new_n1214), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n1210), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n988), .A2(new_n1214), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1219), .A2(KEYINPUT126), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n988), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1221));
  NAND3_X1  g795(.A1(new_n1220), .A2(KEYINPUT127), .A3(new_n1221), .ZN(new_n1222));
  AND2_X1   g796(.A1(new_n1218), .A2(new_n1222), .ZN(G308));
  NAND2_X1  g797(.A1(new_n1220), .A2(new_n1221), .ZN(G225));
endmodule


