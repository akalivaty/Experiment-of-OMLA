

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n551), .A2(n550), .ZN(n677) );
  NAND2_X2 U552 ( .A1(n678), .A2(n677), .ZN(n764) );
  NOR2_X2 U553 ( .A1(G2105), .A2(G2104), .ZN(n548) );
  NAND2_X2 U554 ( .A1(n565), .A2(n564), .ZN(n1015) );
  NOR2_X2 U555 ( .A1(n563), .A2(n562), .ZN(n565) );
  NOR2_X1 U556 ( .A1(n740), .A2(n763), .ZN(n742) );
  AND2_X1 U557 ( .A1(n529), .A2(G2105), .ZN(n994) );
  INV_X1 U558 ( .A(KEYINPUT17), .ZN(n547) );
  NOR2_X1 U559 ( .A1(n797), .A2(n521), .ZN(n798) );
  NOR2_X1 U560 ( .A1(G543), .A2(n539), .ZN(n534) );
  AND2_X1 U561 ( .A1(n760), .A2(n759), .ZN(n518) );
  XNOR2_X1 U562 ( .A(KEYINPUT69), .B(n575), .ZN(n519) );
  AND2_X1 U563 ( .A1(n553), .A2(n552), .ZN(n520) );
  AND2_X1 U564 ( .A1(n879), .A2(n811), .ZN(n521) );
  OR2_X1 U565 ( .A1(n763), .A2(n762), .ZN(n522) );
  OR2_X1 U566 ( .A1(n751), .A2(n750), .ZN(n523) );
  INV_X1 U567 ( .A(KEYINPUT31), .ZN(n716) );
  NOR2_X1 U568 ( .A1(G1966), .A2(n763), .ZN(n732) );
  INV_X1 U569 ( .A(KEYINPUT64), .ZN(n741) );
  INV_X1 U570 ( .A(n881), .ZN(n750) );
  NOR2_X1 U571 ( .A1(G164), .A2(G1384), .ZN(n765) );
  XNOR2_X1 U572 ( .A(KEYINPUT17), .B(n548), .ZN(n524) );
  NOR2_X1 U573 ( .A1(n621), .A2(n539), .ZN(n638) );
  INV_X1 U574 ( .A(n873), .ZN(n1016) );
  NOR2_X2 U575 ( .A1(G651), .A2(n621), .ZN(n647) );
  AND2_X1 U576 ( .A1(n528), .A2(n527), .ZN(n531) );
  NAND2_X1 U577 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U578 ( .A(n524), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n525), .A2(G138), .ZN(n526) );
  XNOR2_X1 U580 ( .A(n526), .B(KEYINPUT81), .ZN(n533) );
  INV_X1 U581 ( .A(G2104), .ZN(n529) );
  NOR2_X2 U582 ( .A1(G2105), .A2(n529), .ZN(n999) );
  NAND2_X1 U583 ( .A1(G102), .A2(n999), .ZN(n528) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n993) );
  NAND2_X1 U585 ( .A1(n993), .A2(G114), .ZN(n527) );
  NAND2_X1 U586 ( .A1(G126), .A2(n994), .ZN(n530) );
  NOR2_X1 U587 ( .A1(n533), .A2(n532), .ZN(G164) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n621) );
  NAND2_X1 U589 ( .A1(G51), .A2(n647), .ZN(n536) );
  INV_X1 U590 ( .A(G651), .ZN(n539) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n534), .Z(n641) );
  NAND2_X1 U592 ( .A1(G63), .A2(n641), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U594 ( .A(KEYINPUT6), .B(n537), .ZN(n545) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U596 ( .A1(n642), .A2(G89), .ZN(n538) );
  XNOR2_X1 U597 ( .A(n538), .B(KEYINPUT4), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G76), .A2(n638), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U600 ( .A(KEYINPUT5), .B(n542), .ZN(n543) );
  XNOR2_X1 U601 ( .A(KEYINPUT73), .B(n543), .ZN(n544) );
  NOR2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT7), .B(n546), .Z(G168) );
  XOR2_X1 U604 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U605 ( .A(n548), .B(n547), .ZN(n997) );
  NAND2_X1 U606 ( .A1(n997), .A2(G137), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G101), .A2(n999), .ZN(n549) );
  XOR2_X1 U608 ( .A(KEYINPUT23), .B(n549), .Z(n550) );
  NAND2_X1 U609 ( .A1(G113), .A2(n993), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G125), .A2(n994), .ZN(n552) );
  AND2_X1 U611 ( .A1(n677), .A2(n520), .ZN(G160) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U613 ( .A1(G7), .A2(G661), .ZN(n554) );
  XOR2_X1 U614 ( .A(n554), .B(KEYINPUT10), .Z(n1028) );
  NAND2_X1 U615 ( .A1(n1028), .A2(G567), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  NAND2_X1 U617 ( .A1(G56), .A2(n641), .ZN(n556) );
  XNOR2_X1 U618 ( .A(KEYINPUT14), .B(n556), .ZN(n557) );
  INV_X1 U619 ( .A(n557), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n642), .A2(G81), .ZN(n558) );
  XNOR2_X1 U621 ( .A(n558), .B(KEYINPUT12), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G68), .A2(n638), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT13), .B(n561), .Z(n562) );
  NAND2_X1 U625 ( .A1(n647), .A2(G43), .ZN(n564) );
  INV_X1 U626 ( .A(G860), .ZN(n595) );
  OR2_X1 U627 ( .A1(n1015), .A2(n595), .ZN(G153) );
  NAND2_X1 U628 ( .A1(G52), .A2(n647), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G64), .A2(n641), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G90), .A2(n642), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G77), .A2(n638), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U634 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U635 ( .A1(n572), .A2(n571), .ZN(G171) );
  INV_X1 U636 ( .A(G171), .ZN(G301) );
  NAND2_X1 U637 ( .A1(G66), .A2(n641), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G79), .A2(n638), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT70), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G54), .A2(n647), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT71), .B(n574), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G92), .A2(n642), .ZN(n575) );
  NOR2_X1 U643 ( .A1(n576), .A2(n519), .ZN(n577) );
  AND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT15), .ZN(n582) );
  XNOR2_X2 U647 ( .A(n582), .B(KEYINPUT72), .ZN(n873) );
  NOR2_X1 U648 ( .A1(n1016), .A2(G868), .ZN(n584) );
  INV_X1 U649 ( .A(G868), .ZN(n659) );
  NOR2_X1 U650 ( .A1(n659), .A2(G301), .ZN(n583) );
  NOR2_X1 U651 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G91), .A2(n642), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G78), .A2(n638), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G65), .A2(n641), .ZN(n587) );
  XNOR2_X1 U656 ( .A(KEYINPUT67), .B(n587), .ZN(n588) );
  NOR2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n647), .A2(G53), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(G299) );
  NOR2_X1 U660 ( .A1(G286), .A2(n659), .ZN(n593) );
  NOR2_X1 U661 ( .A1(G868), .A2(G299), .ZN(n592) );
  NOR2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U663 ( .A(KEYINPUT74), .B(n594), .ZN(G297) );
  NAND2_X1 U664 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n596), .A2(n873), .ZN(n597) );
  XNOR2_X1 U666 ( .A(n597), .B(KEYINPUT16), .ZN(n598) );
  XOR2_X1 U667 ( .A(KEYINPUT75), .B(n598), .Z(G148) );
  NOR2_X1 U668 ( .A1(G868), .A2(n1015), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n873), .A2(G868), .ZN(n599) );
  NOR2_X1 U670 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G123), .A2(n994), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n993), .A2(G111), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G135), .A2(n997), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G99), .A2(n999), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n986) );
  XNOR2_X1 U680 ( .A(n986), .B(G2096), .ZN(n609) );
  INV_X1 U681 ( .A(G2100), .ZN(n962) );
  NAND2_X1 U682 ( .A1(n609), .A2(n962), .ZN(G156) );
  NAND2_X1 U683 ( .A1(n873), .A2(G559), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n1015), .B(n610), .ZN(n656) );
  NOR2_X1 U685 ( .A1(n656), .A2(G860), .ZN(n617) );
  NAND2_X1 U686 ( .A1(G55), .A2(n647), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G67), .A2(n641), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G93), .A2(n642), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G80), .A2(n638), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n658) );
  XNOR2_X1 U693 ( .A(n617), .B(n658), .ZN(G145) );
  NAND2_X1 U694 ( .A1(G49), .A2(n647), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G74), .A2(G651), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n641), .A2(n620), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n621), .A2(G87), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(G288) );
  NAND2_X1 U700 ( .A1(n641), .A2(G60), .ZN(n630) );
  NAND2_X1 U701 ( .A1(G85), .A2(n642), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G72), .A2(n638), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G47), .A2(n647), .ZN(n626) );
  XNOR2_X1 U705 ( .A(KEYINPUT65), .B(n626), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n631), .B(KEYINPUT66), .ZN(G290) );
  NAND2_X1 U709 ( .A1(G88), .A2(n642), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G75), .A2(n638), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G50), .A2(n647), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G62), .A2(n641), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U715 ( .A1(n637), .A2(n636), .ZN(G166) );
  XOR2_X1 U716 ( .A(KEYINPUT76), .B(KEYINPUT2), .Z(n640) );
  NAND2_X1 U717 ( .A1(G73), .A2(n638), .ZN(n639) );
  XNOR2_X1 U718 ( .A(n640), .B(n639), .ZN(n646) );
  NAND2_X1 U719 ( .A1(G61), .A2(n641), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G86), .A2(n642), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n647), .A2(G48), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(G305) );
  XNOR2_X1 U725 ( .A(n658), .B(G288), .ZN(n655) );
  XOR2_X1 U726 ( .A(KEYINPUT77), .B(KEYINPUT19), .Z(n651) );
  XNOR2_X1 U727 ( .A(G290), .B(G166), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U729 ( .A(G299), .B(n652), .Z(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(G305), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(n1014) );
  XOR2_X1 U732 ( .A(n656), .B(n1014), .Z(n657) );
  NAND2_X1 U733 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U736 ( .A(KEYINPUT78), .B(n662), .Z(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U743 ( .A(KEYINPUT68), .B(G57), .Z(G237) );
  NAND2_X1 U744 ( .A1(G661), .A2(G483), .ZN(n675) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(KEYINPUT79), .Z(n668) );
  NAND2_X1 U746 ( .A1(G132), .A2(G82), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U748 ( .A1(n669), .A2(G218), .ZN(n670) );
  NAND2_X1 U749 ( .A1(G96), .A2(n670), .ZN(n949) );
  NAND2_X1 U750 ( .A1(n949), .A2(G2106), .ZN(n674) );
  NAND2_X1 U751 ( .A1(G108), .A2(G120), .ZN(n671) );
  NOR2_X1 U752 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G69), .A2(n672), .ZN(n948) );
  NAND2_X1 U754 ( .A1(G567), .A2(n948), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(n950) );
  NOR2_X1 U756 ( .A1(n675), .A2(n950), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n676), .B(KEYINPUT80), .ZN(n819) );
  NAND2_X1 U758 ( .A1(G36), .A2(n819), .ZN(G176) );
  XOR2_X1 U759 ( .A(G166), .B(KEYINPUT82), .Z(G303) );
  INV_X1 U760 ( .A(n765), .ZN(n679) );
  AND2_X1 U761 ( .A1(G40), .A2(n520), .ZN(n678) );
  NOR2_X4 U762 ( .A1(n679), .A2(n764), .ZN(n703) );
  INV_X2 U763 ( .A(n703), .ZN(n721) );
  NAND2_X1 U764 ( .A1(G1348), .A2(n721), .ZN(n681) );
  NAND2_X1 U765 ( .A1(G2067), .A2(n703), .ZN(n680) );
  NAND2_X1 U766 ( .A1(n681), .A2(n680), .ZN(n687) );
  AND2_X1 U767 ( .A1(n721), .A2(G1341), .ZN(n682) );
  NOR2_X1 U768 ( .A1(n682), .A2(n1015), .ZN(n685) );
  INV_X1 U769 ( .A(G1996), .ZN(n974) );
  NOR2_X1 U770 ( .A1(n721), .A2(n974), .ZN(n683) );
  XOR2_X1 U771 ( .A(n683), .B(KEYINPUT26), .Z(n684) );
  AND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n688) );
  NOR2_X1 U773 ( .A1(n873), .A2(n688), .ZN(n686) );
  NOR2_X1 U774 ( .A1(n687), .A2(n686), .ZN(n690) );
  AND2_X1 U775 ( .A1(n873), .A2(n688), .ZN(n689) );
  NOR2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n696) );
  NAND2_X1 U777 ( .A1(n721), .A2(G1956), .ZN(n693) );
  NAND2_X1 U778 ( .A1(n703), .A2(G2072), .ZN(n691) );
  XOR2_X1 U779 ( .A(KEYINPUT27), .B(n691), .Z(n692) );
  NAND2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U781 ( .A(n694), .B(KEYINPUT91), .ZN(n697) );
  INV_X1 U782 ( .A(G299), .ZN(n868) );
  NAND2_X1 U783 ( .A1(n697), .A2(n868), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U785 ( .A1(n697), .A2(n868), .ZN(n698) );
  XOR2_X1 U786 ( .A(n698), .B(KEYINPUT28), .Z(n699) );
  NAND2_X1 U787 ( .A1(n700), .A2(n699), .ZN(n702) );
  XOR2_X1 U788 ( .A(KEYINPUT29), .B(KEYINPUT92), .Z(n701) );
  XNOR2_X1 U789 ( .A(n702), .B(n701), .ZN(n708) );
  NOR2_X1 U790 ( .A1(n703), .A2(G1961), .ZN(n704) );
  XNOR2_X1 U791 ( .A(n704), .B(KEYINPUT90), .ZN(n706) );
  XOR2_X1 U792 ( .A(G2078), .B(KEYINPUT25), .Z(n917) );
  NOR2_X1 U793 ( .A1(n721), .A2(n917), .ZN(n705) );
  NOR2_X1 U794 ( .A1(n706), .A2(n705), .ZN(n709) );
  OR2_X1 U795 ( .A1(n709), .A2(G301), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n708), .A2(n707), .ZN(n719) );
  NAND2_X1 U797 ( .A1(n709), .A2(G301), .ZN(n710) );
  XNOR2_X1 U798 ( .A(n710), .B(KEYINPUT93), .ZN(n715) );
  NAND2_X1 U799 ( .A1(G8), .A2(n721), .ZN(n763) );
  NOR2_X1 U800 ( .A1(G2084), .A2(n721), .ZN(n729) );
  NOR2_X1 U801 ( .A1(n732), .A2(n729), .ZN(n711) );
  NAND2_X1 U802 ( .A1(G8), .A2(n711), .ZN(n712) );
  XNOR2_X1 U803 ( .A(n712), .B(KEYINPUT30), .ZN(n713) );
  NOR2_X1 U804 ( .A1(n713), .A2(G168), .ZN(n714) );
  NOR2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n717) );
  XNOR2_X1 U806 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n719), .A2(n718), .ZN(n730) );
  NAND2_X1 U808 ( .A1(n730), .A2(G286), .ZN(n720) );
  XNOR2_X1 U809 ( .A(n720), .B(KEYINPUT94), .ZN(n726) );
  NOR2_X1 U810 ( .A1(G1971), .A2(n763), .ZN(n723) );
  NOR2_X1 U811 ( .A1(G2090), .A2(n721), .ZN(n722) );
  NOR2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n724), .A2(G303), .ZN(n725) );
  NAND2_X1 U814 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U815 ( .A1(n727), .A2(G8), .ZN(n728) );
  XNOR2_X1 U816 ( .A(n728), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U817 ( .A1(G8), .A2(n729), .ZN(n734) );
  INV_X1 U818 ( .A(n730), .ZN(n731) );
  NOR2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U820 ( .A1(n734), .A2(n733), .ZN(n754) );
  NAND2_X1 U821 ( .A1(G1976), .A2(G288), .ZN(n864) );
  AND2_X1 U822 ( .A1(n754), .A2(n864), .ZN(n735) );
  AND2_X1 U823 ( .A1(n753), .A2(n735), .ZN(n739) );
  INV_X1 U824 ( .A(n864), .ZN(n737) );
  NOR2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n746) );
  NOR2_X1 U826 ( .A1(G303), .A2(G1971), .ZN(n736) );
  NOR2_X1 U827 ( .A1(n746), .A2(n736), .ZN(n865) );
  NOR2_X1 U828 ( .A1(n737), .A2(n865), .ZN(n738) );
  NOR2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U830 ( .A(n742), .B(n741), .ZN(n744) );
  INV_X1 U831 ( .A(KEYINPUT33), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT95), .ZN(n752) );
  NAND2_X1 U834 ( .A1(n746), .A2(KEYINPUT33), .ZN(n747) );
  XNOR2_X1 U835 ( .A(KEYINPUT96), .B(n747), .ZN(n748) );
  NOR2_X1 U836 ( .A1(n763), .A2(n748), .ZN(n749) );
  XOR2_X1 U837 ( .A(KEYINPUT97), .B(n749), .Z(n751) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n881) );
  OR2_X2 U839 ( .A1(n752), .A2(n523), .ZN(n760) );
  NAND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n757) );
  NOR2_X1 U841 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U842 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n758), .A2(n763), .ZN(n759) );
  NOR2_X1 U845 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XOR2_X1 U846 ( .A(n761), .B(KEYINPUT24), .Z(n762) );
  NAND2_X1 U847 ( .A1(n518), .A2(n522), .ZN(n799) );
  NOR2_X1 U848 ( .A1(n765), .A2(n764), .ZN(n811) );
  NAND2_X1 U849 ( .A1(G140), .A2(n997), .ZN(n767) );
  NAND2_X1 U850 ( .A1(G104), .A2(n999), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U852 ( .A(KEYINPUT34), .B(n768), .ZN(n774) );
  NAND2_X1 U853 ( .A1(n994), .A2(G128), .ZN(n769) );
  XNOR2_X1 U854 ( .A(n769), .B(KEYINPUT84), .ZN(n771) );
  NAND2_X1 U855 ( .A1(G116), .A2(n993), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U857 ( .A(n772), .B(KEYINPUT35), .Z(n773) );
  NOR2_X1 U858 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U859 ( .A(KEYINPUT36), .B(n775), .Z(n776) );
  XNOR2_X1 U860 ( .A(KEYINPUT85), .B(n776), .ZN(n1011) );
  XNOR2_X1 U861 ( .A(G2067), .B(KEYINPUT37), .ZN(n809) );
  NOR2_X1 U862 ( .A1(n1011), .A2(n809), .ZN(n834) );
  NAND2_X1 U863 ( .A1(n811), .A2(n834), .ZN(n807) );
  NAND2_X1 U864 ( .A1(G131), .A2(n997), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G95), .A2(n999), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G107), .A2(n993), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G119), .A2(n994), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n988) );
  XOR2_X1 U871 ( .A(G1991), .B(KEYINPUT86), .Z(n921) );
  NOR2_X1 U872 ( .A1(n988), .A2(n921), .ZN(n794) );
  NAND2_X1 U873 ( .A1(G117), .A2(n993), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G129), .A2(n994), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G105), .A2(n999), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n785), .B(KEYINPUT87), .ZN(n786) );
  XNOR2_X1 U878 ( .A(n786), .B(KEYINPUT38), .ZN(n787) );
  NOR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U880 ( .A(n789), .B(KEYINPUT88), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G141), .A2(n997), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U883 ( .A(KEYINPUT89), .B(n792), .ZN(n800) );
  NOR2_X1 U884 ( .A1(n974), .A2(n800), .ZN(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n836) );
  INV_X1 U886 ( .A(n836), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n795), .A2(n811), .ZN(n801) );
  NAND2_X1 U888 ( .A1(n807), .A2(n801), .ZN(n797) );
  XOR2_X1 U889 ( .A(G1986), .B(G290), .Z(n796) );
  XNOR2_X1 U890 ( .A(KEYINPUT83), .B(n796), .ZN(n879) );
  NAND2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n814) );
  INV_X1 U892 ( .A(n800), .ZN(n1008) );
  NOR2_X1 U893 ( .A1(G1996), .A2(n1008), .ZN(n839) );
  INV_X1 U894 ( .A(n801), .ZN(n804) );
  AND2_X1 U895 ( .A1(n988), .A2(n921), .ZN(n830) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U897 ( .A1(n830), .A2(n802), .ZN(n803) );
  NOR2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n839), .A2(n805), .ZN(n806) );
  XNOR2_X1 U900 ( .A(n806), .B(KEYINPUT39), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n1011), .A2(n809), .ZN(n845) );
  NAND2_X1 U903 ( .A1(n810), .A2(n845), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n816) );
  XNOR2_X1 U906 ( .A(KEYINPUT98), .B(KEYINPUT40), .ZN(n815) );
  XNOR2_X1 U907 ( .A(n816), .B(n815), .ZN(G329) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n1028), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(G188) );
  NAND2_X1 U914 ( .A1(n994), .A2(G124), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n820), .B(KEYINPUT44), .ZN(n822) );
  NAND2_X1 U916 ( .A1(G136), .A2(n997), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT103), .ZN(n825) );
  NAND2_X1 U919 ( .A1(G100), .A2(n999), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n993), .A2(G112), .ZN(n826) );
  XOR2_X1 U922 ( .A(KEYINPUT104), .B(n826), .Z(n827) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT105), .B(n829), .Z(G162) );
  XNOR2_X1 U925 ( .A(G160), .B(G2084), .ZN(n832) );
  NOR2_X1 U926 ( .A1(n830), .A2(n986), .ZN(n831) );
  NAND2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U930 ( .A(KEYINPUT112), .B(n837), .ZN(n843) );
  XOR2_X1 U931 ( .A(G2090), .B(G162), .Z(n838) );
  NOR2_X1 U932 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U933 ( .A(KEYINPUT113), .B(n840), .Z(n841) );
  XNOR2_X1 U934 ( .A(n841), .B(KEYINPUT51), .ZN(n842) );
  NOR2_X1 U935 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U936 ( .A(n844), .B(KEYINPUT114), .ZN(n846) );
  NAND2_X1 U937 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U938 ( .A(KEYINPUT115), .B(n847), .Z(n859) );
  NAND2_X1 U939 ( .A1(G139), .A2(n997), .ZN(n849) );
  NAND2_X1 U940 ( .A1(G103), .A2(n999), .ZN(n848) );
  NAND2_X1 U941 ( .A1(n849), .A2(n848), .ZN(n854) );
  NAND2_X1 U942 ( .A1(G115), .A2(n993), .ZN(n851) );
  NAND2_X1 U943 ( .A1(G127), .A2(n994), .ZN(n850) );
  NAND2_X1 U944 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U945 ( .A(KEYINPUT47), .B(n852), .Z(n853) );
  NOR2_X1 U946 ( .A1(n854), .A2(n853), .ZN(n983) );
  XOR2_X1 U947 ( .A(G2072), .B(n983), .Z(n856) );
  XOR2_X1 U948 ( .A(G164), .B(G2078), .Z(n855) );
  NOR2_X1 U949 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U950 ( .A(KEYINPUT50), .B(n857), .Z(n858) );
  NOR2_X1 U951 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U952 ( .A(KEYINPUT52), .B(n860), .ZN(n861) );
  INV_X1 U953 ( .A(KEYINPUT55), .ZN(n938) );
  NAND2_X1 U954 ( .A1(n861), .A2(n938), .ZN(n862) );
  NAND2_X1 U955 ( .A1(n862), .A2(G29), .ZN(n946) );
  XNOR2_X1 U956 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n863) );
  XOR2_X1 U957 ( .A(G16), .B(n863), .Z(n887) );
  AND2_X1 U958 ( .A1(G303), .A2(G1971), .ZN(n867) );
  NAND2_X1 U959 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U960 ( .A1(n867), .A2(n866), .ZN(n877) );
  XOR2_X1 U961 ( .A(G301), .B(G1961), .Z(n872) );
  XOR2_X1 U962 ( .A(n868), .B(G1956), .Z(n870) );
  XNOR2_X1 U963 ( .A(n1015), .B(G1341), .ZN(n869) );
  NOR2_X1 U964 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U965 ( .A1(n872), .A2(n871), .ZN(n875) );
  XOR2_X1 U966 ( .A(n873), .B(G1348), .Z(n874) );
  NOR2_X1 U967 ( .A1(n875), .A2(n874), .ZN(n876) );
  NAND2_X1 U968 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U969 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U970 ( .A(KEYINPUT122), .B(n880), .ZN(n885) );
  XNOR2_X1 U971 ( .A(G1966), .B(G168), .ZN(n882) );
  NAND2_X1 U972 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U973 ( .A(KEYINPUT57), .B(n883), .ZN(n884) );
  NAND2_X1 U974 ( .A1(n885), .A2(n884), .ZN(n886) );
  NAND2_X1 U975 ( .A1(n887), .A2(n886), .ZN(n915) );
  INV_X1 U976 ( .A(G16), .ZN(n913) );
  XOR2_X1 U977 ( .A(G1976), .B(G23), .Z(n889) );
  XOR2_X1 U978 ( .A(G1971), .B(G22), .Z(n888) );
  NAND2_X1 U979 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U980 ( .A(G24), .B(G1986), .ZN(n890) );
  NOR2_X1 U981 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U982 ( .A(KEYINPUT58), .B(n892), .Z(n910) );
  XOR2_X1 U983 ( .A(G1966), .B(G21), .Z(n904) );
  XOR2_X1 U984 ( .A(G1348), .B(KEYINPUT59), .Z(n893) );
  XNOR2_X1 U985 ( .A(G4), .B(n893), .ZN(n901) );
  XOR2_X1 U986 ( .A(G1956), .B(G20), .Z(n896) );
  XOR2_X1 U987 ( .A(G19), .B(KEYINPUT124), .Z(n894) );
  XNOR2_X1 U988 ( .A(n894), .B(G1341), .ZN(n895) );
  NAND2_X1 U989 ( .A1(n896), .A2(n895), .ZN(n898) );
  XNOR2_X1 U990 ( .A(G6), .B(G1981), .ZN(n897) );
  NOR2_X1 U991 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n899), .B(KEYINPUT125), .ZN(n900) );
  NOR2_X1 U993 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U994 ( .A(KEYINPUT60), .B(n902), .ZN(n903) );
  NAND2_X1 U995 ( .A1(n904), .A2(n903), .ZN(n907) );
  XOR2_X1 U996 ( .A(KEYINPUT123), .B(G1961), .Z(n905) );
  XNOR2_X1 U997 ( .A(G5), .B(n905), .ZN(n906) );
  NOR2_X1 U998 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U999 ( .A(KEYINPUT126), .B(n908), .Z(n909) );
  NOR2_X1 U1000 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1001 ( .A(KEYINPUT61), .B(n911), .ZN(n912) );
  NAND2_X1 U1002 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1003 ( .A1(n915), .A2(n914), .ZN(n944) );
  XNOR2_X1 U1004 ( .A(G2090), .B(G35), .ZN(n931) );
  XOR2_X1 U1005 ( .A(G2072), .B(G33), .Z(n916) );
  NAND2_X1 U1006 ( .A1(G28), .A2(n916), .ZN(n927) );
  XOR2_X1 U1007 ( .A(n974), .B(G32), .Z(n919) );
  XNOR2_X1 U1008 ( .A(n917), .B(G27), .ZN(n918) );
  NOR2_X1 U1009 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1010 ( .A(KEYINPUT116), .B(n920), .ZN(n925) );
  XOR2_X1 U1011 ( .A(n921), .B(G25), .Z(n923) );
  XNOR2_X1 U1012 ( .A(G2067), .B(G26), .ZN(n922) );
  NOR2_X1 U1013 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1014 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1015 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1016 ( .A(KEYINPUT117), .B(n928), .Z(n929) );
  XNOR2_X1 U1017 ( .A(n929), .B(KEYINPUT53), .ZN(n930) );
  NOR2_X1 U1018 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1019 ( .A(KEYINPUT118), .B(n932), .ZN(n935) );
  XOR2_X1 U1020 ( .A(G2084), .B(G34), .Z(n933) );
  XNOR2_X1 U1021 ( .A(KEYINPUT54), .B(n933), .ZN(n934) );
  NAND2_X1 U1022 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1023 ( .A(n936), .B(KEYINPUT119), .ZN(n937) );
  XOR2_X1 U1024 ( .A(n938), .B(n937), .Z(n940) );
  INV_X1 U1025 ( .A(G29), .ZN(n939) );
  NAND2_X1 U1026 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1027 ( .A1(G11), .A2(n941), .ZN(n942) );
  XNOR2_X1 U1028 ( .A(KEYINPUT120), .B(n942), .ZN(n943) );
  NOR2_X1 U1029 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1030 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1031 ( .A(KEYINPUT62), .B(n947), .Z(G311) );
  XNOR2_X1 U1032 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1033 ( .A(G132), .ZN(G219) );
  INV_X1 U1034 ( .A(G120), .ZN(G236) );
  INV_X1 U1035 ( .A(G108), .ZN(G238) );
  INV_X1 U1036 ( .A(G96), .ZN(G221) );
  INV_X1 U1037 ( .A(G82), .ZN(G220) );
  INV_X1 U1038 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(G325) );
  INV_X1 U1040 ( .A(G325), .ZN(G261) );
  INV_X1 U1041 ( .A(n950), .ZN(G319) );
  XOR2_X1 U1042 ( .A(G2454), .B(KEYINPUT99), .Z(n952) );
  XNOR2_X1 U1043 ( .A(G1348), .B(G2446), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(n952), .B(n951), .ZN(n959) );
  XOR2_X1 U1045 ( .A(G2451), .B(G2430), .Z(n954) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G2427), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n954), .B(n953), .ZN(n955) );
  XOR2_X1 U1048 ( .A(n955), .B(G2443), .Z(n957) );
  XNOR2_X1 U1049 ( .A(G2435), .B(G2438), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n957), .B(n956), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n959), .B(n958), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n960), .A2(G14), .ZN(n961) );
  XOR2_X1 U1053 ( .A(KEYINPUT100), .B(n961), .Z(G401) );
  XNOR2_X1 U1054 ( .A(G2678), .B(n962), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G2067), .B(G2084), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(n964), .B(n963), .ZN(n965) );
  XOR2_X1 U1057 ( .A(n965), .B(KEYINPUT101), .Z(n967) );
  XNOR2_X1 U1058 ( .A(G2090), .B(KEYINPUT42), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n967), .B(n966), .ZN(n971) );
  XOR2_X1 U1060 ( .A(G2096), .B(KEYINPUT43), .Z(n969) );
  XNOR2_X1 U1061 ( .A(G2078), .B(G2072), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1063 ( .A(n971), .B(n970), .Z(G227) );
  XNOR2_X1 U1064 ( .A(G1986), .B(G1981), .ZN(n982) );
  XOR2_X1 U1065 ( .A(G1971), .B(G1956), .Z(n973) );
  XNOR2_X1 U1066 ( .A(G1991), .B(G1966), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n973), .B(n972), .ZN(n978) );
  XOR2_X1 U1068 ( .A(KEYINPUT102), .B(KEYINPUT41), .Z(n976) );
  XOR2_X1 U1069 ( .A(n974), .B(G1961), .Z(n975) );
  XNOR2_X1 U1070 ( .A(n976), .B(n975), .ZN(n977) );
  XOR2_X1 U1071 ( .A(n978), .B(n977), .Z(n980) );
  XNOR2_X1 U1072 ( .A(G1976), .B(G2474), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n980), .B(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n982), .B(n981), .ZN(G229) );
  XNOR2_X1 U1075 ( .A(G164), .B(n983), .ZN(n992) );
  XOR2_X1 U1076 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n985), .B(n984), .ZN(n987) );
  XOR2_X1 U1079 ( .A(n987), .B(n986), .Z(n990) );
  XNOR2_X1 U1080 ( .A(G160), .B(n988), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n992), .B(n991), .ZN(n1007) );
  NAND2_X1 U1083 ( .A1(G118), .A2(n993), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(G130), .A2(n994), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n1005) );
  NAND2_X1 U1086 ( .A1(n997), .A2(G142), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n998), .B(KEYINPUT106), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(G106), .A2(n999), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT45), .B(n1002), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT107), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(n1007), .B(n1006), .Z(n1010) );
  XOR2_X1 U1094 ( .A(n1008), .B(G162), .Z(n1009) );
  XNOR2_X1 U1095 ( .A(n1010), .B(n1009), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NOR2_X1 U1097 ( .A1(G37), .A2(n1013), .ZN(G395) );
  XNOR2_X1 U1098 ( .A(n1015), .B(n1014), .ZN(n1018) );
  XOR2_X1 U1099 ( .A(G301), .B(n1016), .Z(n1017) );
  XNOR2_X1 U1100 ( .A(n1018), .B(n1017), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(n1019), .B(G286), .ZN(n1020) );
  NOR2_X1 U1102 ( .A1(G37), .A2(n1020), .ZN(n1021) );
  XNOR2_X1 U1103 ( .A(KEYINPUT110), .B(n1021), .ZN(G397) );
  NOR2_X1 U1104 ( .A1(G227), .A2(G229), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(n1022), .B(KEYINPUT49), .ZN(n1023) );
  NOR2_X1 U1106 ( .A1(G401), .A2(n1023), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(G319), .A2(n1024), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(KEYINPUT111), .B(n1025), .ZN(n1027) );
  NOR2_X1 U1109 ( .A1(G395), .A2(G397), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(G225) );
  INV_X1 U1111 ( .A(G225), .ZN(G308) );
  INV_X1 U1112 ( .A(n1028), .ZN(G223) );
endmodule

