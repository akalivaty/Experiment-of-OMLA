//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  OR2_X1    g000(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  AOI21_X1  g002(.A(G36gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n205), .A2(new_n206), .A3(G29gat), .ZN(new_n207));
  OR3_X1    g006(.A1(new_n204), .A2(KEYINPUT15), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT15), .B1(new_n204), .B2(new_n207), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n209), .B2(new_n210), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT17), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(G1gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G1gat), .B2(new_n214), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(G8gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n212), .A2(new_n218), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT18), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n220), .A2(KEYINPUT18), .A3(new_n221), .A4(new_n222), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n212), .B(new_n218), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n221), .B(KEYINPUT13), .Z(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G113gat), .B(G141gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(G169gat), .B(G197gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT12), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n225), .A2(new_n226), .A3(new_n229), .A4(new_n236), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G141gat), .ZN(new_n242));
  INV_X1    g041(.A(G148gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n245));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G162gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G155gat), .ZN(new_n249));
  INV_X1    g048(.A(G155gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G162gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT78), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n247), .A2(KEYINPUT78), .A3(new_n252), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT79), .ZN(new_n258));
  AND2_X1   g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n244), .A2(KEYINPUT79), .A3(new_n246), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n265));
  OAI21_X1  g064(.A(G155gat), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT2), .ZN(new_n267));
  INV_X1    g066(.A(new_n252), .ZN(new_n268));
  AND4_X1   g067(.A1(new_n257), .A2(new_n263), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n252), .B1(new_n261), .B2(new_n262), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n257), .B1(new_n270), .B2(new_n267), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n256), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n273));
  INV_X1    g072(.A(G113gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(G120gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  INV_X1    g075(.A(G120gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(G113gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n275), .A2(new_n278), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282));
  XNOR2_X1  g081(.A(G127gat), .B(G134gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n274), .A2(G120gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n277), .A2(G113gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n272), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT5), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n295), .B(new_n256), .C1(new_n269), .C2(new_n271), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n284), .A2(new_n289), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n290), .B(new_n256), .C1(new_n269), .C2(new_n271), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT4), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n298), .A2(new_n301), .A3(new_n292), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n293), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G1gat), .B(G29gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT0), .ZN(new_n307));
  XNOR2_X1  g106(.A(G57gat), .B(G85gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n299), .B(KEYINPUT4), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n311), .A2(KEYINPUT5), .A3(new_n292), .A4(new_n298), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n305), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT6), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n310), .B1(new_n305), .B2(new_n312), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT86), .B1(new_n316), .B2(new_n317), .ZN(new_n321));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G197gat), .B(G204gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(G211gat), .A2(G218gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n326), .B1(new_n325), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(new_n322), .A3(new_n324), .A4(new_n328), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT74), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G183gat), .ZN(new_n340));
  INV_X1    g139(.A(G190gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT28), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT28), .B1(new_n342), .B2(new_n343), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT65), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT65), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(G169gat), .A3(G176gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n358), .A2(KEYINPUT67), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT67), .B1(new_n358), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n347), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n359), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT24), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n349), .A2(new_n351), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(KEYINPUT64), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n341), .A2(G183gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n337), .A2(G190gat), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT24), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n365), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n365), .A2(new_n370), .A3(new_n373), .A4(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n362), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n380), .B(KEYINPUT75), .Z(new_n381));
  NOR2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n362), .B2(new_n378), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n336), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n362), .A2(new_n378), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n381), .ZN(new_n386));
  INV_X1    g185(.A(new_n380), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n386), .B(new_n334), .C1(new_n379), .C2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  NAND3_X1  g190(.A1(new_n384), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  OR3_X1    g192(.A1(new_n382), .A2(new_n336), .A3(new_n383), .ZN(new_n394));
  INV_X1    g193(.A(new_n379), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n395), .A2(new_n380), .B1(new_n385), .B2(new_n381), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n334), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT38), .B1(new_n397), .B2(KEYINPUT37), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n384), .A2(new_n388), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(KEYINPUT37), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n393), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n320), .A2(new_n321), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n320), .A2(KEYINPUT87), .A3(new_n321), .A4(new_n404), .ZN(new_n408));
  INV_X1    g207(.A(new_n403), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n399), .A2(KEYINPUT37), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT38), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT31), .B(G50gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT29), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n334), .B1(new_n296), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n255), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(new_n253), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n263), .A2(new_n267), .A3(new_n268), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT81), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n270), .A2(new_n257), .A3(new_n267), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT3), .B1(new_n334), .B2(new_n417), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n416), .B1(new_n418), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n334), .A2(new_n417), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n295), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n416), .B1(new_n429), .B2(new_n272), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n424), .B2(new_n295), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(new_n335), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n427), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n427), .B2(new_n432), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n415), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT82), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(new_n415), .C1(new_n434), .C2(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n427), .A2(new_n432), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n415), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n427), .B(new_n432), .C1(KEYINPUT83), .C2(new_n433), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n415), .B1(new_n441), .B2(new_n442), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n445), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n440), .A2(new_n451), .A3(KEYINPUT85), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT85), .B1(new_n440), .B2(new_n451), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT39), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n291), .A2(new_n292), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n311), .A2(new_n298), .ZN(new_n458));
  INV_X1    g257(.A(new_n292), .ZN(new_n459));
  AOI211_X1 g258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n456), .A3(new_n459), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n309), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n455), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n313), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n388), .A4(new_n391), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n401), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT77), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n392), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n392), .A2(new_n467), .A3(new_n468), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n460), .A2(new_n462), .A3(new_n455), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n464), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n454), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n412), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT70), .B1(new_n284), .B2(new_n289), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n284), .A2(KEYINPUT70), .A3(new_n289), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n342), .A2(new_n343), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT28), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n344), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n358), .A2(KEYINPUT67), .A3(new_n359), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n349), .A2(new_n351), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n357), .A2(new_n353), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n359), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n484), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n376), .A2(new_n377), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n478), .B(new_n480), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G227gat), .ZN(new_n494));
  INV_X1    g293(.A(G233gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT70), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n362), .A2(new_n497), .A3(new_n297), .A4(new_n378), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n493), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n493), .A2(KEYINPUT71), .A3(new_n496), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT33), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n496), .ZN(new_n506));
  AOI211_X1 g305(.A(new_n477), .B(new_n479), .C1(new_n362), .C2(new_n378), .ZN(new_n507));
  INV_X1    g306(.A(new_n498), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT34), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n496), .B1(new_n493), .B2(new_n498), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G15gat), .B(G43gat), .Z(new_n515));
  XNOR2_X1  g314(.A(G71gat), .B(G99gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n505), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n511), .B(KEYINPUT34), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT33), .B1(new_n501), .B2(new_n502), .ZN(new_n520));
  INV_X1    g319(.A(new_n517), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n503), .A2(KEYINPUT32), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n518), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n518), .B2(new_n522), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(KEYINPUT72), .A3(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n514), .B1(new_n505), .B2(new_n517), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n523), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n525), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n441), .A2(G22gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n427), .A2(new_n432), .A3(new_n433), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n438), .B1(new_n541), .B2(new_n415), .ZN(new_n542));
  INV_X1    g341(.A(new_n439), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n445), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT84), .B1(new_n449), .B2(new_n445), .ZN(new_n545));
  OAI22_X1  g344(.A1(new_n542), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n440), .A2(new_n451), .A3(KEYINPUT85), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n316), .ZN(new_n551));
  INV_X1    g350(.A(new_n317), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n315), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n401), .A2(KEYINPUT76), .A3(new_n465), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT76), .B1(new_n401), .B2(new_n465), .ZN(new_n555));
  INV_X1    g354(.A(new_n471), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n469), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n538), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n476), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n558), .B(new_n528), .C1(new_n452), .C2(new_n453), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT35), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n528), .B1(new_n452), .B2(new_n453), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n552), .A2(new_n319), .A3(new_n314), .A4(new_n313), .ZN(new_n565));
  INV_X1    g364(.A(new_n315), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n321), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT35), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n472), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT88), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n564), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n534), .B1(new_n548), .B2(new_n549), .ZN(new_n572));
  INV_X1    g371(.A(new_n466), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n573), .B(new_n568), .C1(new_n469), .C2(new_n556), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n574), .B1(new_n320), .B2(new_n321), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT88), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n563), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n241), .B1(new_n561), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT93), .Z(new_n580));
  INV_X1    g379(.A(KEYINPUT41), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G134gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(new_n248), .ZN(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT94), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n589), .A2(new_n591), .A3(G85gat), .A4(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n589), .A2(new_n591), .B1(G85gat), .B2(G92gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT95), .ZN(new_n600));
  XOR2_X1   g399(.A(G99gat), .B(G106gat), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n597), .B2(new_n598), .ZN(new_n604));
  INV_X1    g403(.A(new_n598), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(new_n602), .A3(new_n592), .A4(new_n596), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n606), .A3(KEYINPUT95), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n213), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n580), .A2(new_n581), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n603), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n212), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n587), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n585), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n587), .A3(new_n611), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n614), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n614), .B1(new_n612), .B2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(G71gat), .A2(G78gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G57gat), .B(G64gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT9), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G57gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(G64gat), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT90), .B(G57gat), .Z(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n629), .B2(G64gat), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n621), .B1(KEYINPUT9), .B2(new_n622), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n218), .B1(KEYINPUT21), .B2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT92), .Z(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G127gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n635), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G155gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n642), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT99), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n651));
  OAI211_X1 g450(.A(KEYINPUT10), .B(new_n626), .C1(new_n630), .C2(new_n631), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n610), .B2(new_n653), .ZN(new_n654));
  AOI211_X1 g453(.A(KEYINPUT97), .B(new_n652), .C1(new_n607), .C2(new_n603), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n604), .A2(new_n606), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(new_n632), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n610), .A2(new_n632), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT10), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n650), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n658), .A2(new_n659), .A3(G230gat), .A4(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(G120gat), .B(G148gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT98), .ZN(new_n665));
  XNOR2_X1  g464(.A(G176gat), .B(G204gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n648), .B1(new_n656), .B2(new_n660), .ZN(new_n669));
  INV_X1    g468(.A(new_n667), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n662), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n620), .A2(new_n647), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n578), .A2(new_n553), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g474(.A1(new_n578), .A2(new_n673), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n472), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(KEYINPUT42), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT101), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT42), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  INV_X1    g480(.A(G8gat), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n677), .A2(KEYINPUT100), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT100), .B1(new_n677), .B2(new_n682), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(new_n538), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n676), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n534), .A2(G15gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n676), .B2(new_n689), .ZN(G1326gat));
  OR3_X1    g489(.A1(new_n676), .A2(KEYINPUT102), .A3(new_n550), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT102), .B1(new_n676), .B2(new_n550), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n693), .B(new_n694), .Z(G1327gat));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  AOI211_X1 g495(.A(new_n559), .B(new_n538), .C1(new_n412), .C2(new_n475), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n577), .A2(KEYINPUT103), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n570), .B1(new_n564), .B2(new_n569), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n572), .A2(KEYINPUT88), .A3(new_n575), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n563), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n697), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n696), .B1(new_n704), .B2(new_n619), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n619), .B1(new_n561), .B2(new_n577), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT44), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n647), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n241), .A3(new_n672), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n553), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n706), .A2(new_n710), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G29gat), .A3(new_n712), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT45), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(G1328gat));
  OAI21_X1  g516(.A(G36gat), .B1(new_n711), .B2(new_n472), .ZN(new_n718));
  INV_X1    g517(.A(new_n472), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n206), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT46), .B1(new_n714), .B2(new_n720), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n714), .A2(KEYINPUT46), .A3(new_n720), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n718), .A2(new_n721), .A3(new_n722), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n538), .A3(new_n710), .A4(new_n707), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G43gat), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n534), .A2(G43gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n706), .A2(new_n710), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(KEYINPUT47), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(KEYINPUT104), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(G43gat), .B2(new_n724), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n730), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g530(.A1(new_n705), .A2(new_n454), .A3(new_n710), .A4(new_n707), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G50gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n714), .A2(G50gat), .A3(new_n550), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(KEYINPUT105), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n733), .B(new_n736), .C1(KEYINPUT105), .C2(new_n735), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(new_n732), .B2(G50gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(KEYINPUT48), .ZN(G1331gat));
  XNOR2_X1  g538(.A(new_n553), .B(KEYINPUT106), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n709), .A2(new_n241), .A3(new_n619), .A4(new_n672), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n704), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(new_n629), .ZN(G1332gat));
  NOR3_X1   g542(.A1(new_n704), .A2(new_n472), .A3(new_n741), .ZN(new_n744));
  NOR2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  AND2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n744), .B2(new_n745), .ZN(G1333gat));
  NOR2_X1   g547(.A1(new_n704), .A2(new_n741), .ZN(new_n749));
  INV_X1    g548(.A(G71gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n687), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n749), .A2(KEYINPUT107), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT107), .B1(new_n749), .B2(new_n751), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n704), .A2(new_n534), .A3(new_n741), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n752), .A2(new_n753), .B1(G71gat), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n749), .A2(new_n454), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  INV_X1    g557(.A(new_n672), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n709), .A2(new_n240), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n708), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n712), .ZN(new_n762));
  AOI221_X4 g561(.A(KEYINPUT103), .B1(new_n562), .B2(KEYINPUT35), .C1(new_n699), .C2(new_n700), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n702), .B1(new_n701), .B2(new_n563), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n561), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n709), .A2(new_n240), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n620), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n553), .A2(new_n594), .A3(new_n672), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n762), .B1(new_n771), .B2(new_n772), .ZN(G1336gat));
  AND3_X1   g572(.A1(new_n767), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT51), .B1(new_n767), .B2(KEYINPUT109), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n472), .A2(G92gat), .A3(new_n759), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT108), .Z(new_n777));
  NOR3_X1   g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n705), .A2(new_n719), .A3(new_n707), .A4(new_n760), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT52), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(G92gat), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n783));
  INV_X1    g582(.A(new_n776), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n782), .B(new_n783), .C1(new_n771), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(G1337gat));
  OAI21_X1  g585(.A(G99gat), .B1(new_n761), .B2(new_n687), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n534), .A2(G99gat), .A3(new_n759), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n771), .B2(new_n788), .ZN(G1338gat));
  OR3_X1    g588(.A1(new_n550), .A2(G106gat), .A3(new_n759), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT111), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT112), .Z(new_n792));
  NOR3_X1   g591(.A1(new_n774), .A2(new_n775), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n705), .A2(new_n454), .A3(new_n707), .A4(new_n760), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT53), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n769), .B2(new_n770), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(G106gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(G1339gat));
  OR2_X1    g600(.A1(new_n654), .A2(new_n655), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n658), .A2(new_n659), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT10), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n805), .A3(new_n649), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n669), .A3(KEYINPUT54), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(new_n650), .C1(new_n656), .C2(new_n660), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(KEYINPUT113), .A3(new_n667), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT113), .B1(new_n809), .B2(new_n667), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT55), .B(new_n807), .C1(new_n811), .C2(new_n812), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n815), .A2(new_n240), .A3(new_n671), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n227), .A2(new_n228), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT114), .Z(new_n819));
  AOI21_X1  g618(.A(new_n221), .B1(new_n220), .B2(new_n222), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n235), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n239), .A3(new_n672), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n620), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n815), .A2(new_n671), .A3(new_n816), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n239), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n824), .A2(new_n619), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n647), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n673), .A2(new_n241), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n740), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n829), .A2(new_n472), .A3(new_n572), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n240), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n454), .B1(new_n827), .B2(new_n828), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n832), .A2(new_n472), .A3(new_n553), .A4(new_n528), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n274), .A3(new_n241), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n831), .A2(new_n834), .ZN(G1340gat));
  NAND3_X1  g634(.A1(new_n830), .A2(new_n277), .A3(new_n672), .ZN(new_n836));
  OAI21_X1  g635(.A(G120gat), .B1(new_n833), .B2(new_n759), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT115), .Z(G1341gat));
  NAND3_X1  g638(.A1(new_n830), .A2(new_n640), .A3(new_n709), .ZN(new_n840));
  OAI21_X1  g639(.A(G127gat), .B1(new_n833), .B2(new_n647), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1342gat));
  NAND3_X1  g641(.A1(new_n830), .A2(new_n583), .A3(new_n620), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n833), .B2(new_n619), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1343gat));
  NAND2_X1  g646(.A1(new_n553), .A2(new_n472), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n538), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n454), .A2(KEYINPUT57), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  INV_X1    g650(.A(new_n807), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n809), .A2(new_n667), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(new_n810), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n671), .B1(new_n856), .B2(KEYINPUT55), .ZN(new_n857));
  INV_X1    g656(.A(new_n816), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n851), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n815), .A2(KEYINPUT116), .A3(new_n671), .A4(new_n816), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n240), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n620), .B1(new_n861), .B2(new_n822), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n647), .B1(new_n862), .B2(new_n826), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n850), .B1(new_n863), .B2(new_n828), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n827), .A2(new_n828), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n865), .B2(new_n454), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n849), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G141gat), .B1(new_n867), .B2(new_n241), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n538), .A2(new_n550), .A3(new_n719), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n829), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(G141gat), .A3(new_n241), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT117), .B(new_n849), .C1(new_n864), .C2(new_n866), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n240), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n871), .B1(new_n877), .B2(G141gat), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(new_n870), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n243), .A3(new_n672), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n759), .B1(new_n849), .B2(KEYINPUT118), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(KEYINPUT118), .B2(new_n849), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  INV_X1    g685(.A(new_n826), .ZN(new_n887));
  INV_X1    g686(.A(new_n822), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n241), .B1(new_n824), .B2(new_n851), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n860), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n890), .B2(new_n620), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n891), .A2(new_n647), .B1(new_n241), .B2(new_n673), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n892), .B2(new_n550), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n865), .A2(KEYINPUT57), .A3(new_n454), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT119), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n243), .B1(new_n895), .B2(KEYINPUT119), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n883), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n883), .A2(G148gat), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n875), .A2(new_n876), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n672), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n882), .B1(new_n898), .B2(new_n901), .ZN(G1345gat));
  NAND3_X1  g701(.A1(new_n881), .A2(new_n250), .A3(new_n709), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n900), .A2(new_n709), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n250), .ZN(G1346gat));
  NAND3_X1  g704(.A1(new_n875), .A2(new_n620), .A3(new_n876), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n264), .A2(new_n265), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n881), .A2(new_n907), .A3(new_n620), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1347gat));
  NAND2_X1  g714(.A1(new_n740), .A2(new_n719), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n534), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n832), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(new_n355), .A3(new_n241), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n472), .B(new_n553), .C1(new_n827), .C2(new_n828), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n572), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT121), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n240), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n920), .B1(new_n924), .B2(new_n355), .ZN(G1348gat));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n356), .A3(new_n672), .ZN(new_n926));
  OAI21_X1  g725(.A(G176gat), .B1(new_n919), .B2(new_n759), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1349gat));
  NAND2_X1  g727(.A1(new_n338), .A2(new_n340), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n922), .A2(new_n929), .A3(new_n647), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT122), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n337), .B1(new_n918), .B2(new_n709), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n934), .B1(new_n932), .B2(KEYINPUT60), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n931), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1350gat));
  AOI21_X1  g737(.A(new_n341), .B1(new_n918), .B2(new_n620), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT61), .Z(new_n940));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n341), .A3(new_n620), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n538), .A2(new_n550), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n921), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n240), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n916), .A2(new_n538), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT124), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n947), .B1(new_n893), .B2(new_n894), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n240), .A2(G197gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1352gat));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n944), .A2(new_n951), .A3(new_n672), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  AND2_X1   g752(.A1(new_n948), .A2(new_n672), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n951), .B2(new_n954), .ZN(G1353gat));
  INV_X1    g754(.A(G211gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n893), .A2(new_n894), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n916), .A2(new_n538), .A3(new_n647), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT63), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n956), .A3(new_n709), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1354gat));
  NAND3_X1  g761(.A1(new_n921), .A2(new_n620), .A3(new_n943), .ZN(new_n963));
  INV_X1    g762(.A(G218gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT125), .ZN(new_n966));
  OAI211_X1 g765(.A(G218gat), .B(new_n620), .C1(new_n948), .C2(KEYINPUT126), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  AOI211_X1 g767(.A(new_n968), .B(new_n947), .C1(new_n893), .C2(new_n894), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g771(.A(KEYINPUT127), .B(new_n966), .C1(new_n967), .C2(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


