//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(G469), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT78), .ZN(new_n192));
  INV_X1    g006(.A(G227), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n192), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT79), .A2(G104), .ZN(new_n200));
  AOI21_X1  g014(.A(G107), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(G101), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT3), .A2(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT3), .A2(G107), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(G104), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n202), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n209), .A3(new_n200), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n204), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT80), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT1), .B1(new_n215), .B2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(G146), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  OAI211_X1 g033(.A(G128), .B(new_n216), .C1(new_n217), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(G146), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n221), .B(new_n222), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n204), .A2(new_n212), .A3(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n214), .A2(KEYINPUT10), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  AOI21_X1  g046(.A(G131), .B1(new_n231), .B2(G137), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT11), .A3(G134), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n232), .A2(new_n233), .A3(new_n238), .A4(new_n235), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n232), .B(new_n235), .C1(G134), .C2(new_n234), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n237), .A2(new_n239), .B1(G131), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT10), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n213), .B2(new_n225), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n221), .A2(new_n222), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n250), .A3(KEYINPUT65), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n207), .A2(new_n210), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G101), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n211), .B1(new_n207), .B2(new_n210), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n252), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n229), .A2(new_n241), .A3(new_n243), .A4(new_n258), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n204), .A2(new_n212), .A3(new_n227), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n227), .B1(new_n204), .B2(new_n212), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n225), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n226), .A2(new_n204), .A3(new_n212), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n237), .A2(new_n239), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n240), .A2(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT12), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT12), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n269), .B(new_n241), .C1(new_n262), .C2(new_n263), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n259), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n258), .A2(new_n243), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n224), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n260), .A2(new_n261), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n267), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT81), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n277), .B(new_n267), .C1(new_n272), .C2(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n259), .A2(new_n195), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n196), .A2(new_n271), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n190), .B1(new_n282), .B2(G469), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT74), .B(G902), .Z(new_n284));
  AOI21_X1  g098(.A(new_n195), .B1(new_n279), .B2(new_n259), .ZN(new_n285));
  INV_X1    g099(.A(new_n268), .ZN(new_n286));
  INV_X1    g100(.A(new_n270), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n280), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n188), .B(new_n284), .C1(new_n285), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT9), .B(G234), .ZN(new_n291));
  OAI21_X1  g105(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n187), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G119), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G116), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT5), .ZN(new_n301));
  OAI21_X1  g115(.A(G113), .B1(new_n298), .B2(KEYINPUT5), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n300), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT2), .B(G113), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n301), .A2(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n214), .A2(new_n306), .A3(new_n228), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT85), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n213), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n213), .B2(new_n305), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n214), .A2(new_n313), .A3(new_n306), .A4(new_n228), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n308), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G110), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT8), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n226), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n247), .A2(new_n251), .A3(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G224), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT7), .B1(new_n323), .B2(G953), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n324), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n303), .B(new_n304), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n255), .B(new_n329), .C1(new_n256), .C2(new_n257), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n307), .A2(new_n330), .A3(new_n316), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(G902), .B1(new_n318), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n323), .A2(G953), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT84), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n322), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n307), .A2(new_n330), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n316), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(KEYINPUT6), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n331), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT6), .B1(new_n337), .B2(new_n339), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n336), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G210), .B1(G237), .B2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n333), .A2(new_n343), .A3(new_n345), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n296), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n290), .A2(new_n187), .A3(new_n292), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n294), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT20), .ZN(new_n352));
  XOR2_X1   g166(.A(G113), .B(G122), .Z(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT91), .B(G104), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(G140), .B1(KEYINPUT75), .B2(G125), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT16), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n360));
  INV_X1    g174(.A(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G125), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n360), .B1(new_n362), .B2(KEYINPUT16), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT16), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(new_n361), .A3(KEYINPUT76), .A4(G125), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n359), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G146), .ZN(new_n368));
  INV_X1    g182(.A(G237), .ZN(new_n369));
  INV_X1    g183(.A(G953), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G214), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT87), .A3(new_n215), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n215), .A2(KEYINPUT87), .ZN(new_n373));
  NOR2_X1   g187(.A1(G237), .A2(G953), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(G214), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G131), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT17), .ZN(new_n378));
  INV_X1    g192(.A(G131), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n372), .A2(new_n379), .A3(new_n375), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n366), .A2(new_n218), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(KEYINPUT17), .A3(G131), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n368), .A2(new_n381), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(KEYINPUT18), .A2(G131), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n372), .A2(new_n385), .A3(new_n375), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT75), .A2(G125), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n361), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(G146), .A3(new_n356), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n319), .A2(G140), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n362), .A2(new_n392), .A3(new_n218), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(new_n391), .B2(new_n393), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n387), .B(new_n388), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n388), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n385), .B1(new_n372), .B2(new_n375), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n391), .A2(new_n393), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT88), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n395), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT89), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n355), .B(new_n384), .C1(new_n400), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(new_n399), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n403), .A2(new_n406), .A3(KEYINPUT89), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n390), .A2(KEYINPUT19), .A3(new_n356), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT19), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n362), .A2(new_n392), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n413), .A3(new_n218), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT90), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n367), .A2(G146), .B1(new_n377), .B2(new_n380), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n409), .A2(new_n410), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n408), .B1(new_n417), .B2(new_n355), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n352), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n352), .A3(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n408), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n409), .A2(new_n410), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n355), .B1(new_n425), .B2(new_n384), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n189), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G475), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n370), .B(new_n284), .C1(G234), .C2(G237), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(G898), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n370), .A2(G952), .ZN(new_n433));
  INV_X1    g247(.A(G234), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(new_n369), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n215), .A2(G128), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n223), .A2(G143), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n231), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n299), .A2(KEYINPUT14), .A3(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(G116), .B(G122), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(G107), .B(new_n441), .C1(new_n443), .C2(KEYINPUT14), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n440), .B(new_n444), .C1(G107), .C2(new_n443), .ZN(new_n445));
  INV_X1    g259(.A(new_n437), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n438), .B1(new_n446), .B2(KEYINPUT13), .ZN(new_n448));
  OAI21_X1  g262(.A(G134), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n439), .A2(new_n231), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n442), .B(new_n202), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G217), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n291), .A2(new_n453), .A3(G953), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n445), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(new_n445), .B2(new_n452), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n284), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT92), .ZN(new_n458));
  INV_X1    g272(.A(G478), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(KEYINPUT15), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT92), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n461), .B(new_n284), .C1(new_n455), .C2(new_n456), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n457), .A2(new_n460), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n429), .A2(new_n436), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n351), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n370), .A2(G221), .A3(G234), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT77), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT22), .B(G137), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT23), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n297), .B2(G128), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n474), .B(new_n475), .C1(G119), .C2(new_n223), .ZN(new_n476));
  XNOR2_X1  g290(.A(G119), .B(G128), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT24), .B(G110), .Z(new_n478));
  OAI22_X1  g292(.A1(new_n476), .A2(G110), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n368), .A2(new_n479), .A3(new_n393), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(G110), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n477), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n368), .B2(new_n382), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n472), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n368), .A2(new_n382), .ZN(new_n486));
  INV_X1    g300(.A(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n368), .A2(new_n479), .A3(new_n393), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n471), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n490), .A3(new_n284), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n453), .B1(new_n284), .B2(G234), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(G902), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n267), .A2(new_n252), .ZN(new_n500));
  INV_X1    g314(.A(new_n329), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n231), .A2(G137), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n234), .A2(G134), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n220), .A2(new_n224), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n265), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(KEYINPUT67), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT67), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n265), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n500), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(KEYINPUT68), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n252), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n506), .B(KEYINPUT30), .C1(new_n519), .C2(new_n241), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n500), .A2(KEYINPUT69), .A3(KEYINPUT30), .A4(new_n506), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n501), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n508), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n374), .A2(G210), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT27), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT26), .B(G101), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n499), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n508), .A2(KEYINPUT28), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n508), .A2(KEYINPUT28), .B1(new_n329), .B2(new_n512), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT29), .B1(new_n533), .B2(new_n529), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n512), .A2(KEYINPUT68), .A3(new_n513), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT68), .B1(new_n512), .B2(new_n513), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n524), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n507), .ZN(new_n538));
  INV_X1    g352(.A(new_n529), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(KEYINPUT72), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n530), .A2(new_n534), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n284), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n508), .A2(KEYINPUT28), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n507), .A2(KEYINPUT73), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n500), .A2(new_n545), .A3(new_n501), .A4(new_n506), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n500), .A2(new_n506), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n544), .B(new_n546), .C1(new_n501), .C2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n543), .B1(new_n549), .B2(KEYINPUT28), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n529), .A2(KEYINPUT29), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n542), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n541), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT70), .B1(new_n508), .B2(new_n539), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT70), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n507), .A2(new_n556), .A3(new_n529), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n537), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT31), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n537), .A2(new_n558), .A3(KEYINPUT31), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n554), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(G472), .A2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n553), .A2(G472), .B1(new_n566), .B2(KEYINPUT32), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n563), .B2(new_n565), .ZN(new_n569));
  INV_X1    g383(.A(new_n554), .ZN(new_n570));
  INV_X1    g384(.A(new_n562), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT31), .B1(new_n537), .B2(new_n558), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT71), .A3(new_n564), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n498), .B1(new_n567), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n467), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G101), .ZN(G3));
  NAND2_X1  g393(.A1(new_n573), .A2(new_n284), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n569), .A3(new_n574), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n292), .ZN(new_n584));
  AOI211_X1 g398(.A(KEYINPUT82), .B(new_n584), .C1(new_n283), .C2(new_n289), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n293), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n498), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT93), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n349), .A2(new_n436), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n455), .A2(new_n456), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT33), .Z(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(G478), .A3(new_n284), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n458), .A2(new_n459), .A3(new_n462), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n423), .A2(new_n428), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  NOR3_X1   g415(.A1(new_n590), .A2(new_n596), .A3(new_n465), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n589), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G107), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT94), .B(KEYINPUT35), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n471), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT95), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n488), .A2(new_n489), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n496), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n495), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n466), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n616), .A2(new_n581), .A3(new_n569), .A4(new_n574), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n351), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT37), .B(G110), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G12));
  INV_X1    g434(.A(new_n435), .ZN(new_n621));
  INV_X1    g435(.A(G900), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n430), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n418), .A2(new_n352), .A3(new_n419), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n428), .B(new_n624), .C1(new_n625), .C2(new_n420), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n465), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n349), .A2(new_n627), .A3(new_n614), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n293), .A2(new_n585), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n553), .A2(G472), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n566), .A2(KEYINPUT32), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n576), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n629), .B2(new_n632), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n223), .ZN(G30));
  XOR2_X1   g451(.A(new_n623), .B(KEYINPUT39), .Z(new_n638));
  NAND2_X1  g452(.A1(new_n586), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n639), .A2(KEYINPUT40), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(KEYINPUT40), .ZN(new_n641));
  INV_X1    g455(.A(new_n549), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n559), .B1(new_n529), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n189), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n566), .A2(KEYINPUT32), .B1(G472), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n576), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n347), .A2(new_n348), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT97), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT99), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n647), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n463), .A2(new_n464), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n596), .A2(new_n652), .ZN(new_n653));
  NOR4_X1   g467(.A1(new_n651), .A2(new_n296), .A3(new_n614), .A4(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n640), .A2(new_n641), .A3(new_n646), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT100), .B(G143), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G45));
  INV_X1    g471(.A(new_n349), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n595), .A2(new_n596), .A3(new_n624), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n658), .A2(new_n659), .A3(new_n615), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n632), .A2(new_n586), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  NOR2_X1   g476(.A1(new_n188), .A2(KEYINPUT101), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n285), .A2(new_n288), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n542), .ZN(new_n665));
  OAI221_X1 g479(.A(new_n284), .B1(KEYINPUT101), .B2(new_n188), .C1(new_n285), .C2(new_n288), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n292), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n577), .A2(new_n598), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT41), .B(G113), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G15));
  NAND4_X1  g485(.A1(new_n632), .A2(new_n668), .A3(new_n587), .A4(new_n602), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n577), .A2(KEYINPUT102), .A3(new_n602), .A4(new_n668), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  AND2_X1   g491(.A1(new_n665), .A2(new_n666), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n349), .A3(new_n679), .A4(new_n292), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT103), .B1(new_n667), .B2(new_n658), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n632), .A3(new_n616), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT104), .B(G119), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G21));
  NAND4_X1  g499(.A1(new_n665), .A2(new_n666), .A3(new_n292), .A4(new_n436), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n349), .A2(new_n596), .A3(new_n652), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n550), .A2(KEYINPUT105), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n539), .B1(new_n550), .B2(KEYINPUT105), .ZN(new_n690));
  OAI22_X1  g504(.A1(new_n689), .A2(new_n690), .B1(new_n571), .B2(new_n572), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n580), .A2(G472), .B1(new_n691), .B2(new_n564), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n587), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  INV_X1    g508(.A(new_n692), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n695), .A2(new_n615), .A3(new_n659), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n682), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  NAND2_X1  g512(.A1(new_n573), .A2(new_n564), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n575), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT32), .B1(new_n573), .B2(new_n564), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT106), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n701), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n631), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n705), .A3(new_n630), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n647), .A2(new_n296), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n292), .A3(new_n290), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n659), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n709), .A3(new_n587), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n711));
  INV_X1    g525(.A(new_n708), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n659), .A2(KEYINPUT42), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n577), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT107), .B(G131), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G33));
  NAND3_X1  g531(.A1(new_n577), .A2(new_n627), .A3(new_n712), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G134), .ZN(G36));
  OR2_X1    g533(.A1(new_n282), .A2(KEYINPUT45), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n282), .A2(KEYINPUT45), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(G469), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n190), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(KEYINPUT46), .A3(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n723), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n725), .A2(new_n289), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n730), .A2(new_n292), .A3(new_n638), .ZN(new_n731));
  INV_X1    g545(.A(new_n707), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT43), .B1(new_n429), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n429), .A2(new_n595), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n582), .A3(new_n614), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n732), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n731), .B(new_n739), .C1(new_n738), .C2(new_n737), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G137), .ZN(G39));
  NOR4_X1   g555(.A1(new_n632), .A2(new_n587), .A3(new_n659), .A4(new_n732), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n730), .A2(KEYINPUT47), .A3(new_n292), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT47), .B1(new_n730), .B2(new_n292), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G140), .ZN(G42));
  XNOR2_X1  g560(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n736), .A2(new_n587), .A3(new_n621), .A4(new_n692), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n732), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT115), .Z(new_n750));
  NOR2_X1   g564(.A1(new_n743), .A2(new_n744), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n665), .A2(new_n666), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n292), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT116), .ZN(new_n755));
  INV_X1    g569(.A(new_n646), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n732), .A2(new_n667), .A3(new_n435), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n587), .A3(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n596), .A3(new_n595), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n695), .A2(new_n615), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n736), .A2(new_n757), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n651), .A2(new_n296), .A3(new_n668), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n748), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n766), .B2(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n755), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n754), .A2(KEYINPUT116), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n747), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(KEYINPUT51), .A3(new_n754), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n706), .A2(new_n587), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n761), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT48), .Z(new_n776));
  INV_X1    g590(.A(new_n682), .ZN(new_n777));
  OAI221_X1 g591(.A(new_n433), .B1(new_n758), .B2(new_n597), .C1(new_n777), .C2(new_n748), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n772), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n697), .B1(new_n634), .B2(new_n635), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n697), .B(KEYINPUT112), .C1(new_n634), .C2(new_n635), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n614), .A2(new_n623), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n292), .A3(new_n290), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n687), .B1(new_n786), .B2(KEYINPUT113), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n646), .C1(KEYINPUT113), .C2(new_n786), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n661), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n783), .A2(new_n784), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n790), .B1(new_n781), .B2(new_n789), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n693), .B1(new_n617), .B2(new_n351), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n577), .B2(new_n467), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n652), .B(KEYINPUT111), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(new_n596), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n590), .B1(new_n798), .B2(new_n597), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n583), .A3(new_n586), .A4(new_n587), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n683), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n796), .A2(new_n676), .A3(new_n669), .A4(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n632), .A2(new_n586), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n797), .A2(new_n614), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n732), .A2(new_n804), .A3(new_n626), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n803), .A2(new_n805), .B1(new_n696), .B2(new_n712), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n711), .A2(new_n806), .A3(new_n714), .A4(new_n718), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n794), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n635), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n812), .A2(new_n813), .B1(new_n682), .B2(new_n696), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT52), .A3(new_n661), .A4(new_n788), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n793), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n808), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n811), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n810), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n794), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n780), .A2(new_n824), .B1(G952), .B2(G953), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n735), .A2(new_n498), .A3(new_n296), .A4(new_n584), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT110), .Z(new_n827));
  OAI21_X1  g641(.A(new_n651), .B1(KEYINPUT49), .B2(new_n752), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(KEYINPUT49), .B2(new_n752), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n756), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n825), .A2(new_n830), .ZN(G75));
  NOR2_X1   g645(.A1(new_n370), .A2(G952), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n794), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n816), .B2(new_n808), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n284), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n837), .B2(new_n346), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n341), .A2(new_n342), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(new_n336), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT55), .Z(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n833), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n838), .B2(new_n842), .ZN(G51));
  OAI21_X1  g658(.A(KEYINPUT54), .B1(new_n834), .B2(new_n835), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n823), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n190), .B(KEYINPUT57), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n664), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n722), .B(KEYINPUT118), .Z(new_n849));
  OAI211_X1 g663(.A(new_n542), .B(new_n849), .C1(new_n834), .C2(new_n835), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n820), .A2(new_n822), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT119), .A3(new_n542), .A4(new_n849), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n833), .B1(new_n848), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT120), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n833), .C1(new_n848), .C2(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(G54));
  NAND3_X1  g674(.A1(new_n837), .A2(KEYINPUT58), .A3(G475), .ZN(new_n861));
  INV_X1    g675(.A(new_n418), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(new_n832), .ZN(G60));
  NAND2_X1  g679(.A1(G478), .A2(G902), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT59), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n592), .B1(new_n824), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n846), .A2(new_n592), .A3(new_n867), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n868), .A2(new_n832), .A3(new_n869), .ZN(G63));
  XNOR2_X1  g684(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n871));
  NAND2_X1  g685(.A1(G217), .A2(G902), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n836), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n611), .A2(new_n612), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n485), .A2(new_n490), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n836), .B2(new_n873), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n833), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(G66));
  OAI21_X1  g695(.A(G953), .B1(new_n431), .B2(new_n323), .ZN(new_n882));
  INV_X1    g696(.A(new_n802), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n882), .B1(new_n883), .B2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n839), .B1(G898), .B2(new_n370), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT123), .Z(new_n886));
  XNOR2_X1  g700(.A(new_n884), .B(new_n886), .ZN(G69));
  NAND2_X1  g701(.A1(new_n622), .A2(G953), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT125), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n687), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n731), .A2(new_n891), .A3(new_n774), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n740), .A2(new_n745), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n783), .A2(new_n784), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n715), .A2(new_n718), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n661), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n890), .B1(new_n896), .B2(new_n370), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n522), .A2(new_n523), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n518), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n411), .A2(new_n413), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT124), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n894), .A2(new_n655), .A3(new_n661), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n904), .A2(KEYINPUT62), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n732), .B1(new_n798), .B2(new_n597), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n577), .A2(new_n586), .A3(new_n638), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n740), .A2(new_n745), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n904), .B2(KEYINPUT62), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n901), .B1(new_n910), .B2(new_n370), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(G953), .B1(new_n193), .B2(new_n622), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(G72));
  NAND2_X1  g728(.A1(G472), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT63), .Z(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n910), .B2(new_n802), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n538), .B(KEYINPUT126), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n529), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT127), .B1(new_n530), .B2(new_n540), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n537), .B2(new_n558), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n530), .A2(KEYINPUT127), .A3(new_n540), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n818), .A2(new_n916), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n916), .B1(new_n896), .B2(new_n802), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n918), .A2(new_n529), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n832), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n919), .A2(new_n924), .A3(new_n927), .ZN(G57));
endmodule


