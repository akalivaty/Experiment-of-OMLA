//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n187));
  INV_X1    g001(.A(G469), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G227), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT3), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT4), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n198), .B2(new_n200), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n198), .A2(new_n200), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G101), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT0), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(new_n210), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n213), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n207), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n208), .A2(new_n221), .A3(G128), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n214), .A2(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n212), .A2(G146), .ZN(new_n225));
  AOI21_X1  g039(.A(G128), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n221), .A2(new_n214), .A3(G143), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n229), .B(KEYINPUT64), .C1(new_n208), .C2(G128), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n222), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT77), .B1(new_n196), .B2(G104), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n194), .A3(G107), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n196), .A2(G104), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n201), .A3(KEYINPUT10), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n204), .A2(new_n220), .B1(new_n231), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT78), .B1(new_n226), .B2(new_n227), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n208), .A2(new_n221), .A3(G128), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT78), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n229), .B(new_n244), .C1(new_n208), .C2(G128), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n237), .A2(new_n201), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n239), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT11), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G137), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n252), .A2(new_n254), .A3(new_n258), .A4(new_n255), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(KEYINPUT80), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n192), .B1(new_n249), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n239), .B2(new_n248), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT81), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n246), .A2(new_n247), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n240), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n210), .B1(new_n213), .B2(new_n215), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT64), .B1(new_n268), .B2(new_n229), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n226), .A2(new_n223), .A3(new_n227), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n243), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n247), .ZN(new_n272));
  INV_X1    g086(.A(new_n203), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n219), .A3(new_n207), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n267), .A2(new_n261), .A3(new_n272), .A4(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n260), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n228), .A2(new_n230), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n237), .A2(new_n201), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n243), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n277), .B1(new_n266), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT12), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT12), .ZN(new_n283));
  AOI211_X1 g097(.A(new_n283), .B(new_n277), .C1(new_n266), .C2(new_n280), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n265), .B(new_n276), .C1(new_n282), .C2(new_n284), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n192), .B(KEYINPUT76), .Z(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n266), .A2(new_n280), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n260), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n283), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n281), .A2(KEYINPUT12), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n265), .B1(new_n292), .B2(new_n276), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n264), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n188), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n298));
  INV_X1    g112(.A(new_n192), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n276), .B(new_n299), .C1(new_n282), .C2(new_n284), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n276), .A2(new_n263), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n300), .A2(new_n301), .B1(new_n192), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n292), .A2(new_n262), .A3(KEYINPUT82), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n305), .B2(new_n188), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n282), .A2(new_n284), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n276), .A2(new_n299), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n301), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n302), .A2(new_n192), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n311), .A2(new_n298), .A3(new_n188), .A4(new_n295), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n297), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT2), .A2(G113), .ZN(new_n320));
  NAND2_X1  g134(.A1(KEYINPUT2), .A2(G113), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G116), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT66), .B1(new_n326), .B2(G119), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G116), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(G119), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n327), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n327), .A2(new_n330), .A3(new_n331), .ZN(new_n333));
  INV_X1    g147(.A(new_n324), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n336), .B2(new_n320), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n332), .A2(new_n337), .B1(new_n203), .B2(new_n206), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n274), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n327), .A2(new_n330), .A3(KEYINPUT5), .A4(new_n331), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n326), .A2(KEYINPUT5), .A3(G119), .ZN(new_n342));
  INV_X1    g156(.A(G113), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n247), .A2(new_n340), .A3(new_n332), .A4(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n332), .A2(new_n345), .A3(new_n201), .A4(new_n237), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT84), .ZN(new_n348));
  XNOR2_X1  g162(.A(G110), .B(G122), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n339), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n338), .A2(new_n274), .B1(new_n347), .B2(KEYINPUT84), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT86), .A3(new_n349), .A4(new_n346), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n346), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n349), .B(KEYINPUT85), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n356), .A3(new_n358), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n219), .A2(G125), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n231), .B2(G125), .ZN(new_n363));
  INV_X1    g177(.A(G224), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G953), .ZN(new_n365));
  XOR2_X1   g179(.A(new_n363), .B(new_n365), .Z(new_n366));
  NAND3_X1  g180(.A1(new_n360), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT7), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n362), .B(new_n369), .C1(new_n231), .C2(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n332), .A2(new_n345), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n279), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n347), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n349), .B(KEYINPUT8), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n373), .A2(KEYINPUT87), .A3(new_n378), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n355), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n367), .A2(new_n295), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G210), .B1(G237), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n367), .A2(new_n295), .A3(new_n383), .A4(new_n385), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n319), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n326), .A2(G122), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n196), .B1(new_n390), .B2(KEYINPUT14), .ZN(new_n391));
  XNOR2_X1  g205(.A(G116), .B(G122), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n391), .B(new_n392), .Z(new_n393));
  OAI21_X1  g207(.A(KEYINPUT92), .B1(new_n210), .B2(G143), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT92), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n212), .A3(G128), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n210), .A2(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n251), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT13), .B1(new_n394), .B2(new_n396), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT93), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT13), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT94), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT94), .A4(KEYINPUT13), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n406), .A2(new_n407), .A3(new_n398), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n251), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n392), .B(new_n196), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n397), .A2(new_n251), .A3(new_n398), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT95), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n404), .A2(new_n405), .B1(new_n210), .B2(G143), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n402), .A2(KEYINPUT93), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT93), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n416), .B(KEYINPUT13), .C1(new_n394), .C2(new_n396), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n414), .B(new_n407), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G134), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n420));
  INV_X1    g234(.A(new_n412), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n401), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G217), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n315), .A2(new_n424), .A3(G953), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n401), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n420), .B1(new_n419), .B2(new_n421), .ZN(new_n428));
  AOI211_X1 g242(.A(KEYINPUT95), .B(new_n412), .C1(new_n418), .C2(G134), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n427), .B(new_n425), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n295), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT96), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n437));
  INV_X1    g251(.A(new_n425), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n439), .B2(new_n430), .ZN(new_n440));
  INV_X1    g254(.A(new_n435), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT96), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n295), .B(new_n441), .C1(new_n426), .C2(new_n431), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT97), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(KEYINPUT97), .A3(new_n441), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n436), .A2(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(G234), .A2(G237), .ZN(new_n448));
  INV_X1    g262(.A(G953), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n448), .A2(G952), .A3(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n448), .A2(G902), .A3(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(G898), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G237), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n455), .A2(new_n449), .A3(G214), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(G143), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT18), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT88), .B(G143), .ZN(new_n460));
  OAI221_X1 g274(.A(new_n458), .B1(new_n459), .B2(new_n258), .C1(new_n456), .C2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT90), .ZN(new_n462));
  XNOR2_X1  g276(.A(G125), .B(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n214), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G140), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G125), .ZN(new_n467));
  INV_X1    g281(.A(G125), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G140), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT89), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n465), .B1(new_n471), .B2(G146), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n212), .A2(KEYINPUT88), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n456), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n460), .A2(new_n456), .ZN(new_n475));
  OAI21_X1  g289(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n472), .B1(KEYINPUT18), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n462), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n474), .A2(new_n475), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n258), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n476), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n463), .A2(KEYINPUT16), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n467), .A2(KEYINPUT16), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(new_n214), .ZN(new_n487));
  AOI21_X1  g301(.A(G146), .B1(new_n484), .B2(new_n485), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n483), .B(new_n489), .C1(new_n482), .C2(new_n476), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n479), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G113), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n194), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n479), .A2(new_n490), .A3(new_n493), .ZN(new_n496));
  AOI21_X1  g310(.A(G902), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G475), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n471), .A2(KEYINPUT91), .A3(KEYINPUT19), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n470), .B2(KEYINPUT19), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n471), .B2(KEYINPUT19), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n214), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n487), .B1(new_n481), .B2(new_n476), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n462), .A2(new_n478), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n496), .B1(new_n507), .B2(new_n493), .ZN(new_n508));
  NOR2_X1   g322(.A1(G475), .A2(G902), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n500), .A3(new_n509), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n499), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n389), .A2(new_n447), .A3(new_n454), .A4(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n187), .B1(new_n317), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n383), .A2(new_n295), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n385), .B1(new_n516), .B2(new_n367), .ZN(new_n517));
  INV_X1    g331(.A(new_n388), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n454), .B(new_n318), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n436), .A2(new_n442), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n445), .A2(new_n446), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n311), .A2(new_n188), .A3(new_n295), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT83), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n296), .B1(new_n525), .B2(new_n312), .ZN(new_n526));
  INV_X1    g340(.A(new_n316), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT98), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT32), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n332), .A2(new_n337), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT70), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n260), .A2(new_n219), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n332), .A2(new_n337), .A3(KEYINPUT70), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n251), .A2(G137), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n253), .A2(G134), .ZN(new_n539));
  OAI21_X1  g353(.A(G131), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n259), .A2(new_n540), .A3(KEYINPUT67), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT67), .B1(new_n259), .B2(new_n540), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n271), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT28), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(KEYINPUT68), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n278), .B2(new_n243), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n542), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n537), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n259), .A2(new_n257), .B1(new_n211), .B2(new_n218), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n259), .A2(new_n540), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n271), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n531), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n534), .B1(new_n231), .B2(new_n554), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(KEYINPUT72), .A3(new_n531), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n551), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n546), .B1(new_n561), .B2(KEYINPUT28), .ZN(new_n562));
  XOR2_X1   g376(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n563));
  NAND3_X1  g377(.A1(new_n455), .A2(new_n449), .A3(G210), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT26), .B(G101), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n551), .A2(new_n567), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n549), .B1(new_n548), .B2(new_n542), .ZN(new_n571));
  NOR4_X1   g385(.A1(new_n231), .A2(new_n541), .A3(KEYINPUT68), .A4(new_n543), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n534), .A2(KEYINPUT30), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT30), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n557), .B1(new_n559), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT69), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT69), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n547), .A2(KEYINPUT30), .A3(new_n534), .A4(new_n550), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n576), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n570), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT31), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT69), .B1(new_n574), .B2(new_n577), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n579), .A3(new_n576), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT31), .A3(new_n570), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n568), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(G472), .A2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n530), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT31), .B1(new_n587), .B2(new_n570), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n583), .B(new_n569), .C1(new_n585), .C2(new_n586), .ZN(new_n594));
  OAI22_X1  g408(.A1(new_n593), .A2(new_n594), .B1(new_n567), .B2(new_n562), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT32), .A3(new_n590), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT73), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT29), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n558), .A2(new_n560), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n571), .A2(new_n572), .A3(new_n536), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT28), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n546), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n567), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n585), .B2(new_n586), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n598), .B(new_n603), .C1(new_n604), .C2(new_n567), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n571), .A2(new_n572), .A3(new_n553), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n533), .A2(new_n535), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n551), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n546), .B1(new_n609), .B2(KEYINPUT28), .ZN(new_n610));
  INV_X1    g424(.A(new_n567), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n598), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n597), .B1(new_n614), .B2(G472), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  AOI211_X1 g430(.A(KEYINPUT73), .B(new_n616), .C1(new_n605), .C2(new_n613), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n592), .B(new_n596), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT22), .B(G137), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n449), .A2(G221), .A3(G234), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n210), .A2(G119), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n329), .A2(G128), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT74), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT24), .B(G110), .Z(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT75), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n329), .A2(G128), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n624), .B(new_n630), .C1(new_n631), .C2(KEYINPUT23), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G110), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n489), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n626), .A2(new_n627), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n633), .A2(new_n634), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n487), .B(new_n465), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n622), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n640), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n629), .A2(new_n636), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n621), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n641), .A2(new_n295), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT25), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n641), .A2(KEYINPUT25), .A3(new_n644), .A4(new_n295), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n424), .B1(G234), .B2(new_n295), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(G902), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n641), .A2(new_n644), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n515), .A2(new_n529), .A3(new_n618), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  INV_X1    g470(.A(new_n654), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n317), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n508), .A2(new_n500), .A3(new_n509), .ZN(new_n659));
  OAI22_X1  g473(.A1(new_n659), .A2(new_n510), .B1(new_n498), .B2(new_n497), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n434), .A2(G902), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n438), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n423), .B2(KEYINPUT99), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n430), .A2(new_n663), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  INV_X1    g481(.A(new_n664), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n437), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT33), .ZN(new_n671));
  OR3_X1    g485(.A1(new_n426), .A2(new_n431), .A3(KEYINPUT33), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n662), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n440), .A2(G478), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n660), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n519), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n595), .A2(new_n590), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n616), .B1(new_n595), .B2(new_n295), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n658), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT34), .B(G104), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G6));
  NAND2_X1  g497(.A1(new_n520), .A2(new_n521), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n513), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n519), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n658), .A2(new_n680), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  NAND2_X1  g503(.A1(new_n642), .A2(new_n643), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n622), .A2(KEYINPUT36), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT101), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n690), .B(new_n692), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n649), .A2(new_n650), .B1(new_n652), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n515), .A2(new_n529), .A3(new_n680), .A4(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT37), .B(G110), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n451), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n450), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n684), .A2(new_n513), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n387), .A2(new_n388), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n318), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n694), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n618), .A2(new_n704), .A3(new_n528), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  INV_X1    g523(.A(new_n604), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n567), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n295), .B1(new_n609), .B2(new_n567), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n592), .A2(new_n596), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n715), .B(KEYINPUT102), .Z(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n660), .A2(new_n318), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n447), .A2(new_n695), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n517), .A2(new_n518), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT38), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n720), .A2(KEYINPUT38), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n702), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n528), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n723), .B1(KEYINPUT40), .B2(new_n726), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n726), .A2(KEYINPUT40), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n717), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  OAI211_X1 g544(.A(new_n660), .B(new_n702), .C1(new_n673), .C2(new_n674), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n526), .A3(new_n527), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n618), .A3(new_n707), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  NAND2_X1  g548(.A1(new_n311), .A2(new_n295), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n316), .B(new_n736), .C1(new_n306), .C2(new_n313), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n618), .A2(new_n738), .A3(new_n654), .A4(new_n676), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND4_X1  g555(.A1(new_n618), .A2(new_n686), .A3(new_n654), .A4(new_n738), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  NOR2_X1   g557(.A1(new_n737), .A2(new_n706), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n522), .A2(new_n453), .A3(new_n694), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n618), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT104), .B(G119), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G21));
  NAND2_X1  g562(.A1(new_n610), .A2(KEYINPUT105), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT28), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n547), .A2(new_n534), .A3(new_n550), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n607), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n751), .B1(new_n753), .B2(new_n551), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n750), .B1(new_n754), .B2(new_n546), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n749), .A2(new_n611), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n584), .A2(new_n588), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n591), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(G472), .B1(new_n589), .B2(G902), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n654), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n737), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n720), .A2(new_n447), .A3(new_n718), .A4(new_n453), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NOR3_X1   g579(.A1(new_n679), .A2(new_n758), .A3(new_n694), .ZN(new_n766));
  INV_X1    g580(.A(new_n731), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n744), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  AOI21_X1  g583(.A(new_n616), .B1(new_n605), .B2(new_n613), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n597), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n596), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n596), .A2(new_n772), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n592), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n387), .A2(new_n318), .A3(new_n388), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n526), .A2(new_n527), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n767), .A2(KEYINPUT42), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(new_n654), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n618), .A2(new_n777), .A3(new_n654), .A4(new_n767), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  AND2_X1   g598(.A1(new_n592), .A2(new_n596), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n657), .B1(new_n771), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(KEYINPUT108), .A3(new_n704), .A4(new_n777), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n618), .A2(new_n777), .A3(new_n704), .A4(new_n654), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  AOI21_X1  g606(.A(new_n694), .B1(new_n760), .B2(new_n677), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n671), .A2(new_n672), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n674), .B1(new_n794), .B2(new_n661), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT43), .B1(new_n795), .B2(new_n660), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT43), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n797), .B(new_n513), .C1(new_n673), .C2(new_n674), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n776), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n796), .A2(new_n798), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(KEYINPUT44), .A3(new_n793), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(KEYINPUT110), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n525), .A2(new_n312), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n188), .A2(new_n295), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT45), .B(new_n264), .C1(new_n287), .C2(new_n293), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT109), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n188), .B1(new_n294), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n806), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n805), .B1(new_n811), .B2(KEYINPUT46), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT46), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n813), .B(new_n806), .C1(new_n808), .C2(new_n810), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n316), .B(new_n725), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n804), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n801), .A2(new_n803), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G137), .ZN(G39));
  OAI21_X1  g636(.A(new_n316), .B1(new_n812), .B2(new_n814), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(KEYINPUT47), .B(new_n316), .C1(new_n812), .C2(new_n814), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n654), .A2(new_n776), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n771), .A2(new_n785), .A3(new_n767), .A4(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT111), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(new_n833), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G140), .ZN(G42));
  NAND2_X1  g650(.A1(new_n805), .A2(new_n736), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n839));
  OAI221_X1 g653(.A(new_n513), .B1(new_n674), .B2(new_n673), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n722), .A2(new_n721), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n657), .A2(new_n527), .A3(new_n319), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n716), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n802), .A2(new_n450), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n319), .A3(new_n842), .A4(new_n762), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT50), .Z(new_n847));
  INV_X1    g661(.A(new_n776), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n761), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n837), .A2(new_n316), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n850), .B1(new_n827), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n845), .A2(new_n738), .A3(new_n766), .A4(new_n848), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n654), .A2(new_n848), .A3(new_n450), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n717), .A2(new_n737), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n513), .A3(new_n795), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n847), .A2(new_n852), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n845), .A2(new_n738), .A3(new_n848), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n775), .A2(new_n654), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT48), .Z(new_n864));
  NAND3_X1  g678(.A1(new_n845), .A2(new_n389), .A3(new_n762), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT115), .Z(new_n866));
  INV_X1    g680(.A(G952), .ZN(new_n867));
  INV_X1    g681(.A(new_n675), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n867), .B(G953), .C1(new_n855), .C2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n860), .A2(new_n864), .A3(new_n866), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n720), .A2(new_n447), .A3(new_n718), .ZN(new_n872));
  INV_X1    g686(.A(new_n702), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n695), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n715), .A3(new_n528), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n708), .A2(new_n733), .A3(new_n768), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n317), .A2(new_n703), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n618), .B(new_n707), .C1(new_n879), .C2(new_n732), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n768), .A4(new_n875), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n790), .A2(new_n787), .B1(new_n779), .B2(new_n782), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n764), .A2(new_n739), .A3(new_n742), .A4(new_n746), .ZN(new_n884));
  INV_X1    g698(.A(new_n777), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n684), .A2(new_n694), .A3(new_n660), .A4(new_n873), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n618), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n766), .A2(new_n767), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n882), .A2(new_n883), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n655), .A2(new_n681), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT113), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n655), .A2(KEYINPUT113), .A3(new_n681), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n686), .A2(KEYINPUT114), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n685), .B2(new_n519), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n658), .A3(new_n680), .A4(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n894), .A2(new_n696), .A3(new_n895), .A4(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n871), .B1(new_n891), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n791), .A2(new_n783), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n618), .A2(new_n745), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n903), .A2(new_n744), .B1(new_n762), .B2(new_n763), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n887), .A2(new_n888), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n777), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n904), .A2(new_n906), .A3(new_n739), .A4(new_n742), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n655), .A2(KEYINPUT113), .A3(new_n681), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT113), .B1(new_n655), .B2(new_n681), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n696), .A2(new_n899), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n908), .A2(new_n912), .A3(KEYINPUT53), .A4(new_n882), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n901), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n901), .A2(new_n913), .A3(KEYINPUT54), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n859), .B(new_n870), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(G952), .A2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n844), .B1(new_n918), .B2(new_n919), .ZN(G75));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n295), .B1(new_n901), .B2(new_n913), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(KEYINPUT116), .A3(G210), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n360), .A2(new_n361), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n366), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT55), .Z(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(KEYINPUT56), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT116), .B1(new_n922), .B2(G210), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n449), .A2(G952), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT56), .B1(new_n922), .B2(G210), .ZN(new_n933));
  INV_X1    g747(.A(new_n926), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n921), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n933), .A2(new_n934), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n914), .A2(G210), .A3(G902), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT116), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n923), .A3(new_n927), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n937), .A2(new_n941), .A3(KEYINPUT117), .A4(new_n932), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n936), .A2(new_n942), .ZN(G51));
  XNOR2_X1  g757(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n806), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n916), .A2(new_n917), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n311), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n922), .A2(new_n808), .A3(new_n810), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n931), .B1(new_n947), .B2(new_n948), .ZN(G54));
  AND2_X1   g763(.A1(KEYINPUT58), .A2(G475), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n922), .A2(new_n508), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n508), .B1(new_n922), .B2(new_n950), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n931), .ZN(G60));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT59), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n916), .A2(new_n917), .A3(new_n955), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n794), .B(KEYINPUT119), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n957), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n916), .A2(new_n917), .A3(new_n955), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n932), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT120), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT120), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n958), .A2(new_n963), .A3(new_n932), .A4(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n914), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n641), .A2(new_n644), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n931), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n693), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n968), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G66));
  OR2_X1    g788(.A1(new_n900), .A2(new_n884), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n449), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n452), .B2(new_n364), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(KEYINPUT121), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(KEYINPUT121), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n924), .B1(G898), .B2(new_n449), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT122), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n979), .B(new_n981), .ZN(G69));
  OAI21_X1  g796(.A(new_n580), .B1(KEYINPUT30), .B2(new_n556), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT123), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n501), .A2(new_n504), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(G900), .A2(G953), .ZN(new_n987));
  AOI22_X1  g801(.A1(new_n832), .A2(new_n834), .B1(new_n820), .B2(new_n817), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n708), .A2(new_n733), .A3(new_n768), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n880), .A2(new_n991), .A3(new_n768), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n816), .A2(new_n654), .A3(new_n872), .A4(new_n775), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n883), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n986), .B(new_n987), .C1(new_n996), .C2(G953), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n993), .A2(KEYINPUT62), .A3(new_n729), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT62), .B1(new_n993), .B2(new_n729), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n726), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n685), .A2(new_n675), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n786), .A2(new_n1002), .A3(new_n848), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n834), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n833), .B1(new_n827), .B2(new_n830), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n821), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(KEYINPUT125), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n993), .A2(new_n729), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT62), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n998), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT125), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1012), .A2(new_n988), .A3(new_n1013), .A4(new_n1004), .ZN(new_n1014));
  AOI21_X1  g828(.A(G953), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n997), .B1(new_n1015), .B2(new_n986), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n997), .A2(KEYINPUT126), .ZN(new_n1017));
  OAI21_X1  g831(.A(G953), .B1(new_n190), .B2(new_n699), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1016), .B(new_n1019), .ZN(G72));
  XNOR2_X1  g834(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n616), .A2(new_n295), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1021), .B(new_n1022), .Z(new_n1023));
  OAI21_X1  g837(.A(new_n1023), .B1(new_n996), .B2(new_n975), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n604), .A3(new_n611), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1023), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n710), .A2(new_n611), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1026), .B1(new_n1027), .B2(new_n582), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n931), .B1(new_n914), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1023), .B1(new_n1031), .B2(new_n975), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1030), .B1(new_n1032), .B2(new_n712), .ZN(G57));
endmodule


