

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U320 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U321 ( .A(n372), .B(n371), .ZN(n375) );
  XNOR2_X1 U322 ( .A(n370), .B(KEYINPUT90), .ZN(n371) );
  INV_X1 U323 ( .A(n482), .ZN(n401) );
  XNOR2_X1 U324 ( .A(n362), .B(n290), .ZN(n363) );
  XOR2_X1 U325 ( .A(n355), .B(n354), .Z(n563) );
  AND2_X1 U326 ( .A1(G228GAT), .A2(G233GAT), .ZN(n288) );
  AND2_X1 U327 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U328 ( .A(G218GAT), .B(G106GAT), .Z(n290) );
  INV_X1 U329 ( .A(KEYINPUT25), .ZN(n370) );
  XNOR2_X1 U330 ( .A(n356), .B(n288), .ZN(n357) );
  XNOR2_X1 U331 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n458) );
  NAND2_X1 U332 ( .A1(n401), .A2(n479), .ZN(n402) );
  XNOR2_X1 U333 ( .A(n364), .B(n363), .ZN(n368) );
  XNOR2_X1 U334 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U335 ( .A(n297), .B(n289), .ZN(n298) );
  XNOR2_X1 U336 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U337 ( .A(KEYINPUT36), .B(n542), .Z(n462) );
  XOR2_X1 U338 ( .A(KEYINPUT76), .B(n560), .Z(n542) );
  XOR2_X1 U339 ( .A(n419), .B(n418), .Z(n578) );
  XNOR2_X1 U340 ( .A(n437), .B(n436), .ZN(n496) );
  XNOR2_X1 U341 ( .A(n463), .B(G218GAT), .ZN(n464) );
  XNOR2_X1 U342 ( .A(n468), .B(G204GAT), .ZN(n469) );
  XNOR2_X1 U343 ( .A(n438), .B(G50GAT), .ZN(n439) );
  XNOR2_X1 U344 ( .A(n465), .B(n464), .ZN(G1355GAT) );
  XNOR2_X1 U345 ( .A(n470), .B(n469), .ZN(G1353GAT) );
  XNOR2_X1 U346 ( .A(n440), .B(n439), .ZN(G1331GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n292) );
  XNOR2_X1 U348 ( .A(KEYINPUT64), .B(KEYINPUT10), .ZN(n291) );
  XNOR2_X1 U349 ( .A(n292), .B(n291), .ZN(n307) );
  XOR2_X1 U350 ( .A(KEYINPUT74), .B(G218GAT), .Z(n294) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n330) );
  XOR2_X1 U353 ( .A(G50GAT), .B(G162GAT), .Z(n356) );
  XOR2_X1 U354 ( .A(n330), .B(n356), .Z(n299) );
  XOR2_X1 U355 ( .A(KEYINPUT11), .B(KEYINPUT73), .Z(n296) );
  XNOR2_X1 U356 ( .A(G134GAT), .B(KEYINPUT65), .ZN(n295) );
  XNOR2_X1 U357 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U358 ( .A(G29GAT), .B(G43GAT), .Z(n301) );
  XNOR2_X1 U359 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n406) );
  XOR2_X1 U361 ( .A(G92GAT), .B(G85GAT), .Z(n303) );
  XNOR2_X1 U362 ( .A(G99GAT), .B(G106GAT), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n303), .B(n302), .ZN(n430) );
  XNOR2_X1 U364 ( .A(n406), .B(n430), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n307), .B(n306), .ZN(n560) );
  XOR2_X1 U367 ( .A(KEYINPUT86), .B(G57GAT), .Z(n309) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n317) );
  NAND2_X1 U370 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U371 ( .A(KEYINPUT5), .B(G85GAT), .Z(n311) );
  XNOR2_X1 U372 ( .A(G148GAT), .B(G155GAT), .ZN(n310) );
  XNOR2_X1 U373 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U374 ( .A(G29GAT), .B(G162GAT), .Z(n312) );
  XNOR2_X1 U375 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U378 ( .A(n318), .B(KEYINPUT1), .Z(n322) );
  XOR2_X1 U379 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n320) );
  XNOR2_X1 U380 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n366) );
  XNOR2_X1 U382 ( .A(n366), .B(KEYINPUT6), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n327) );
  XNOR2_X1 U384 ( .A(G127GAT), .B(G134GAT), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n323), .B(KEYINPUT0), .ZN(n324) );
  XOR2_X1 U386 ( .A(n324), .B(KEYINPUT80), .Z(n326) );
  XNOR2_X1 U387 ( .A(G113GAT), .B(G120GAT), .ZN(n325) );
  XOR2_X1 U388 ( .A(n326), .B(n325), .Z(n345) );
  XOR2_X1 U389 ( .A(n327), .B(n345), .Z(n516) );
  XOR2_X1 U390 ( .A(G176GAT), .B(G64GAT), .Z(n422) );
  XOR2_X1 U391 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n329) );
  XNOR2_X1 U392 ( .A(G8GAT), .B(G92GAT), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n331) );
  XOR2_X1 U394 ( .A(n331), .B(n330), .Z(n340) );
  XOR2_X1 U395 ( .A(G204GAT), .B(G211GAT), .Z(n333) );
  XNOR2_X1 U396 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n358) );
  XOR2_X1 U398 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n335) );
  XNOR2_X1 U399 ( .A(KEYINPUT83), .B(KEYINPUT18), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U401 ( .A(n336), .B(KEYINPUT82), .Z(n338) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(G183GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n358), .B(n344), .ZN(n339) );
  XOR2_X1 U405 ( .A(n340), .B(n339), .Z(n341) );
  XNOR2_X1 U406 ( .A(n422), .B(n341), .ZN(n343) );
  NAND2_X1 U407 ( .A1(G226GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n505) );
  XOR2_X1 U409 ( .A(n345), .B(n344), .Z(n355) );
  XOR2_X1 U410 ( .A(G176GAT), .B(G71GAT), .Z(n347) );
  NAND2_X1 U411 ( .A1(G227GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U413 ( .A(n348), .B(G99GAT), .Z(n353) );
  XOR2_X1 U414 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n350) );
  XNOR2_X1 U415 ( .A(G15GAT), .B(G190GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U417 ( .A(G43GAT), .B(n351), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  NAND2_X1 U419 ( .A1(n505), .A2(n563), .ZN(n369) );
  XOR2_X1 U420 ( .A(G22GAT), .B(G155GAT), .Z(n393) );
  XOR2_X1 U421 ( .A(n359), .B(n393), .Z(n364) );
  XOR2_X1 U422 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n361) );
  XNOR2_X1 U423 ( .A(KEYINPUT23), .B(KEYINPUT84), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U425 ( .A(G78GAT), .B(KEYINPUT70), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n365), .B(G148GAT), .ZN(n431) );
  XNOR2_X1 U427 ( .A(n431), .B(n366), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n472) );
  NAND2_X1 U429 ( .A1(n369), .A2(n472), .ZN(n372) );
  INV_X1 U430 ( .A(n505), .ZN(n518) );
  XOR2_X1 U431 ( .A(n518), .B(KEYINPUT27), .Z(n379) );
  NOR2_X1 U432 ( .A1(n563), .A2(n472), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n373), .B(KEYINPUT26), .ZN(n546) );
  NAND2_X1 U434 ( .A1(n379), .A2(n546), .ZN(n374) );
  NAND2_X1 U435 ( .A1(n375), .A2(n374), .ZN(n376) );
  NAND2_X1 U436 ( .A1(n516), .A2(n376), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n377), .B(KEYINPUT91), .ZN(n383) );
  XOR2_X1 U438 ( .A(n472), .B(KEYINPUT66), .Z(n378) );
  XOR2_X1 U439 ( .A(KEYINPUT28), .B(n378), .Z(n523) );
  INV_X1 U440 ( .A(n523), .ZN(n531) );
  INV_X1 U441 ( .A(n563), .ZN(n528) );
  INV_X1 U442 ( .A(n516), .ZN(n502) );
  NAND2_X1 U443 ( .A1(n379), .A2(n502), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n380), .B(KEYINPUT89), .ZN(n526) );
  NAND2_X1 U445 ( .A1(n528), .A2(n526), .ZN(n381) );
  NOR2_X1 U446 ( .A1(n531), .A2(n381), .ZN(n382) );
  NOR2_X1 U447 ( .A1(n383), .A2(n382), .ZN(n482) );
  XOR2_X1 U448 ( .A(KEYINPUT78), .B(G64GAT), .Z(n385) );
  XNOR2_X1 U449 ( .A(G127GAT), .B(G183GAT), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n400) );
  XOR2_X1 U451 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n387) );
  XNOR2_X1 U452 ( .A(KEYINPUT15), .B(KEYINPUT79), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n392) );
  XNOR2_X1 U454 ( .A(G71GAT), .B(G57GAT), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n388), .B(KEYINPUT13), .ZN(n423) );
  XOR2_X1 U456 ( .A(KEYINPUT77), .B(n423), .Z(n390) );
  NAND2_X1 U457 ( .A1(G231GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n398) );
  XOR2_X1 U460 ( .A(G211GAT), .B(n393), .Z(n396) );
  XNOR2_X1 U461 ( .A(G15GAT), .B(G1GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n394), .B(G8GAT), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n405), .B(G78GAT), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U466 ( .A(n400), .B(n399), .Z(n479) );
  INV_X1 U467 ( .A(n479), .ZN(n582) );
  XNOR2_X1 U468 ( .A(n402), .B(KEYINPUT94), .ZN(n403) );
  NOR2_X1 U469 ( .A1(n462), .A2(n403), .ZN(n404) );
  XOR2_X1 U470 ( .A(KEYINPUT37), .B(n404), .Z(n515) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n419) );
  XOR2_X1 U472 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n408) );
  NAND2_X1 U473 ( .A1(G229GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U475 ( .A(n409), .B(KEYINPUT30), .Z(n417) );
  XOR2_X1 U476 ( .A(G22GAT), .B(G141GAT), .Z(n411) );
  XNOR2_X1 U477 ( .A(G50GAT), .B(G36GAT), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U479 ( .A(KEYINPUT67), .B(G113GAT), .Z(n413) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(G197GAT), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  INV_X1 U484 ( .A(n578), .ZN(n447) );
  XOR2_X1 U485 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n421) );
  XNOR2_X1 U486 ( .A(G120GAT), .B(G204GAT), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n435) );
  XOR2_X1 U488 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U489 ( .A1(G230GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U491 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n427) );
  XNOR2_X1 U492 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U495 ( .A(n431), .B(n430), .Z(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U497 ( .A(n435), .B(n434), .Z(n445) );
  INV_X1 U498 ( .A(n445), .ZN(n467) );
  NOR2_X1 U499 ( .A1(n447), .A2(n467), .ZN(n483) );
  NAND2_X1 U500 ( .A1(n515), .A2(n483), .ZN(n437) );
  XNOR2_X1 U501 ( .A(KEYINPUT95), .B(KEYINPUT38), .ZN(n436) );
  NAND2_X1 U502 ( .A1(n496), .A2(n531), .ZN(n440) );
  XOR2_X1 U503 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n438) );
  NOR2_X1 U504 ( .A1(n479), .A2(n462), .ZN(n442) );
  XNOR2_X1 U505 ( .A(KEYINPUT45), .B(KEYINPUT107), .ZN(n441) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n443) );
  NOR2_X1 U507 ( .A1(n578), .A2(n443), .ZN(n444) );
  NAND2_X1 U508 ( .A1(n445), .A2(n444), .ZN(n456) );
  XNOR2_X1 U509 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n454) );
  INV_X1 U510 ( .A(KEYINPUT41), .ZN(n446) );
  XNOR2_X1 U511 ( .A(n446), .B(n445), .ZN(n534) );
  NOR2_X1 U512 ( .A1(n534), .A2(n447), .ZN(n448) );
  XNOR2_X1 U513 ( .A(n448), .B(KEYINPUT46), .ZN(n449) );
  NOR2_X1 U514 ( .A1(n582), .A2(n449), .ZN(n450) );
  XNOR2_X1 U515 ( .A(n450), .B(KEYINPUT104), .ZN(n451) );
  NAND2_X1 U516 ( .A1(n451), .A2(n560), .ZN(n452) );
  XNOR2_X1 U517 ( .A(n452), .B(KEYINPUT47), .ZN(n453) );
  XNOR2_X1 U518 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U519 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n457), .B(KEYINPUT48), .ZN(n527) );
  NAND2_X1 U521 ( .A1(n527), .A2(n505), .ZN(n459) );
  NOR2_X1 U522 ( .A1(n502), .A2(n460), .ZN(n471) );
  NAND2_X1 U523 ( .A1(n546), .A2(n471), .ZN(n461) );
  XOR2_X1 U524 ( .A(n461), .B(KEYINPUT123), .Z(n466) );
  NOR2_X1 U525 ( .A1(n462), .A2(n466), .ZN(n465) );
  XNOR2_X1 U526 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n463) );
  INV_X1 U527 ( .A(n466), .ZN(n581) );
  NAND2_X1 U528 ( .A1(n581), .A2(n467), .ZN(n470) );
  XOR2_X1 U529 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n468) );
  INV_X1 U530 ( .A(G190GAT), .ZN(n478) );
  XOR2_X1 U531 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n476) );
  AND2_X1 U532 ( .A1(n542), .A2(n563), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U534 ( .A(KEYINPUT55), .B(n473), .ZN(n564) );
  NAND2_X1 U535 ( .A1(n474), .A2(n564), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT34), .B(KEYINPUT93), .Z(n486) );
  NOR2_X1 U539 ( .A1(n479), .A2(n542), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  NOR2_X1 U541 ( .A1(n482), .A2(n481), .ZN(n500) );
  NAND2_X1 U542 ( .A1(n483), .A2(n500), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT92), .B(n484), .Z(n491) );
  NAND2_X1 U544 ( .A1(n502), .A2(n491), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n491), .A2(n505), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U550 ( .A1(n491), .A2(n563), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U552 ( .A1(n491), .A2(n531), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NAND2_X1 U555 ( .A1(n502), .A2(n496), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n496), .A2(n505), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n496), .A2(n563), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  NOR2_X1 U563 ( .A1(n578), .A2(n534), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n499), .B(KEYINPUT98), .ZN(n514) );
  NAND2_X1 U565 ( .A1(n514), .A2(n500), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(KEYINPUT99), .ZN(n509) );
  NAND2_X1 U567 ( .A1(n502), .A2(n509), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n509), .A2(n505), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT100), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n563), .A2(n509), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT102), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n531), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n513) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT101), .Z(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n522) );
  NOR2_X1 U580 ( .A1(n516), .A2(n522), .ZN(n517) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n522), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT103), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NOR2_X1 U585 ( .A1(n528), .A2(n522), .ZN(n521) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U588 ( .A(G106GAT), .B(n524), .Z(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT44), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT109), .Z(n533) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n547) );
  NOR2_X1 U592 ( .A1(n528), .A2(n547), .ZN(n529) );
  XOR2_X1 U593 ( .A(KEYINPUT108), .B(n529), .Z(n530) );
  NOR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n543), .A2(n578), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT110), .B(KEYINPUT49), .Z(n536) );
  INV_X1 U598 ( .A(n534), .ZN(n569) );
  NAND2_X1 U599 ( .A1(n543), .A2(n569), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(n537), .ZN(G1341GAT) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(KEYINPUT111), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U604 ( .A1(n543), .A2(n582), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT113), .Z(n550) );
  INV_X1 U611 ( .A(n546), .ZN(n548) );
  NOR2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n558), .A2(n578), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XOR2_X1 U616 ( .A(KEYINPUT114), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U617 ( .A1(n558), .A2(n569), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n556) );
  NAND2_X1 U621 ( .A1(n558), .A2(n582), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  INV_X1 U624 ( .A(n558), .ZN(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  AND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n572), .A2(n578), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n567) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT119), .B(n568), .Z(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  XOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT121), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n582), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT124), .B(n577), .Z(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
endmodule

