//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n610,
    new_n611, new_n612, new_n613, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n655, new_n658, new_n660, new_n661,
    new_n662, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT67), .B(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G137), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n476), .B1(new_n479), .B2(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n474), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(new_n469), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G125), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(KEYINPUT68), .B(new_n482), .C1(new_n487), .C2(new_n476), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n473), .B1(new_n481), .B2(new_n488), .ZN(G160));
  AND3_X1   g064(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT3), .B1(new_n466), .B2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(new_n469), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n469), .A2(G112), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n492), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G136), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT70), .B1(new_n497), .B2(G136), .ZN(new_n501));
  OAI221_X1 g076(.A(new_n494), .B1(new_n495), .B2(new_n496), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n502), .B(new_n503), .ZN(G162));
  AND2_X1   g079(.A1(KEYINPUT72), .A2(G114), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT72), .A2(G114), .ZN(new_n506));
  OAI21_X1  g081(.A(G2105), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(G126), .A2(G2105), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n490), .B2(new_n491), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n469), .B(G138), .C1(new_n490), .C2(new_n491), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT4), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT4), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT4), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(new_n519), .B1(new_n477), .B2(new_n478), .ZN(new_n520));
  INV_X1    g095(.A(G2105), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT67), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G2105), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n522), .A2(new_n524), .A3(G138), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n513), .B1(new_n515), .B2(new_n526), .ZN(G164));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  AND3_X1   g105(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(G543), .B1(KEYINPUT74), .B2(KEYINPUT5), .ZN(new_n532));
  AND2_X1   g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(KEYINPUT6), .A2(G651), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G88), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n529), .A2(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(G75), .A2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n531), .A2(new_n532), .ZN(new_n539));
  INV_X1    g114(.A(G62), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n537), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(KEYINPUT75), .A3(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(G303));
  INV_X1    g121(.A(G303), .ZN(G166));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT76), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT7), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n551), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n550), .B1(new_n549), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g130(.A(G63), .B(G651), .C1(new_n531), .C2(new_n532), .ZN(new_n556));
  OAI211_X1 g131(.A(G51), .B(G543), .C1(new_n533), .C2(new_n534), .ZN(new_n557));
  INV_X1    g132(.A(G89), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n535), .C2(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT77), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n549), .A2(new_n552), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT7), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n556), .A2(new_n557), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  NAND2_X1  g141(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n567));
  INV_X1    g142(.A(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(G89), .A3(new_n528), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n560), .A2(new_n573), .ZN(G168));
  INV_X1    g149(.A(G52), .ZN(new_n575));
  INV_X1    g150(.A(G90), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n529), .A2(new_n575), .B1(new_n535), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n571), .A2(G64), .ZN(new_n578));
  NAND2_X1  g153(.A1(G77), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n577), .B1(new_n581), .B2(KEYINPUT78), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n583), .A3(G651), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(G171));
  AOI22_X1  g160(.A1(new_n571), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G651), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G43), .ZN(new_n589));
  INV_X1    g164(.A(G81), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n529), .A2(new_n589), .B1(new_n535), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G860), .ZN(G153));
  NAND4_X1  g168(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g169(.A1(G1), .A2(G3), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT8), .ZN(new_n596));
  NAND4_X1  g171(.A1(G319), .A2(G483), .A3(G661), .A4(new_n596), .ZN(G188));
  INV_X1    g172(.A(G53), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n529), .A2(KEYINPUT9), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT9), .B1(new_n529), .B2(new_n598), .ZN(new_n600));
  NAND2_X1  g175(.A1(G78), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G65), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n539), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n599), .A2(new_n600), .B1(G651), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G91), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n535), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT79), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(G299));
  NAND2_X1  g183(.A1(new_n582), .A2(new_n584), .ZN(G301));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n610));
  NAND2_X1  g185(.A1(G168), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n560), .A2(new_n573), .A3(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G286));
  INV_X1    g189(.A(G49), .ZN(new_n615));
  INV_X1    g190(.A(G87), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n529), .A2(new_n615), .B1(new_n535), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G651), .C1(new_n571), .C2(G74), .ZN(new_n619));
  OAI21_X1  g194(.A(G651), .B1(new_n571), .B2(G74), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT81), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n617), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(G288));
  NAND2_X1  g198(.A1(G73), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(G61), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n539), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G651), .ZN(new_n627));
  INV_X1    g202(.A(new_n535), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G86), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n528), .A2(G48), .A3(G543), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(G305));
  INV_X1    g206(.A(G47), .ZN(new_n632));
  INV_X1    g207(.A(G85), .ZN(new_n633));
  OAI22_X1  g208(.A1(new_n529), .A2(new_n632), .B1(new_n535), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT82), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n636), .B1(new_n535), .B2(new_n633), .C1(new_n632), .C2(new_n529), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n571), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(new_n587), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(G290));
  NAND2_X1  g216(.A1(G301), .A2(G868), .ZN(new_n642));
  INV_X1    g217(.A(G92), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n535), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT10), .ZN(new_n645));
  NAND2_X1  g220(.A1(G79), .A2(G543), .ZN(new_n646));
  INV_X1    g221(.A(G66), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n539), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n528), .A2(G543), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n648), .A2(G651), .B1(new_n649), .B2(G54), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n642), .B1(G868), .B2(new_n652), .ZN(G284));
  OAI21_X1  g228(.A(new_n642), .B1(G868), .B2(new_n652), .ZN(G321));
  NOR2_X1   g229(.A1(G299), .A2(G868), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n613), .B2(G868), .ZN(G297));
  AOI21_X1  g231(.A(new_n655), .B1(new_n613), .B2(G868), .ZN(G280));
  XOR2_X1   g232(.A(KEYINPUT83), .B(G559), .Z(new_n658));
  OAI21_X1  g233(.A(new_n652), .B1(G860), .B2(new_n658), .ZN(G148));
  AND2_X1   g234(.A1(new_n652), .A2(new_n658), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G868), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(G868), .B2(new_n592), .ZN(G323));
  XNOR2_X1  g238(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g239(.A1(new_n479), .A2(new_n471), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT12), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT13), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n497), .A2(G135), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n493), .A2(G123), .ZN(new_n670));
  OAI221_X1 g245(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n469), .C2(G111), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2096), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n673), .ZN(G156));
  INV_X1    g249(.A(KEYINPUT14), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2427), .B(G2438), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2430), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT15), .B(G2435), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n678), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2451), .B(G2454), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT16), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1341), .B(G1348), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n680), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2443), .B(G2446), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G14), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(G401));
  XOR2_X1   g265(.A(G2084), .B(G2090), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT84), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2067), .B(G2678), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT85), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G2072), .B(G2078), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT18), .Z(new_n699));
  OAI21_X1  g274(.A(KEYINPUT17), .B1(new_n692), .B2(new_n694), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n695), .B1(new_n700), .B2(new_n696), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n696), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G2100), .ZN(new_n704));
  INV_X1    g279(.A(G2100), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n699), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT86), .B(G2096), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n707), .A2(new_n709), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(G227));
  XOR2_X1   g288(.A(G1971), .B(G1976), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT19), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1956), .B(G2474), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1961), .B(G1966), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n715), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(new_n718), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT20), .Z(new_n722));
  AOI211_X1 g297(.A(new_n720), .B(new_n722), .C1(new_n715), .C2(new_n719), .ZN(new_n723));
  XOR2_X1   g298(.A(G1991), .B(G1996), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT88), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n723), .B(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(G1981), .B(G1986), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT87), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n727), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(G229));
  XNOR2_X1  g308(.A(new_n502), .B(KEYINPUT71), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G35), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n735), .B2(new_n737), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2090), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G20), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT100), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT23), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G299), .B2(G16), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1956), .ZN(new_n749));
  INV_X1    g324(.A(new_n740), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT99), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n750), .A2(new_n751), .A3(G2090), .A4(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n743), .A2(KEYINPUT101), .A3(new_n749), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n741), .A2(G2090), .ZN(new_n755));
  NOR2_X1   g330(.A1(G4), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n652), .B2(G16), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT93), .Z(new_n758));
  INV_X1    g333(.A(G1348), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT24), .ZN(new_n762));
  INV_X1    g337(.A(G34), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G160), .B2(new_n736), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G2084), .ZN(new_n767));
  OR2_X1    g342(.A1(G29), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n497), .A2(G139), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n770), .B(new_n771), .C1(new_n469), .C2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(new_n736), .ZN(new_n774));
  INV_X1    g349(.A(G2072), .ZN(new_n775));
  NOR2_X1   g350(.A1(G27), .A2(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G164), .B2(G29), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n774), .A2(new_n775), .B1(G2078), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT30), .B(G28), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n779), .A2(new_n736), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n672), .B2(new_n736), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n766), .A2(G2084), .ZN(new_n785));
  AND4_X1   g360(.A1(new_n767), .A2(new_n778), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n760), .A2(new_n761), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n736), .A2(G26), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT28), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n497), .A2(G140), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n469), .A2(G116), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n493), .A2(G128), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2067), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n744), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n744), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G1966), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n744), .A2(G5), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G171), .B2(new_n744), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n799), .B(new_n802), .C1(G1961), .C2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n736), .A2(G32), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n497), .A2(G141), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT95), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n471), .A2(G105), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT96), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT96), .ZN(new_n811));
  NAND3_X1  g386(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT26), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n810), .A2(new_n811), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n493), .A2(G129), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n808), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n806), .B1(new_n819), .B2(G29), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT27), .B(G1996), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(G16), .A2(G19), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n592), .B2(G16), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G1341), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n774), .B2(new_n775), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(G1341), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n777), .A2(G2078), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n804), .A2(G1961), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n801), .A2(G1966), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n822), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NOR4_X1   g407(.A1(new_n755), .A2(new_n787), .A3(new_n805), .A4(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n753), .A2(new_n749), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n751), .B1(new_n741), .B2(G2090), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n754), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n744), .A2(G6), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G305), .B2(G16), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT90), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT32), .B(G1981), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT91), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n841), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n744), .A2(G22), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G166), .B2(new_n744), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT92), .Z(new_n847));
  AOI21_X1  g422(.A(new_n844), .B1(G1971), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n744), .A2(G23), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n622), .B2(new_n744), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT33), .Z(new_n851));
  INV_X1    g426(.A(G1976), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n848), .B(new_n853), .C1(G1971), .C2(new_n847), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT34), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n736), .A2(G25), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n493), .A2(G119), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT89), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n469), .A2(G107), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n497), .A2(G131), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n857), .B1(new_n865), .B2(new_n736), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G1991), .Z(new_n867));
  XOR2_X1   g442(.A(new_n866), .B(new_n867), .Z(new_n868));
  MUX2_X1   g443(.A(G24), .B(G290), .S(G16), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G1986), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n854), .B2(KEYINPUT34), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT36), .B1(new_n856), .B2(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n854), .A2(KEYINPUT34), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n874), .A2(new_n875), .A3(new_n855), .A4(new_n871), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n838), .B1(new_n873), .B2(new_n876), .ZN(G311));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n876), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n878), .A2(new_n754), .A3(new_n837), .A4(new_n833), .ZN(G150));
  NAND2_X1  g454(.A1(G80), .A2(G543), .ZN(new_n880));
  INV_X1    g455(.A(G67), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n539), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G651), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  OAI211_X1 g459(.A(G55), .B(G543), .C1(new_n533), .C2(new_n534), .ZN(new_n885));
  INV_X1    g460(.A(G93), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n884), .B(new_n885), .C1(new_n535), .C2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n571), .A2(G93), .A3(new_n528), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n884), .B1(new_n889), .B2(new_n885), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n883), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G860), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT37), .Z(new_n893));
  NAND2_X1  g468(.A1(new_n652), .A2(G559), .ZN(new_n894));
  XOR2_X1   g469(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n592), .ZN(new_n899));
  OAI211_X1 g474(.A(KEYINPUT104), .B(new_n883), .C1(new_n888), .C2(new_n890), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n891), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT104), .A3(new_n592), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n896), .B(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT39), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT105), .ZN(new_n909));
  INV_X1    g484(.A(G860), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n907), .B2(KEYINPUT39), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n893), .B1(new_n909), .B2(new_n911), .ZN(G145));
  XNOR2_X1  g487(.A(new_n864), .B(new_n666), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n493), .A2(G130), .ZN(new_n914));
  OAI221_X1 g489(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(G142), .B2(new_n497), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n913), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n773), .A2(new_n919), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n468), .A2(new_n511), .B1(new_n507), .B2(new_n509), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n516), .B1(new_n525), .B2(new_n468), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n522), .A2(new_n524), .A3(G138), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n923), .A2(new_n485), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n797), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n792), .A2(G164), .A3(new_n796), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n819), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n929), .A2(new_n930), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n920), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n933), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n773), .B(new_n919), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n918), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n939));
  XNOR2_X1  g514(.A(G162), .B(new_n672), .ZN(new_n940));
  INV_X1    g515(.A(G160), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n934), .B(new_n937), .C1(new_n918), .C2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n940), .B(G160), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n934), .A2(new_n937), .A3(new_n918), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n938), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G37), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g526(.A1(G290), .A2(new_n622), .ZN(new_n952));
  NAND3_X1  g527(.A1(G288), .A2(new_n638), .A3(new_n640), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G305), .ZN(new_n955));
  NAND2_X1  g530(.A1(G303), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n544), .A2(new_n545), .A3(G305), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n952), .A2(new_n953), .A3(new_n956), .A4(new_n957), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT42), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n959), .A2(KEYINPUT108), .A3(new_n960), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT108), .B1(new_n959), .B2(new_n960), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n961), .B1(new_n964), .B2(KEYINPUT42), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n661), .B(new_n904), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT41), .ZN(new_n967));
  NAND2_X1  g542(.A1(G299), .A2(new_n651), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(G299), .A2(new_n651), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n970), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(KEYINPUT41), .A3(new_n968), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n966), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n969), .A2(new_n970), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(new_n966), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n965), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(G868), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(G868), .B2(new_n902), .ZN(G295));
  OAI21_X1  g555(.A(new_n979), .B1(G868), .B2(new_n902), .ZN(G331));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n982));
  AOI21_X1  g557(.A(G168), .B1(new_n584), .B2(new_n582), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n613), .B2(G171), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n976), .B1(new_n984), .B2(new_n904), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n560), .A2(new_n573), .A3(KEYINPUT80), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT80), .B1(new_n560), .B2(new_n573), .ZN(new_n987));
  OAI21_X1  g562(.A(G171), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G168), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G301), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n988), .A2(new_n903), .A3(new_n901), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n984), .A2(KEYINPUT109), .A3(new_n904), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n985), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n984), .A2(new_n904), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n974), .B1(new_n996), .B2(new_n991), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n964), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n962), .A2(new_n963), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n976), .A3(new_n991), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n984), .A2(new_n904), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n993), .B2(new_n994), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n999), .B(new_n1000), .C1(new_n1002), .C2(new_n974), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n1003), .A3(new_n949), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n998), .A2(new_n1003), .A3(KEYINPUT111), .A4(new_n949), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n982), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n991), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n985), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n993), .A2(new_n994), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n996), .ZN(new_n1012));
  INV_X1    g587(.A(new_n974), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(new_n999), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1003), .A2(new_n949), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT43), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT44), .B1(new_n1008), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1011), .A2(new_n976), .A3(new_n996), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1013), .B1(new_n1009), .B2(new_n1001), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(G37), .B1(new_n1023), .B2(new_n964), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(KEYINPUT110), .A3(new_n982), .A4(new_n1003), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT43), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n998), .A2(new_n1003), .A3(new_n982), .A4(new_n949), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1020), .A2(new_n1032), .ZN(G397));
  NAND2_X1  g608(.A1(G160), .A2(G40), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(G164), .B2(G1384), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n819), .B(G1996), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n797), .B(G2067), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n864), .B(new_n867), .Z(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(G290), .B(G1986), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1037), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G303), .A2(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n926), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT50), .ZN(new_n1054));
  INV_X1    g629(.A(G40), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1055), .B(new_n473), .C1(new_n481), .C2(new_n488), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n926), .A2(new_n1057), .A3(new_n1052), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G2090), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n514), .A2(KEYINPUT4), .B1(new_n520), .B2(new_n525), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT45), .B(new_n1052), .C1(new_n1061), .C2(new_n513), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT45), .B1(new_n926), .B2(new_n1052), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1053), .A2(KEYINPUT112), .A3(new_n1035), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1056), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1971), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1060), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1051), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n571), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n630), .B1(new_n1074), .B2(new_n587), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT116), .B(G86), .Z(new_n1076));
  NOR2_X1   g651(.A1(new_n535), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(G1981), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n627), .A2(new_n1079), .A3(new_n629), .A4(new_n630), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(KEYINPUT117), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT49), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(G1981), .C1(new_n1075), .C2(new_n1077), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G164), .A2(G1384), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1072), .B1(new_n1056), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1082), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT118), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT49), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1087), .A4(new_n1085), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT114), .B(G1976), .Z(new_n1095));
  NOR2_X1   g670(.A1(new_n622), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(G8), .B(new_n1096), .C1(new_n1034), .C2(new_n1053), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(G8), .B1(new_n1034), .B2(new_n1053), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT115), .B1(G288), .B2(new_n852), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1097), .B(new_n1098), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1090), .A2(new_n1094), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1036), .A2(new_n1063), .A3(new_n1062), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1034), .B1(new_n1106), .B2(new_n1067), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G1971), .ZN(new_n1108));
  OAI211_X1 g683(.A(G8), .B(new_n1050), .C1(new_n1108), .C2(new_n1060), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1073), .A2(new_n1105), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1072), .B1(KEYINPUT122), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1062), .B1(new_n1065), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1086), .A2(KEYINPUT120), .A3(KEYINPUT45), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1056), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1966), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1119));
  INV_X1    g694(.A(G2084), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1117), .A2(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1113), .B1(new_n1121), .B2(G168), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1111), .A2(KEYINPUT122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1121), .A2(new_n1072), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1122), .A2(new_n1124), .B1(new_n1126), .B2(new_n989), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1110), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G2078), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1107), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT123), .B(G1961), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1059), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(KEYINPUT53), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n470), .A2(G40), .A3(new_n472), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n480), .A2(new_n469), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1065), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1062), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1129), .B1(new_n1133), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1132), .B(new_n1056), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1130), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1059), .A2(new_n1134), .B1(new_n1140), .B2(new_n1062), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(KEYINPUT126), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G301), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1115), .A2(new_n1116), .A3(new_n1056), .A4(new_n1137), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1135), .ZN(new_n1150));
  OAI21_X1  g725(.A(G301), .B1(new_n1133), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT54), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1145), .A2(new_n1153), .A3(G301), .A4(new_n1146), .ZN(new_n1154));
  OAI21_X1  g729(.A(G171), .B1(new_n1133), .B2(new_n1150), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1142), .B1(new_n1144), .B2(new_n1130), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n1158), .B2(G301), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1148), .A2(new_n1152), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1128), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT56), .B(G2072), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1107), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(G1956), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1059), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n1166));
  XNOR2_X1  g741(.A(G299), .B(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1163), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1034), .A2(new_n1053), .ZN(new_n1170));
  INV_X1    g745(.A(G2067), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n759), .A2(new_n1059), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(new_n651), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1168), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n1175));
  INV_X1    g750(.A(G1996), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1056), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n1106), .B2(new_n1067), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT58), .B(G1341), .Z(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1170), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n592), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT59), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1184), .B(new_n592), .C1(new_n1178), .C2(new_n1181), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1106), .A2(new_n1067), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1187), .A2(new_n1056), .A3(new_n1162), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1167), .A2(new_n1165), .ZN(new_n1189));
  OAI21_X1  g764(.A(KEYINPUT61), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1183), .A2(new_n1186), .B1(new_n1190), .B2(new_n1169), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1167), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(KEYINPUT61), .B1(new_n1194), .B2(new_n1168), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1175), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1194), .A2(KEYINPUT61), .A3(new_n1168), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n1169), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1185), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1197), .A2(new_n1200), .A3(KEYINPUT121), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1172), .A2(KEYINPUT60), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(new_n652), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1205), .B1(KEYINPUT60), .B2(new_n1172), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1196), .A2(new_n1203), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1161), .B1(new_n1174), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT119), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n622), .A2(new_n852), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1100), .B1(new_n1213), .B2(new_n1080), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1210), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1216), .A2(new_n1109), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1209), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g793(.A1(new_n1210), .A2(new_n1212), .B1(new_n1079), .B2(new_n955), .ZN(new_n1219));
  OAI221_X1 g794(.A(KEYINPUT119), .B1(new_n1216), .B2(new_n1109), .C1(new_n1219), .C2(new_n1100), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1121), .A2(G168), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1222), .A2(new_n1112), .A3(new_n1124), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1126), .A2(new_n989), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1226));
  OAI21_X1  g801(.A(KEYINPUT62), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1127), .A2(new_n1125), .A3(new_n1228), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n1110), .A2(new_n1155), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NOR3_X1   g806(.A1(new_n1121), .A2(G286), .A3(new_n1072), .ZN(new_n1232));
  NAND4_X1  g807(.A1(new_n1073), .A2(new_n1105), .A3(new_n1232), .A4(new_n1109), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT63), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1233), .B(new_n1234), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1221), .A2(new_n1231), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1045), .B1(new_n1208), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1037), .B1(new_n1039), .B2(new_n819), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1037), .A2(new_n1176), .ZN(new_n1239));
  XNOR2_X1  g814(.A(new_n1239), .B(KEYINPUT46), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g816(.A(new_n1241), .B(KEYINPUT47), .ZN(new_n1242));
  INV_X1    g817(.A(new_n1037), .ZN(new_n1243));
  NOR3_X1   g818(.A1(new_n1243), .A2(G1986), .A3(G290), .ZN(new_n1244));
  XOR2_X1   g819(.A(new_n1244), .B(KEYINPUT48), .Z(new_n1245));
  OAI21_X1  g820(.A(new_n1245), .B1(new_n1042), .B2(new_n1243), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n865), .A2(new_n867), .ZN(new_n1247));
  OAI22_X1  g822(.A1(new_n1040), .A2(new_n1247), .B1(G2067), .B2(new_n797), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1248), .A2(new_n1037), .ZN(new_n1249));
  AND3_X1   g824(.A1(new_n1242), .A2(new_n1246), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1237), .A2(new_n1250), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g826(.A1(G401), .A2(new_n461), .ZN(new_n1253));
  INV_X1    g827(.A(new_n1253), .ZN(new_n1254));
  OAI21_X1  g828(.A(KEYINPUT127), .B1(G227), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1256));
  OAI211_X1 g830(.A(new_n1256), .B(new_n1253), .C1(new_n711), .C2(new_n712), .ZN(new_n1257));
  AND3_X1   g831(.A1(new_n1255), .A2(new_n732), .A3(new_n1257), .ZN(new_n1258));
  AND3_X1   g832(.A1(new_n1258), .A2(new_n1030), .A3(new_n950), .ZN(G308));
  NAND3_X1  g833(.A1(new_n1258), .A2(new_n1030), .A3(new_n950), .ZN(G225));
endmodule


