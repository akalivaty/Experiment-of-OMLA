//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n212), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT66), .B(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(KEYINPUT67), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n228), .A2(KEYINPUT67), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n209), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n221), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n202), .A2(G68), .ZN(new_n248));
  INV_X1    g0048(.A(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n247), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  INV_X1    g0055(.A(new_n213), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n261), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(G226), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G222), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G223), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(new_n264), .C1(G77), .C2(new_n267), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(G200), .B2(new_n273), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT68), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT8), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT8), .A2(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n207), .A2(G33), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n279), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n213), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n207), .A3(G1), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G50), .ZN(new_n293));
  INV_X1    g0093(.A(new_n287), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n206), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n293), .B1(new_n297), .B2(G50), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n277), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n289), .A2(new_n298), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n303), .A2(KEYINPUT9), .A3(new_n300), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n276), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n273), .A2(G200), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT76), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n276), .B(new_n308), .C1(new_n302), .C2(new_n304), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n263), .B1(G244), .B2(new_n265), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G232), .A2(G1698), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n269), .A2(G238), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n267), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT71), .B(G107), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n264), .C1(new_n267), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G179), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n320), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT8), .B(G58), .Z(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT72), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT15), .B(G87), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n325), .A2(new_n326), .B1(new_n284), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n287), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n291), .A2(new_n223), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OR3_X1    g0132(.A1(new_n291), .A2(new_n287), .A3(KEYINPUT73), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT73), .B1(new_n291), .B2(new_n287), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n333), .A2(G77), .A3(new_n295), .A4(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT74), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n323), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n320), .A2(G200), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n313), .A2(G190), .A3(new_n319), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n332), .A2(new_n336), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n256), .A2(new_n257), .ZN(new_n343));
  INV_X1    g0143(.A(G232), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G1698), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n267), .B(new_n345), .C1(G226), .C2(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n262), .B1(new_n350), .B2(new_n227), .ZN(new_n351));
  OR3_X1    g0151(.A1(new_n348), .A2(new_n351), .A3(KEYINPUT13), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT13), .B1(new_n348), .B2(new_n351), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G169), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT14), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(new_n357), .A3(G169), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n356), .B(new_n358), .C1(new_n359), .C2(new_n354), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT12), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n291), .A2(new_n361), .A3(new_n249), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(KEYINPUT77), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT12), .B1(new_n292), .B2(new_n225), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(KEYINPUT77), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n333), .A2(G68), .A3(new_n295), .A4(new_n334), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(KEYINPUT78), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n225), .A2(new_n207), .ZN(new_n369));
  INV_X1    g0169(.A(new_n278), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n370), .A2(new_n202), .B1(new_n284), .B2(new_n223), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n287), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT11), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT78), .B1(new_n366), .B2(new_n367), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n342), .A2(KEYINPUT75), .B1(new_n360), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n352), .A2(G190), .A3(new_n353), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n354), .A2(G200), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT79), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n376), .A2(new_n380), .A3(KEYINPUT79), .A4(new_n379), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n299), .A2(new_n301), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n266), .A2(new_n359), .A3(new_n272), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT70), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n273), .A2(new_n322), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n338), .A2(new_n341), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AND4_X1   g0193(.A1(new_n312), .A2(new_n378), .A3(new_n385), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT82), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT66), .A2(G68), .ZN(new_n396));
  AND2_X1   g0196(.A1(KEYINPUT66), .A2(G68), .ZN(new_n397));
  AND2_X1   g0197(.A1(KEYINPUT68), .A2(G58), .ZN(new_n398));
  NOR2_X1   g0198(.A1(KEYINPUT68), .A2(G58), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n396), .A2(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n207), .B1(new_n400), .B2(new_n215), .ZN(new_n401));
  INV_X1    g0201(.A(G159), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n370), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n395), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n403), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n201), .B1(new_n225), .B2(new_n280), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT82), .B(new_n405), .C1(new_n406), .C2(new_n207), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT3), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT80), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT80), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT3), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n412), .A3(G33), .ZN(new_n413));
  INV_X1    g0213(.A(G33), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT3), .ZN(new_n415));
  AOI21_X1  g0215(.A(G20), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n249), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n415), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(G33), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT7), .B1(new_n421), .B2(G20), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT81), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n418), .A2(KEYINPUT81), .A3(new_n422), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n408), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT84), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n409), .A2(G33), .ZN(new_n428));
  AOI21_X1  g0228(.A(G20), .B1(new_n428), .B2(new_n415), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(KEYINPUT7), .ZN(new_n430));
  OAI211_X1 g0230(.A(KEYINPUT84), .B(new_n417), .C1(new_n267), .C2(G20), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(KEYINPUT85), .B(new_n428), .C1(new_n420), .C2(G33), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n410), .A2(new_n412), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT85), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n414), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n433), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n226), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n404), .A2(new_n407), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n426), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n425), .A2(new_n440), .A3(new_n287), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n283), .A2(new_n292), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n283), .B2(new_n297), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n265), .A2(G232), .B1(new_n258), .B2(new_n261), .ZN(new_n444));
  INV_X1    g0244(.A(G87), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n414), .A2(new_n445), .ZN(new_n446));
  MUX2_X1   g0246(.A(G223), .B(G226), .S(G1698), .Z(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n421), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n444), .B1(new_n448), .B2(new_n343), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n274), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(G200), .B2(new_n449), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n441), .A2(new_n443), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT18), .ZN(new_n455));
  INV_X1    g0255(.A(new_n443), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n418), .A2(new_n422), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n418), .A2(KEYINPUT81), .A3(new_n422), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n294), .B1(new_n461), .B2(new_n408), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n456), .B1(new_n462), .B2(new_n440), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n447), .A2(new_n413), .A3(new_n415), .ZN(new_n464));
  INV_X1    g0264(.A(new_n446), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n343), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n262), .B1(new_n350), .B2(new_n344), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n322), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n359), .B(new_n444), .C1(new_n448), .C2(new_n343), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT86), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n455), .B1(new_n463), .B2(new_n473), .ZN(new_n474));
  AOI211_X1 g0274(.A(new_n455), .B(new_n473), .C1(new_n441), .C2(new_n443), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(KEYINPUT87), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n441), .B2(new_n443), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n477), .A2(KEYINPUT87), .A3(KEYINPUT18), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n454), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n394), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT24), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n421), .A2(new_n207), .A3(G87), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT95), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n421), .A2(KEYINPUT95), .A3(new_n207), .A4(G87), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(KEYINPUT22), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n267), .ZN(new_n488));
  OR4_X1    g0288(.A1(KEYINPUT22), .A2(new_n488), .A3(G20), .A4(new_n445), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT89), .B(G116), .ZN(new_n491));
  OR4_X1    g0291(.A1(KEYINPUT96), .A2(new_n491), .A3(G20), .A4(new_n414), .ZN(new_n492));
  INV_X1    g0292(.A(new_n491), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(new_n207), .A3(G33), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT96), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n317), .A2(G20), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(KEYINPUT23), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n482), .B1(new_n490), .B2(new_n500), .ZN(new_n501));
  AOI211_X1 g0301(.A(KEYINPUT24), .B(new_n499), .C1(new_n487), .C2(new_n489), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n287), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G107), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT25), .B1(new_n291), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n504), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n414), .A2(G1), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n291), .A2(new_n287), .A3(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n506), .A2(new_n507), .B1(new_n509), .B2(G107), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n413), .A2(new_n415), .ZN(new_n512));
  INV_X1    g0312(.A(G257), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G1698), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(G250), .B2(G1698), .ZN(new_n515));
  INV_X1    g0315(.A(G294), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n512), .A2(new_n515), .B1(new_n414), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(KEYINPUT5), .B(G41), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n260), .A2(G1), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n343), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n264), .A2(new_n517), .B1(new_n522), .B2(G264), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n258), .A2(new_n519), .A3(new_n518), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n359), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n527), .B2(G169), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT97), .B1(new_n511), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT97), .ZN(new_n531));
  AOI211_X1 g0331(.A(new_n531), .B(new_n528), .C1(new_n503), .C2(new_n510), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n526), .A2(new_n274), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(G200), .B2(new_n526), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n503), .A2(new_n510), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n258), .A2(new_n519), .ZN(new_n538));
  INV_X1    g0338(.A(G250), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n519), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n343), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G238), .A2(G1698), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n224), .B2(G1698), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n421), .A2(new_n544), .B1(G33), .B2(new_n493), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n542), .B1(new_n545), .B2(new_n343), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n322), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(G179), .B2(new_n546), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n421), .A2(new_n207), .A3(G68), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  INV_X1    g0351(.A(G97), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n317), .A2(new_n445), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n347), .A2(new_n207), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n284), .A2(KEYINPUT19), .A3(new_n552), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n287), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT91), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n327), .B(KEYINPUT90), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n291), .A2(new_n287), .A3(new_n508), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT90), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n327), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(KEYINPUT91), .A3(new_n509), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n327), .A2(new_n291), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n558), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT92), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n557), .A2(new_n287), .B1(new_n291), .B2(new_n327), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT92), .B1(new_n571), .B2(new_n566), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n549), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT93), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n509), .A2(G87), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n546), .A2(G200), .ZN(new_n577));
  INV_X1    g0377(.A(new_n546), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n573), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n568), .A2(new_n569), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n571), .A2(KEYINPUT92), .A3(new_n566), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n548), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND4_X1   g0384(.A1(new_n571), .A2(new_n579), .A3(new_n575), .A4(new_n577), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT93), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n224), .A2(G1698), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT4), .B1(new_n421), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G283), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n269), .A2(KEYINPUT4), .A3(G244), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n539), .B2(new_n269), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n593), .B2(new_n488), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n264), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n524), .B1(new_n521), .B2(new_n513), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(G190), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT88), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n597), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G200), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n292), .A2(G97), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n509), .B2(G97), .ZN(new_n603));
  XNOR2_X1  g0403(.A(G97), .B(G107), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT6), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n605), .A2(new_n552), .A3(G107), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n608), .A2(new_n207), .B1(new_n223), .B2(new_n370), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n432), .A2(new_n437), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n318), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n601), .B(new_n603), .C1(new_n611), .C2(new_n294), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n603), .B1(new_n611), .B2(new_n294), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n600), .A2(new_n322), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n595), .A2(new_n359), .A3(new_n597), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n599), .A2(new_n612), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT94), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n491), .A2(G20), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n590), .B(new_n207), .C1(G33), .C2(new_n552), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n287), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n620), .A2(KEYINPUT20), .A3(new_n287), .A4(new_n621), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G116), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n508), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n333), .A2(new_n334), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n290), .A2(G1), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n491), .A2(G20), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n626), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  MUX2_X1   g0432(.A(G257), .B(G264), .S(G1698), .Z(new_n633));
  AOI22_X1  g0433(.A1(new_n421), .A2(new_n633), .B1(G303), .B2(new_n488), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n343), .ZN(new_n635));
  INV_X1    g0435(.A(G270), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n524), .B1(new_n521), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(G169), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n619), .B1(new_n632), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT21), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n635), .A2(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G179), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n632), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(G190), .ZN(new_n646));
  INV_X1    g0446(.A(G200), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n646), .B(new_n632), .C1(new_n647), .C2(new_n641), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT21), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n619), .B(new_n649), .C1(new_n632), .C2(new_n638), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n640), .A2(new_n645), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n618), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n587), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n481), .A2(new_n537), .A3(new_n653), .ZN(G372));
  XNOR2_X1  g0454(.A(new_n312), .B(KEYINPUT98), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n360), .A2(new_n377), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n381), .A2(new_n337), .A3(new_n323), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n477), .A2(KEYINPUT18), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n658), .A2(new_n454), .B1(new_n659), .B2(new_n475), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n390), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n481), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n598), .B(KEYINPUT88), .Z(new_n663));
  INV_X1    g0463(.A(new_n601), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n613), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n617), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n663), .A2(new_n665), .B1(new_n613), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n584), .A2(new_n585), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n536), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n640), .A2(new_n650), .A3(new_n645), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n511), .B2(new_n529), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n584), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n614), .A2(new_n617), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n587), .A2(KEYINPUT26), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT26), .B1(new_n668), .B2(new_n675), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n661), .B1(new_n662), .B2(new_n681), .ZN(G369));
  INV_X1    g0482(.A(new_n511), .ZN(new_n683));
  INV_X1    g0483(.A(new_n630), .ZN(new_n684));
  OR3_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .A3(G20), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT27), .B1(new_n684), .B2(G20), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n537), .B1(new_n683), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n511), .A2(new_n529), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n632), .A2(new_n690), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n671), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n651), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT99), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n689), .B(KEYINPUT100), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n511), .A2(new_n529), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n671), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n689), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n537), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n701), .A2(new_n703), .A3(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n210), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n553), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n219), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n653), .A2(new_n533), .A3(new_n536), .A4(new_n702), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n595), .A2(new_n597), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n523), .A3(new_n578), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT30), .B1(new_n717), .B2(new_n642), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n578), .A2(new_n523), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n643), .A2(new_n719), .A3(new_n720), .A4(new_n716), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n546), .A2(new_n359), .ZN(new_n723));
  OR4_X1    g0523(.A1(new_n527), .A2(new_n716), .A3(new_n641), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n689), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  XOR2_X1   g0527(.A(KEYINPUT101), .B(KEYINPUT31), .Z(new_n728));
  NOR2_X1   g0528(.A1(new_n702), .A2(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n726), .A2(new_n727), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n715), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n533), .A2(new_n704), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n584), .B1(new_n734), .B2(new_n670), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n587), .A2(new_n675), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT102), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT26), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n675), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n586), .B2(new_n581), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT102), .B1(new_n741), .B2(KEYINPUT26), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n668), .A2(KEYINPUT26), .A3(new_n675), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n689), .B1(new_n735), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT29), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n680), .A2(new_n702), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT29), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n733), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n714), .B1(new_n750), .B2(G1), .ZN(G364));
  NOR2_X1   g0551(.A1(new_n290), .A2(G20), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G45), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT103), .Z(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n755), .A2(new_n206), .A3(new_n709), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n698), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G330), .B2(new_n696), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n322), .A2(KEYINPUT105), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n207), .B1(KEYINPUT105), .B2(new_n322), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n213), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(G20), .A3(new_n274), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(G329), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n207), .A2(new_n359), .A3(new_n274), .A4(G200), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n267), .B(new_n767), .C1(G322), .C2(new_n768), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n207), .A2(new_n274), .A3(new_n647), .A4(G179), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n207), .B1(new_n764), .B2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n770), .A2(G303), .B1(new_n772), .B2(G294), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n207), .A2(new_n359), .A3(G190), .A4(G200), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT106), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n774), .B1(G311), .B2(new_n780), .ZN(new_n781));
  NOR4_X1   g0581(.A1(new_n207), .A2(new_n647), .A3(G179), .A4(G190), .ZN(new_n782));
  NAND3_X1  g0582(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n274), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n782), .A2(G283), .B1(G326), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n783), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI211_X1 g0588(.A(new_n781), .B(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n782), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n504), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n488), .B(new_n791), .C1(new_n280), .C2(new_n768), .ZN(new_n792));
  INV_X1    g0592(.A(new_n770), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n766), .A2(G159), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n445), .A2(new_n793), .B1(new_n794), .B2(KEYINPUT32), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n787), .A2(new_n249), .B1(new_n771), .B2(new_n552), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n780), .A2(G77), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n794), .A2(KEYINPUT32), .B1(G50), .B2(new_n784), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n792), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n763), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n207), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT104), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n763), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n220), .A2(new_n260), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n708), .A2(new_n421), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(new_n260), .C2(new_n253), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n708), .A2(new_n488), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n809), .A2(G355), .B1(new_n627), .B2(new_n708), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n805), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n756), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n801), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n696), .B2(new_n804), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n758), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n337), .A2(new_n689), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n338), .A2(new_n817), .A3(new_n341), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT108), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n323), .A2(new_n337), .A3(new_n689), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n338), .A2(new_n817), .A3(KEYINPUT108), .A4(new_n341), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n680), .A2(KEYINPUT109), .A3(new_n702), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n677), .B1(new_n741), .B2(KEYINPUT26), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n573), .B1(new_n669), .B2(new_n672), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n702), .B(new_n823), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT109), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n823), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n824), .A2(new_n829), .B1(new_n747), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n733), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n756), .B1(new_n831), .B2(new_n733), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(KEYINPUT110), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(KEYINPUT110), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n762), .A2(new_n802), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT107), .Z(new_n837));
  OAI21_X1  g0637(.A(new_n756), .B1(new_n837), .B2(G77), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n780), .A2(new_n493), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n793), .A2(new_n504), .B1(new_n840), .B2(new_n787), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G303), .B2(new_n784), .ZN(new_n842));
  INV_X1    g0642(.A(G311), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n488), .B1(new_n765), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G294), .B2(new_n768), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n790), .A2(new_n445), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G97), .B2(new_n772), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n839), .A2(new_n842), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n768), .A2(G143), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  INV_X1    g0651(.A(new_n784), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n849), .B1(new_n787), .B2(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G159), .B2(new_n780), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT34), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n512), .B1(G132), .B2(new_n766), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n770), .A2(G50), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n790), .A2(new_n249), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n280), .B2(new_n772), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n854), .A2(KEYINPUT34), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n848), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n838), .B1(new_n862), .B2(new_n762), .ZN(new_n863));
  INV_X1    g0663(.A(new_n802), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n823), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n835), .A2(new_n865), .ZN(G384));
  INV_X1    g0666(.A(new_n608), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n867), .A2(KEYINPUT35), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(KEYINPUT35), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n868), .A2(G116), .A3(new_n214), .A4(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(KEYINPUT111), .B(KEYINPUT36), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n217), .A2(G77), .A3(new_n218), .A4(new_n400), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n206), .B(G13), .C1(new_n873), .C2(new_n248), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n659), .A2(new_n475), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n687), .ZN(new_n877));
  INV_X1    g0677(.A(new_n426), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n439), .B1(new_n459), .B2(new_n460), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n462), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n443), .ZN(new_n881));
  INV_X1    g0681(.A(new_n687), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT112), .B1(new_n480), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n452), .B(KEYINPUT17), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT87), .B1(new_n477), .B2(KEYINPUT18), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(new_n659), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n887), .B2(new_n478), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT112), .ZN(new_n889));
  INV_X1    g0689(.A(new_n883), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n473), .A2(new_n687), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .A3(new_n452), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n441), .A2(new_n443), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n452), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n892), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n895), .A2(new_n900), .A3(KEYINPUT38), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n480), .A2(KEYINPUT112), .A3(new_n883), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT113), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n903), .B1(new_n884), .B2(new_n891), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT113), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n902), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n338), .A2(new_n689), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n827), .A2(new_n828), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n827), .A2(new_n828), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n377), .A2(new_n689), .ZN(new_n918));
  INV_X1    g0718(.A(new_n360), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n385), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n381), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n377), .B2(new_n360), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n877), .B1(new_n912), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n360), .A2(new_n377), .A3(new_n690), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT114), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n899), .B1(new_n897), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(new_n898), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n896), .B(new_n882), .C1(new_n876), .C2(new_n454), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n912), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n926), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n746), .A2(new_n481), .A3(new_n749), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n939), .A2(new_n661), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(G330), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT38), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT113), .B1(new_n892), .B2(new_n904), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n908), .B(new_n903), .C1(new_n884), .C2(new_n891), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n726), .A2(new_n728), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n715), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n823), .B1(new_n920), .B2(new_n922), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT40), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT115), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n933), .B1(new_n892), .B2(new_n904), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n952), .A2(KEYINPUT40), .A3(new_n823), .A4(new_n924), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT40), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n961), .B(new_n954), .C1(new_n715), .C2(new_n951), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(KEYINPUT115), .C1(new_n910), .C2(new_n933), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n956), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n481), .A2(new_n952), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n942), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n941), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n206), .B2(new_n752), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n941), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n875), .B1(new_n969), .B2(new_n970), .ZN(G367));
  INV_X1    g0771(.A(new_n805), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n210), .B2(new_n327), .ZN(new_n973));
  INV_X1    g0773(.A(new_n807), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n243), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n756), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n790), .A2(new_n223), .ZN(new_n977));
  INV_X1    g0777(.A(new_n768), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n267), .B1(new_n765), .B2(new_n851), .C1(new_n978), .C2(new_n850), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n977), .B(new_n979), .C1(G159), .C2(new_n786), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n771), .A2(new_n249), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n784), .A2(G143), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n280), .C2(new_n770), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n980), .B(new_n983), .C1(new_n202), .C2(new_n779), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n421), .B1(G317), .B2(new_n766), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT46), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n793), .B2(new_n491), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(new_n779), .C2(new_n840), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n790), .A2(new_n552), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G294), .B2(new_n786), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n768), .A2(G303), .B1(G311), .B2(new_n784), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT119), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT119), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n986), .A2(new_n627), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n770), .A2(new_n994), .B1(new_n772), .B2(new_n318), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n992), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n984), .B1(new_n988), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n976), .B1(new_n998), .B2(new_n762), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n576), .A2(new_n690), .ZN(new_n1000));
  MUX2_X1   g0800(.A(new_n668), .B(new_n584), .S(new_n1000), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n999), .B1(new_n1001), .B2(new_n804), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n755), .A2(new_n206), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n706), .A2(new_n703), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n740), .A2(new_n702), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n667), .B1(new_n614), .B2(new_n702), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT45), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT118), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1005), .B(new_n1009), .C1(new_n1012), .C2(KEYINPUT44), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1012), .A2(KEYINPUT44), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n699), .B(KEYINPUT99), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n701), .A2(new_n1011), .A3(new_n1016), .A4(new_n1015), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n706), .B1(new_n693), .B2(new_n705), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(new_n698), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n750), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n750), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n709), .B(KEYINPUT41), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1004), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT117), .Z(new_n1029));
  NAND3_X1  g0829(.A1(new_n537), .A2(new_n705), .A3(new_n1008), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT42), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n740), .B1(new_n533), .B2(new_n1007), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n702), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1030), .A2(KEYINPUT42), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1029), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT116), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1036), .B(new_n1038), .Z(new_n1039));
  NOR2_X1   g0839(.A1(new_n701), .A2(new_n1009), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1002), .B1(new_n1027), .B2(new_n1043), .ZN(G387));
  AOI21_X1  g0844(.A(new_n710), .B1(new_n1022), .B2(new_n750), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n750), .B2(new_n1022), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n693), .A2(new_n804), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n807), .B1(new_n240), .B2(new_n260), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n809), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n711), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n324), .A2(new_n202), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT50), .Z(new_n1052));
  AOI21_X1  g0852(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n711), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1050), .A2(new_n1054), .B1(new_n504), .B2(new_n708), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n756), .B1(new_n1055), .B2(new_n805), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n793), .A2(new_n223), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n989), .B(new_n1057), .C1(new_n784), .C2(G159), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n421), .B1(new_n850), .B2(new_n765), .C1(new_n978), .C2(new_n202), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n780), .B2(G68), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n281), .A2(new_n282), .A3(new_n786), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n564), .A2(new_n772), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n421), .B1(G326), .B2(new_n766), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n793), .A2(new_n516), .B1(new_n840), .B2(new_n771), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n784), .A2(G322), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n768), .A2(G317), .B1(G311), .B2(new_n786), .ZN(new_n1067));
  INV_X1    g0867(.A(G303), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1066), .B(new_n1067), .C1(new_n779), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1065), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1064), .B1(new_n491), .B2(new_n790), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1063), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1056), .B1(new_n1076), .B2(new_n762), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1022), .A2(new_n1004), .B1(new_n1047), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT120), .B1(new_n1046), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1046), .A2(KEYINPUT120), .A3(new_n1078), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(G393));
  NAND3_X1  g0882(.A1(new_n1019), .A2(new_n1020), .A3(new_n1004), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n972), .B1(new_n552), .B2(new_n210), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n974), .A2(new_n247), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n756), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n768), .A2(G311), .B1(G317), .B2(new_n784), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT52), .Z(new_n1088));
  AOI211_X1 g0888(.A(new_n267), .B(new_n791), .C1(G322), .C2(new_n766), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n787), .A2(new_n1068), .B1(new_n771), .B2(new_n491), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G283), .B2(new_n770), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n780), .A2(G294), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n780), .A2(new_n324), .B1(G50), .B2(new_n786), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT121), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n768), .A2(G159), .B1(G150), .B2(new_n784), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT51), .Z(new_n1097));
  NOR2_X1   g0897(.A1(new_n771), .A2(new_n223), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1098), .B(new_n846), .C1(new_n225), .C2(new_n770), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n512), .B1(G143), .B2(new_n766), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1097), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1093), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1086), .B1(new_n1102), .B2(new_n762), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1008), .B2(new_n804), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1023), .A2(new_n709), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1019), .A2(new_n1020), .B1(new_n750), .B2(new_n1022), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1083), .B(new_n1104), .C1(new_n1105), .C2(new_n1106), .ZN(G390));
  AOI21_X1  g0907(.A(new_n913), .B1(new_n824), .B2(new_n829), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n927), .B1(new_n1108), .B2(new_n923), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n935), .B(new_n1109), .C1(new_n912), .C2(new_n936), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n923), .B(KEYINPUT122), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n820), .A2(new_n822), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n745), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1111), .B1(new_n1113), .B2(new_n914), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n933), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n907), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n927), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n823), .A2(G330), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n715), .B2(new_n730), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n924), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1110), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n934), .B1(new_n948), .B2(KEYINPUT39), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n1109), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1119), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n952), .A2(new_n924), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1122), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(new_n1003), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n837), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n812), .B1(new_n1130), .B2(new_n283), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n787), .A2(new_n851), .B1(new_n771), .B2(new_n402), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n780), .B2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT124), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n770), .A2(G150), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT53), .Z(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n267), .B1(new_n765), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G132), .B2(new_n768), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n782), .A2(G50), .B1(G128), .B2(new_n784), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1135), .A2(new_n1137), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n488), .B1(new_n765), .B2(new_n516), .C1(new_n978), .C2(new_n627), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n858), .B(new_n1143), .C1(G87), .C2(new_n770), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n852), .A2(new_n840), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1098), .B(new_n1145), .C1(new_n318), .C2(new_n786), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n552), .C2(new_n779), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1131), .B1(new_n1148), .B2(new_n763), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n1124), .B2(new_n802), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1129), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1111), .B1(new_n953), .B2(new_n1119), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1152), .A2(new_n1121), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n913), .B1(new_n745), .B2(new_n1112), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1127), .B1(new_n924), .B2(new_n1120), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1153), .A2(new_n1154), .B1(new_n1155), .B2(new_n917), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT123), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n965), .B2(G330), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n662), .A2(new_n953), .A3(KEYINPUT123), .A4(new_n942), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n939), .B(new_n661), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1128), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1122), .B(new_n1161), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n709), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1151), .A2(new_n1165), .ZN(G378));
  INV_X1    g0966(.A(KEYINPUT125), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n824), .A2(new_n829), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n923), .B1(new_n1168), .B2(new_n914), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n948), .A2(new_n1169), .B1(new_n876), .B2(new_n687), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1124), .B2(new_n927), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n955), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n961), .B1(new_n912), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n942), .B1(new_n960), .B2(new_n963), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n390), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n655), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n386), .A2(new_n882), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1173), .A2(new_n1174), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1171), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1173), .A2(new_n1174), .A3(new_n1180), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1178), .B(new_n1179), .Z(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT115), .B1(new_n1116), .B2(new_n962), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n963), .ZN(new_n1187));
  OAI21_X1  g0987(.A(G330), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1185), .B1(new_n1188), .B2(new_n956), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n938), .A2(new_n1184), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1003), .B1(new_n1183), .B2(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n787), .A2(new_n552), .B1(new_n852), .B2(new_n627), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1192), .B(new_n1057), .C1(new_n280), .C2(new_n782), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n978), .A2(new_n504), .B1(new_n840), .B2(new_n765), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n512), .A2(new_n259), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1194), .A2(new_n981), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(new_n560), .C2(new_n779), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G50), .B1(new_n414), .B2(new_n259), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1197), .A2(new_n1198), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n786), .A2(G132), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n852), .B2(new_n1138), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G150), .B2(new_n772), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G128), .A2(new_n768), .B1(new_n770), .B2(new_n1133), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n851), .C2(new_n779), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n782), .A2(G159), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1200), .B1(new_n1198), .B2(new_n1197), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n762), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(new_n756), .C1(G50), .C2(new_n837), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1185), .B2(new_n802), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1167), .B1(new_n1191), .B2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1181), .A2(new_n1182), .A3(new_n1171), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n937), .A2(new_n928), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1189), .A2(new_n1184), .B1(new_n1217), .B2(new_n1170), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1004), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1214), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(KEYINPUT125), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1215), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1183), .A2(new_n1190), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1160), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1164), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1225), .A3(KEYINPUT57), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1190), .A2(new_n1183), .B1(new_n1164), .B2(new_n1224), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n709), .C1(KEYINPUT57), .C2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1222), .A2(new_n1228), .ZN(G375));
  NAND2_X1  g1029(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1162), .A2(new_n1026), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1156), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1111), .A2(new_n802), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n793), .A2(new_n552), .B1(new_n491), .B2(new_n787), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n977), .B(new_n1234), .C1(G294), .C2(new_n784), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n780), .A2(new_n318), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n488), .B1(new_n765), .B2(new_n1068), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G283), .B2(new_n768), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1062), .A3(new_n1236), .A4(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n978), .A2(new_n851), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n512), .B(new_n1240), .C1(G128), .C2(new_n766), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n780), .A2(G150), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n793), .A2(new_n402), .B1(new_n202), .B2(new_n771), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n786), .B2(new_n1133), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n782), .A2(new_n280), .B1(G132), .B2(new_n784), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1241), .A2(new_n1242), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n763), .B1(new_n1239), .B2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n812), .B(new_n1247), .C1(new_n249), .C2(new_n1130), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1232), .A2(new_n1004), .B1(new_n1233), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1231), .A2(new_n1249), .ZN(G381));
  OR4_X1    g1050(.A1(G384), .A2(G387), .A3(G390), .A4(G381), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1080), .A2(new_n815), .A3(new_n1081), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G378), .A2(new_n1251), .A3(G375), .A4(new_n1252), .ZN(G407));
  INV_X1    g1053(.A(G378), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n688), .A2(G213), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G375), .C2(new_n1257), .ZN(G409));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  INV_X1    g1059(.A(G390), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT126), .B1(G387), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1081), .ZN(new_n1262));
  OAI21_X1  g1062(.A(G396), .B1(new_n1262), .B2(new_n1079), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1252), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1025), .B1(new_n1023), .B2(new_n750), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1042), .B(new_n1041), .C1(new_n1265), .C2(new_n1004), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1266), .A2(new_n1002), .A3(G390), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G390), .B1(new_n1266), .B2(new_n1002), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1261), .A2(new_n1264), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1264), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(new_n1260), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(new_n1002), .A3(G390), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1270), .A2(KEYINPUT126), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1222), .A2(new_n1228), .A3(G378), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1227), .A2(new_n1026), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1254), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1256), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1156), .A2(new_n1160), .A3(KEYINPUT60), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n709), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1162), .A2(KEYINPUT60), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1230), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(G384), .A3(new_n1249), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1249), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n835), .B(new_n865), .C1(new_n1284), .C2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(G2897), .A3(new_n1256), .ZN(new_n1290));
  INV_X1    g1090(.A(G2897), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1286), .B(new_n1288), .C1(new_n1291), .C2(new_n1255), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1275), .B1(new_n1280), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1289), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1295), .B1(new_n1280), .B2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n1256), .B(new_n1289), .C1(new_n1276), .C2(new_n1279), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1295), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1274), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1296), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1302), .B(new_n1275), .C1(new_n1280), .C2(new_n1293), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1274), .B1(KEYINPUT63), .B2(new_n1299), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1259), .B1(new_n1301), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1294), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1280), .A2(new_n1296), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1307), .A2(new_n1310), .A3(new_n1274), .A4(new_n1302), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1312), .A2(new_n1294), .A3(new_n1297), .ZN(new_n1313));
  OAI211_X1 g1113(.A(KEYINPUT127), .B(new_n1311), .C1(new_n1313), .C2(new_n1274), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1306), .A2(new_n1314), .ZN(G405));
  NAND2_X1  g1115(.A1(G375), .A2(new_n1254), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1276), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1317), .B(new_n1289), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1318), .B(new_n1274), .ZN(G402));
endmodule


