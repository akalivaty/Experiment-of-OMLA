//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND3_X1  g0012(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n212), .B1(new_n213), .B2(new_n216), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1698), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G226), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G97), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n247), .A2(new_n248), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  INV_X1    g0053(.A(G232), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n250), .B(new_n251), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(G1), .B(G13), .C1(new_n246), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n206), .A2(G274), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT68), .B(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n266), .B2(G238), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n259), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n259), .B2(new_n267), .ZN(new_n271));
  OAI21_X1  g0071(.A(G200), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n259), .A2(new_n267), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  OAI211_X1 g0075(.A(G190), .B(new_n269), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G1), .A2(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n246), .A2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G77), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G68), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n283), .A2(G50), .B1(G20), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n280), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT72), .B(KEYINPUT11), .Z(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G20), .A3(new_n284), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT12), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n290), .A2(new_n207), .A3(G1), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n279), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n207), .A2(KEYINPUT69), .A3(G1), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT69), .B1(new_n207), .B2(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n300), .A2(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n272), .A2(new_n276), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(G169), .B1(new_n270), .B2(new_n271), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT14), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(G169), .C1(new_n270), .C2(new_n271), .ZN(new_n308));
  OAI211_X1 g0108(.A(G179), .B(new_n269), .C1(new_n274), .C2(new_n275), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n302), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(KEYINPUT73), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n275), .B1(new_n259), .B2(new_n267), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n270), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(KEYINPUT14), .B2(new_n305), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n302), .B1(new_n317), .B2(new_n308), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT73), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n318), .A2(new_n319), .A3(new_n304), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n299), .A2(new_n322), .ZN(new_n323));
  AOI211_X1 g0123(.A(new_n279), .B(new_n295), .C1(new_n323), .C2(KEYINPUT76), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(new_n295), .B2(new_n321), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT7), .B1(new_n330), .B2(new_n207), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  NOR4_X1   g0132(.A1(new_n328), .A2(new_n329), .A3(new_n332), .A4(G20), .ZN(new_n333));
  OAI21_X1  g0133(.A(G68), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT74), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G58), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n284), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n338), .B2(new_n201), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n283), .A2(G159), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT74), .B(G68), .C1(new_n331), .C2(new_n333), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n336), .A2(KEYINPUT16), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT75), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n247), .A2(new_n207), .A3(new_n248), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n332), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n248), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n284), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n341), .B1(new_n350), .B2(KEYINPUT74), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n351), .A2(new_n336), .A3(KEYINPUT75), .A4(KEYINPUT16), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n280), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT16), .B1(new_n334), .B2(new_n342), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n327), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n249), .A2(G223), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  INV_X1    g0158(.A(G226), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n357), .B(new_n358), .C1(new_n253), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n258), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n263), .B1(new_n266), .B2(G232), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G179), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n363), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT18), .B1(new_n356), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT18), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n354), .B(new_n280), .C1(new_n346), .C2(new_n352), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n369), .B(new_n366), .C1(new_n370), .C2(new_n327), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n361), .A2(new_n373), .A3(new_n362), .ZN(new_n374));
  AOI21_X1  g0174(.A(G200), .B1(new_n361), .B2(new_n362), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n326), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n372), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n343), .A2(new_n342), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n350), .A2(KEYINPUT74), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT75), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n381));
  INV_X1    g0181(.A(new_n352), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n355), .B(new_n279), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n376), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(KEYINPUT17), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n368), .A2(new_n371), .A3(new_n377), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n295), .A2(G50), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n300), .B2(G50), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n322), .A2(new_n281), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n283), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n280), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT9), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT10), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n261), .A2(new_n262), .ZN(new_n396));
  INV_X1    g0196(.A(new_n260), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n359), .B2(new_n265), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n249), .A2(G222), .B1(new_n330), .B2(G77), .ZN(new_n400));
  INV_X1    g0200(.A(G223), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n253), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n402), .B2(new_n258), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G190), .ZN(new_n404));
  INV_X1    g0204(.A(G200), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n394), .A2(new_n395), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n404), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT10), .B1(new_n408), .B2(new_n393), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n403), .A2(G179), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n365), .B2(new_n403), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n391), .B2(new_n388), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n249), .A2(G232), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n252), .A2(G238), .A3(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n330), .A2(G107), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n258), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n257), .A2(G244), .A3(new_n264), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n398), .A2(KEYINPUT70), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT70), .B1(new_n398), .B2(new_n419), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n373), .B(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n398), .A2(new_n419), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT70), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n420), .B1(new_n258), .B2(new_n417), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n423), .B1(new_n427), .B2(G200), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n322), .A2(new_n283), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n280), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G77), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n295), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n300), .B2(new_n434), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(G179), .B(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n427), .B2(new_n365), .ZN(new_n440));
  INV_X1    g0240(.A(new_n437), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n410), .A2(new_n413), .A3(new_n443), .ZN(new_n444));
  NOR4_X1   g0244(.A1(new_n313), .A2(new_n320), .A3(new_n386), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT21), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n291), .A2(G20), .ZN(new_n447));
  INV_X1    g0247(.A(G116), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n206), .A2(G33), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n280), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n452), .B2(new_n448), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n246), .A2(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  AOI21_X1  g0255(.A(G20), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n207), .A2(new_n448), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n279), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT20), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT20), .B(new_n279), .C1(new_n456), .C2(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n365), .B1(new_n453), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n252), .A2(G264), .A3(G1698), .ZN(new_n464));
  INV_X1    g0264(.A(G1698), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n252), .A2(G257), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G303), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n464), .B(new_n466), .C1(new_n467), .C2(new_n252), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n258), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n206), .B(G45), .C1(new_n470), .C2(G41), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(KEYINPUT5), .B2(new_n261), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(KEYINPUT81), .A3(G270), .A4(new_n257), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(G274), .C1(KEYINPUT5), .C2(new_n261), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT68), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G41), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT5), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G270), .B(new_n257), .C1(new_n479), .C2(new_n471), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n469), .A2(new_n474), .A3(new_n475), .A4(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n463), .A2(new_n483), .A3(KEYINPUT83), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT83), .B1(new_n463), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n446), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n483), .A2(new_n314), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n453), .A2(new_n462), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n463), .A2(new_n483), .A3(KEYINPUT21), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n463), .A2(new_n483), .A3(KEYINPUT82), .A4(KEYINPUT21), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n483), .A2(new_n405), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G190), .B2(new_n483), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n488), .ZN(new_n497));
  AND4_X1   g0297(.A1(new_n486), .A2(new_n489), .A3(new_n494), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n291), .A2(G20), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n500), .A2(KEYINPUT25), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(KEYINPUT25), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n502), .C1(new_n499), .C2(new_n451), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT23), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n207), .B2(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n499), .A2(KEYINPUT23), .A3(G20), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n246), .A2(new_n448), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n207), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n252), .A2(new_n207), .A3(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT22), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT22), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n252), .A2(new_n512), .A3(new_n207), .A4(G87), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n514), .A2(KEYINPUT24), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n280), .B1(new_n514), .B2(KEYINPUT24), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n503), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n479), .A2(new_n471), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n258), .ZN(new_n520));
  OAI211_X1 g0320(.A(G250), .B(new_n465), .C1(new_n328), .C2(new_n329), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n522));
  INV_X1    g0322(.A(G294), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n246), .C2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n520), .A2(G264), .B1(new_n258), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G179), .A3(new_n475), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT84), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n258), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n473), .A2(G264), .A3(new_n257), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n475), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n526), .A2(new_n527), .B1(G169), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n530), .A2(new_n527), .A3(G169), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n518), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n525), .A2(KEYINPUT85), .A3(new_n373), .A4(new_n475), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT85), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n530), .B2(new_n405), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n530), .A2(G190), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n517), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n397), .A2(G45), .ZN(new_n541));
  OAI21_X1  g0341(.A(G250), .B1(new_n262), .B2(G1), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n257), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G244), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n544));
  OAI211_X1 g0344(.A(G238), .B(new_n465), .C1(new_n328), .C2(new_n329), .ZN(new_n545));
  INV_X1    g0345(.A(new_n507), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n547), .A2(KEYINPUT79), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT79), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n544), .A2(new_n545), .A3(new_n549), .A4(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n258), .ZN(new_n551));
  OAI211_X1 g0351(.A(G200), .B(new_n543), .C1(new_n548), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n452), .A2(G87), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n207), .B1(new_n251), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(G87), .A2(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n499), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n207), .B(G68), .C1(new_n328), .C2(new_n329), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n554), .B1(new_n251), .B2(G20), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n279), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n430), .A2(new_n447), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n553), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n543), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n550), .A2(new_n258), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n547), .A2(KEYINPUT79), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n552), .B(new_n565), .C1(new_n569), .C2(new_n373), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n451), .A2(G97), .ZN(new_n571));
  INV_X1    g0371(.A(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n447), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT78), .ZN(new_n575));
  OAI21_X1  g0375(.A(G107), .B1(new_n331), .B2(new_n333), .ZN(new_n576));
  XNOR2_X1  g0376(.A(G97), .B(G107), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n499), .A2(KEYINPUT6), .A3(G97), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G20), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n283), .A2(KEYINPUT77), .A3(G77), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT77), .B1(new_n283), .B2(G77), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n576), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n575), .B1(new_n587), .B2(new_n279), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n580), .B1(new_n577), .B2(new_n578), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n589), .B2(new_n207), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n499), .B1(new_n348), .B2(new_n349), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n575), .B(new_n279), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n574), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n252), .B2(G250), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n465), .ZN(new_n597));
  OAI21_X1  g0397(.A(G244), .B1(new_n328), .B2(new_n329), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n595), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n595), .A2(G1698), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(G244), .C1(new_n329), .C2(new_n328), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n455), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n258), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(G257), .B(new_n257), .C1(new_n479), .C2(new_n471), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n475), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(G179), .A3(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n598), .A2(new_n595), .B1(G33), .B2(G283), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n608), .B(new_n601), .C1(new_n465), .C2(new_n596), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n605), .B1(new_n609), .B2(new_n258), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n607), .B1(new_n610), .B2(new_n365), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n594), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n279), .B1(new_n590), .B2(new_n591), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT78), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n614), .A2(new_n592), .B1(new_n573), .B2(new_n571), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n603), .A2(new_n373), .A3(new_n606), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n610), .B2(G200), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n543), .B1(new_n548), .B2(new_n551), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n314), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n365), .B(new_n543), .C1(new_n548), .C2(new_n551), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n296), .A2(new_n430), .A3(new_n450), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n562), .A2(new_n564), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT80), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n562), .A2(KEYINPUT80), .A3(new_n564), .A4(new_n622), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n620), .A2(new_n621), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n570), .A2(new_n612), .A3(new_n618), .A4(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n445), .A2(new_n498), .A3(new_n540), .A4(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n310), .A2(new_n311), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n304), .B1(new_n630), .B2(new_n442), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n377), .A3(new_n385), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n368), .A2(new_n371), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT89), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n632), .A2(KEYINPUT89), .A3(new_n633), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n410), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n612), .A2(new_n618), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n621), .B(new_n623), .C1(new_n569), .C2(G179), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n570), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n639), .A2(new_n640), .A3(new_n539), .A4(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n642), .A2(new_n539), .A3(new_n618), .A4(new_n612), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT86), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n533), .A2(new_n489), .A3(new_n486), .A4(new_n494), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n570), .A2(new_n641), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n603), .A2(G179), .A3(new_n606), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n365), .B1(new_n603), .B2(new_n606), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT88), .B1(new_n651), .B2(new_n615), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT88), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n594), .A2(new_n653), .A3(new_n611), .ZN(new_n654));
  AOI211_X1 g0454(.A(KEYINPUT26), .B(new_n648), .C1(new_n652), .C2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n627), .A2(new_n594), .A3(new_n570), .A4(new_n611), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n641), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n647), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n445), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n638), .A2(new_n413), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT90), .ZN(G369));
  INV_X1    g0465(.A(new_n498), .ZN(new_n666));
  INV_X1    g0466(.A(new_n291), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .A3(G20), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT27), .B1(new_n667), .B2(G20), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n488), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n489), .A2(new_n486), .A3(new_n494), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n517), .A2(new_n673), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT91), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n540), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n533), .B2(new_n673), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n676), .A2(new_n673), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n540), .A3(new_n682), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n533), .A2(new_n672), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT92), .Z(G399));
  INV_X1    g0492(.A(new_n210), .ZN(new_n693));
  INV_X1    g0493(.A(new_n261), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n556), .A2(new_n499), .A3(new_n448), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n216), .B2(new_n696), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  INV_X1    g0501(.A(new_n610), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n487), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n619), .A2(new_n525), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT93), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n704), .A2(KEYINPUT93), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n610), .B1(new_n475), .B2(new_n525), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n314), .A3(new_n483), .A4(new_n569), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n707), .B2(new_n708), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n672), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n498), .A2(new_n540), .A3(new_n628), .A4(new_n673), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n714), .A3(KEYINPUT31), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(new_n672), .C1(new_n709), .C2(new_n712), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n715), .A2(G330), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n672), .B1(new_n647), .B2(new_n661), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n656), .A2(KEYINPUT26), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT26), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n648), .B1(new_n652), .B2(new_n654), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n721), .B(new_n659), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n489), .A2(new_n486), .A3(new_n494), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n644), .B1(new_n725), .B2(new_n533), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT29), .B(new_n673), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n718), .B1(new_n720), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n701), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n290), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n206), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n695), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n678), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n736), .B2(new_n680), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n207), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT95), .Z(new_n740));
  NOR2_X1   g0540(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n740), .ZN(new_n742));
  OR2_X1    g0542(.A1(KEYINPUT96), .A2(G169), .ZN(new_n743));
  NAND2_X1  g0543(.A1(KEYINPUT96), .A2(G169), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n207), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n278), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n210), .A2(new_n252), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT94), .ZN(new_n749));
  INV_X1    g0549(.A(G355), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n749), .A2(new_n750), .B1(G116), .B2(new_n210), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n693), .A2(new_n252), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n243), .A2(G45), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n216), .A2(new_n262), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n747), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  NOR2_X1   g0558(.A1(new_n314), .A2(new_n405), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n207), .A2(G190), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n330), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n207), .A2(new_n373), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n759), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n314), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n765), .A2(G326), .B1(new_n768), .B2(G311), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n763), .A2(new_n766), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n405), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n760), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G322), .A2(new_n771), .B1(new_n774), .B2(G283), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n373), .A2(G179), .A3(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n207), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n762), .B(new_n776), .C1(G294), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n763), .A2(new_n772), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n760), .A2(new_n314), .A3(new_n405), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n786), .A2(G303), .B1(G329), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  INV_X1    g0595(.A(new_n761), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G50), .A2(new_n765), .B1(new_n796), .B2(G68), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n779), .A2(G97), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n330), .B1(new_n768), .B2(G77), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n773), .A2(new_n499), .ZN(new_n801));
  INV_X1    g0601(.A(G87), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n337), .A2(new_n770), .B1(new_n781), .B2(new_n802), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n780), .A2(new_n792), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n746), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n757), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n733), .B1(new_n741), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n737), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NOR2_X1   g0610(.A1(new_n442), .A2(new_n673), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n441), .A2(new_n672), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n438), .A2(new_n442), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT101), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT101), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n438), .A2(new_n442), .A3(new_n815), .A4(new_n812), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n811), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n719), .A2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n672), .B(new_n817), .C1(new_n647), .C2(new_n661), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n733), .B1(new_n821), .B2(new_n718), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n718), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n746), .A2(new_n738), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n734), .B1(new_n824), .B2(new_n434), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G143), .A2(new_n771), .B1(new_n796), .B2(G150), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n765), .A2(G137), .B1(new_n768), .B2(G159), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n779), .A2(G58), .B1(new_n774), .B2(G68), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n785), .B2(new_n202), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n252), .B1(new_n790), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT100), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n330), .B1(new_n785), .B2(new_n499), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT99), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n796), .A2(G283), .B1(new_n774), .B2(G87), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n467), .B2(new_n764), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n798), .B1(new_n448), .B2(new_n767), .C1(new_n523), .C2(new_n770), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n840), .B(new_n841), .C1(G311), .C2(new_n791), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n833), .A2(new_n836), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n738), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n825), .B1(new_n806), .B2(new_n843), .C1(new_n818), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n823), .A2(new_n845), .ZN(G384));
  INV_X1    g0646(.A(KEYINPUT35), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n448), .B(new_n213), .C1(new_n589), .C2(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n848), .A2(KEYINPUT102), .B1(new_n847), .B2(new_n589), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(KEYINPUT102), .B2(new_n848), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT36), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n215), .B(G77), .C1(new_n337), .C2(new_n284), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n202), .A2(G68), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n206), .B(G13), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT40), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n383), .A2(new_n384), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n380), .A2(KEYINPUT16), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n327), .B1(new_n353), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n857), .B1(new_n859), .B2(new_n670), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n367), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n670), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n370), .A2(new_n327), .B1(new_n366), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n857), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n859), .A2(new_n670), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n386), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT108), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT108), .A4(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n386), .B(new_n863), .C1(new_n370), .C2(new_n327), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT106), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n876), .B(new_n376), .C1(new_n353), .C2(new_n355), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT106), .B1(new_n383), .B2(new_n384), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n864), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT107), .A3(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n866), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT107), .B1(new_n879), .B2(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n875), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n715), .A2(new_n717), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n311), .A2(new_n672), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n630), .A2(new_n303), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT104), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n312), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n630), .A2(KEYINPUT105), .A3(new_n673), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n318), .B2(new_n672), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n817), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n887), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT109), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n856), .B1(new_n886), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n867), .A2(new_n869), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n884), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n870), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n856), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n856), .A2(KEYINPUT109), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n887), .A2(new_n445), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n679), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n874), .A2(new_n885), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n903), .B2(new_n870), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n630), .A2(new_n672), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n633), .A2(new_n863), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n893), .A2(new_n897), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT103), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n442), .A2(new_n672), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n922), .B1(new_n820), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n662), .A2(new_n673), .A3(new_n818), .ZN(new_n925));
  INV_X1    g0725(.A(new_n923), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(KEYINPUT103), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n921), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n919), .B1(new_n928), .B2(new_n904), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n918), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n720), .A2(new_n445), .A3(new_n727), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n931), .A2(new_n413), .A3(new_n638), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n911), .A2(new_n933), .B1(new_n206), .B2(new_n730), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n911), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n855), .B1(new_n934), .B2(new_n935), .ZN(G367));
  OAI21_X1  g0736(.A(new_n639), .B1(new_n615), .B2(new_n673), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n612), .B2(new_n673), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT110), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(new_n533), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n672), .B1(new_n940), .B2(new_n612), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n688), .A2(new_n937), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT42), .Z(new_n943));
  INV_X1    g0743(.A(KEYINPUT43), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n673), .A2(new_n565), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n659), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n642), .B2(new_n945), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n941), .A2(new_n943), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n944), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n685), .ZN(new_n951));
  INV_X1    g0751(.A(new_n939), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n950), .B(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n695), .B(KEYINPUT41), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n688), .B1(new_n684), .B2(new_n687), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n680), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n690), .A2(new_n938), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT45), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n690), .A2(new_n938), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT44), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(KEYINPUT111), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT112), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n685), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n959), .A2(new_n961), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT111), .B1(new_n951), .B2(KEYINPUT112), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n728), .B(new_n957), .C1(new_n964), .C2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n955), .B1(new_n968), .B2(new_n728), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n954), .B1(new_n969), .B2(new_n732), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n753), .A2(new_n234), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n747), .B1(new_n210), .B2(new_n429), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G150), .A2(new_n771), .B1(new_n768), .B2(G50), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT113), .B(G137), .Z(new_n974));
  OAI221_X1 g0774(.A(new_n973), .B1(new_n793), .B2(new_n761), .C1(new_n790), .C2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n778), .A2(new_n284), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n330), .B1(new_n782), .B2(G58), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n765), .A2(G143), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(new_n434), .C2(new_n773), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n975), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT114), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G294), .A2(new_n796), .B1(new_n771), .B2(G303), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n774), .A2(G97), .ZN(new_n983));
  INV_X1    g0783(.A(G311), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n983), .C1(new_n984), .C2(new_n764), .ZN(new_n985));
  AND2_X1   g0785(.A1(KEYINPUT46), .A2(G116), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n985), .B1(new_n786), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(G283), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n330), .B1(new_n767), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT46), .B1(new_n782), .B2(G116), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(G107), .C2(new_n779), .ZN(new_n991));
  INV_X1    g0791(.A(G317), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n987), .B(new_n991), .C1(new_n992), .C2(new_n790), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n981), .A2(KEYINPUT47), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n746), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT47), .B1(new_n981), .B2(new_n993), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n733), .B1(new_n971), .B2(new_n972), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n947), .B2(new_n742), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT115), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n970), .A2(new_n999), .ZN(G387));
  NAND2_X1  g0800(.A1(new_n957), .A2(new_n732), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n684), .A2(new_n740), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n330), .B1(new_n773), .B2(new_n448), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n779), .A2(G283), .B1(new_n782), .B2(G294), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n765), .A2(G322), .B1(new_n768), .B2(G303), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n984), .B2(new_n761), .C1(new_n992), .C2(new_n770), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT49), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1003), .B(new_n1010), .C1(G326), .C2(new_n791), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G159), .A2(new_n765), .B1(new_n782), .B2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n202), .B2(new_n770), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n796), .A2(new_n322), .B1(new_n768), .B2(G68), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n779), .A2(new_n430), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1014), .A2(new_n252), .A3(new_n983), .A4(new_n1015), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1013), .B(new_n1016), .C1(G150), .C2(new_n791), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n746), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n321), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  AOI211_X1 g0820(.A(G45), .B(new_n697), .C1(G68), .C2(G77), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n753), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT116), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n231), .B2(new_n262), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(G107), .B2(new_n210), .C1(new_n698), .C2(new_n749), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n734), .B1(new_n1025), .B2(new_n747), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n728), .A2(new_n957), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n695), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n728), .A2(new_n957), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1001), .B1(new_n1002), .B2(new_n1027), .C1(new_n1029), .C2(new_n1030), .ZN(G393));
  OAI21_X1  g0831(.A(new_n747), .B1(new_n572), .B2(new_n210), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n240), .B2(new_n752), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n791), .A2(G322), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n988), .A2(new_n781), .B1(new_n761), .B2(new_n467), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G294), .B2(new_n768), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n252), .B(new_n801), .C1(G116), .C2(new_n779), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n764), .A2(new_n992), .B1(new_n770), .B2(new_n984), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT52), .Z(new_n1040));
  OAI22_X1  g0840(.A1(new_n202), .A2(new_n761), .B1(new_n781), .B2(new_n284), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n322), .B2(new_n768), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n252), .B1(new_n773), .B2(new_n802), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G77), .B2(new_n779), .ZN(new_n1044));
  INV_X1    g0844(.A(G143), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1042), .B(new_n1044), .C1(new_n1045), .C2(new_n790), .ZN(new_n1046));
  INV_X1    g0846(.A(G150), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n764), .A2(new_n1047), .B1(new_n770), .B2(new_n793), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT51), .Z(new_n1049));
  OAI22_X1  g0849(.A1(new_n1038), .A2(new_n1040), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n734), .B(new_n1033), .C1(new_n746), .C2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n952), .B2(new_n740), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n965), .B(new_n951), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n731), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n696), .B1(new_n1053), .B2(new_n1028), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1054), .B1(new_n968), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(G390));
  INV_X1    g0857(.A(new_n824), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n330), .B1(new_n773), .B2(new_n284), .C1(new_n778), .C2(new_n434), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n499), .A2(new_n761), .B1(new_n770), .B2(new_n448), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n764), .A2(new_n988), .B1(new_n767), .B2(new_n572), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n802), .B2(new_n785), .C1(new_n523), .C2(new_n790), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT118), .Z(new_n1064));
  OAI221_X1 g0864(.A(new_n252), .B1(new_n974), .B2(new_n761), .C1(new_n793), .C2(new_n778), .ZN(new_n1065));
  INV_X1    g0865(.A(G128), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT54), .B(G143), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n764), .A2(new_n1066), .B1(new_n767), .B2(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n770), .A2(new_n834), .B1(new_n773), .B2(new_n202), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1065), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n781), .A2(new_n1047), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT53), .ZN(new_n1072));
  INV_X1    g0872(.A(G125), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1070), .B(new_n1072), .C1(new_n1073), .C2(new_n790), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1064), .A2(KEYINPUT119), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n746), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT119), .B1(new_n1064), .B2(new_n1074), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n733), .B1(new_n322), .B2(new_n1058), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n872), .A2(new_n873), .B1(new_n883), .B2(new_n884), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n914), .B1(new_n1079), .B2(new_n912), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n1080), .B2(new_n738), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n913), .B(new_n915), .C1(new_n928), .C2(new_n917), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n917), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n673), .B1(new_n724), .B2(new_n726), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n814), .A2(new_n816), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n926), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n920), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n886), .A2(new_n1083), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1082), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n718), .A2(new_n898), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT117), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1087), .A2(new_n1083), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1079), .A2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n820), .A2(new_n922), .A3(new_n923), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT103), .B1(new_n925), .B2(new_n926), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n920), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1083), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1095), .B1(new_n1080), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1093), .B1(new_n1100), .B2(new_n1090), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1089), .A2(KEYINPUT117), .A3(new_n1091), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1092), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1081), .B1(new_n1103), .B2(new_n732), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n887), .A2(new_n445), .A3(G330), .ZN(new_n1105));
  AND4_X1   g0905(.A1(new_n413), .A2(new_n931), .A3(new_n1105), .A4(new_n638), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n715), .A2(G330), .A3(new_n717), .A4(new_n818), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n921), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1090), .A2(new_n1108), .A3(new_n1086), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1090), .A2(new_n1108), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1106), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n695), .B1(new_n1103), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1100), .A2(new_n1090), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT117), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1093), .B(new_n1090), .C1(new_n1082), .C2(new_n1088), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n1114), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1104), .B1(new_n1115), .B2(new_n1120), .ZN(G378));
  OAI21_X1  g0921(.A(G330), .B1(new_n901), .B2(new_n907), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n903), .A2(new_n870), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1098), .A2(new_n1124), .B1(new_n633), .B2(new_n863), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1083), .B1(new_n913), .B2(new_n915), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n410), .A2(new_n413), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n392), .A2(new_n670), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1130));
  XNOR2_X1  g0930(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1125), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1131), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n918), .B2(new_n929), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1123), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n918), .A2(new_n929), .A3(new_n1133), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1131), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n1122), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n732), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n733), .B1(new_n1058), .B2(G50), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n694), .A2(new_n252), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G50), .B(new_n1142), .C1(new_n246), .C2(new_n256), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT120), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G107), .A2(new_n771), .B1(new_n768), .B2(new_n430), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1142), .B(new_n1145), .C1(new_n790), .C2(new_n988), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n434), .A2(new_n781), .B1(new_n761), .B2(new_n572), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n764), .A2(new_n448), .B1(new_n773), .B2(new_n337), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1146), .A2(new_n976), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1144), .B1(KEYINPUT58), .B2(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n764), .A2(new_n1073), .B1(new_n761), .B2(new_n834), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n768), .A2(G137), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n1066), .B2(new_n770), .C1(new_n781), .C2(new_n1067), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(G150), .C2(new_n779), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n791), .A2(G124), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G33), .B(G41), .C1(new_n774), .C2(G159), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT59), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1158), .C1(new_n1154), .C2(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1150), .B1(KEYINPUT58), .B2(new_n1149), .C1(new_n1156), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1141), .B1(new_n1161), .B2(new_n746), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1131), .B2(new_n844), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1140), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n932), .A2(new_n1105), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1103), .B2(new_n1114), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1138), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1122), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT57), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n695), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1119), .A2(new_n1106), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT57), .B1(new_n1171), .B2(new_n1139), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1164), .B1(new_n1170), .B2(new_n1172), .ZN(G375));
  NAND3_X1  g0973(.A1(new_n1112), .A2(new_n732), .A3(new_n1109), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n733), .B1(new_n1058), .B2(G68), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n770), .A2(new_n974), .B1(new_n764), .B2(new_n834), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n761), .A2(new_n1067), .B1(new_n767), .B2(new_n1047), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n330), .B1(new_n774), .B2(G58), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(new_n202), .C2(new_n778), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n785), .A2(new_n793), .B1(new_n1066), .B2(new_n790), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n785), .A2(new_n572), .B1(new_n467), .B2(new_n790), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G116), .A2(new_n796), .B1(new_n771), .B2(G283), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n765), .A2(G294), .B1(new_n768), .B2(G107), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n252), .B1(new_n774), .B2(G77), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1015), .A4(new_n1185), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n1180), .A2(new_n1181), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1175), .B1(new_n1187), .B2(new_n746), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n920), .B2(new_n844), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT121), .B1(new_n1174), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1174), .A2(KEYINPUT121), .A3(new_n1189), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1112), .A2(new_n1109), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1165), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n955), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1113), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT122), .ZN(G381));
  NAND3_X1  g0999(.A1(new_n970), .A2(new_n999), .A3(new_n1056), .ZN(new_n1200));
  OR2_X1    g1000(.A1(G393), .A2(G396), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1200), .A2(G381), .A3(G384), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1081), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(new_n1204), .B2(new_n731), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n696), .B1(new_n1204), .B2(new_n1113), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n1119), .ZN(new_n1207));
  AND2_X1   g1007(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1202), .B(new_n1207), .C1(new_n1208), .C2(new_n1209), .ZN(G407));
  NAND2_X1  g1010(.A1(new_n671), .A2(G213), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1207), .B(new_n1212), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(G407), .A2(new_n1213), .A3(G213), .ZN(G409));
  INV_X1    g1014(.A(G384), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1113), .A2(new_n695), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1195), .A2(KEYINPUT60), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT60), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1194), .A2(new_n1165), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1216), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1174), .A2(KEYINPUT121), .A3(new_n1189), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(new_n1190), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1215), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1194), .A2(new_n1165), .A3(new_n1218), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1218), .B1(new_n1194), .B2(new_n1165), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n695), .B(new_n1113), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1193), .A3(G384), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT124), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1223), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT125), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT125), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1223), .A2(new_n1227), .A3(new_n1228), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1227), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G384), .B1(new_n1226), .B2(new_n1193), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT124), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1212), .A2(G2897), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1233), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1230), .A2(new_n1236), .A3(new_n1237), .A4(new_n1232), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G378), .B(new_n1164), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1171), .A2(new_n1196), .A3(new_n1139), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1140), .A2(new_n1163), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1207), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1212), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT63), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1211), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1246), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(new_n809), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n970), .A2(new_n999), .A3(new_n1056), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1056), .B1(new_n970), .B2(new_n999), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(G390), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1254), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1200), .A3(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .A4(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1252), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1250), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1246), .A2(new_n1264), .A3(new_n1265), .A4(new_n1249), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1263), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1262), .B1(new_n1271), .B2(new_n1261), .ZN(G405));
  NAND2_X1  g1072(.A1(G375), .A2(new_n1207), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1242), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1235), .B2(new_n1234), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(new_n1249), .A3(new_n1242), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1261), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1275), .A2(new_n1261), .A3(KEYINPUT127), .A4(new_n1276), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1261), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1279), .A2(new_n1280), .A3(new_n1283), .ZN(G402));
endmodule


