

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U322 ( .A(n299), .B(n298), .Z(n290) );
  XNOR2_X1 U323 ( .A(n364), .B(KEYINPUT67), .ZN(n365) );
  XNOR2_X1 U324 ( .A(n366), .B(n365), .ZN(n368) );
  INV_X1 U325 ( .A(KEYINPUT114), .ZN(n369) );
  XNOR2_X1 U326 ( .A(n300), .B(n290), .ZN(n301) );
  XNOR2_X1 U327 ( .A(n302), .B(n301), .ZN(n308) );
  XNOR2_X1 U328 ( .A(n452), .B(KEYINPUT58), .ZN(n453) );
  XNOR2_X1 U329 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  INV_X1 U330 ( .A(KEYINPUT80), .ZN(n309) );
  XNOR2_X1 U331 ( .A(G36GAT), .B(G190GAT), .ZN(n291) );
  XNOR2_X1 U332 ( .A(n291), .B(G218GAT), .ZN(n376) );
  INV_X1 U333 ( .A(KEYINPUT68), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n376), .B(n292), .ZN(n294) );
  XOR2_X1 U335 ( .A(G50GAT), .B(G162GAT), .Z(n427) );
  XNOR2_X1 U336 ( .A(G134GAT), .B(n427), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n302) );
  XOR2_X1 U338 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n296) );
  XNOR2_X1 U339 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n297), .B(KEYINPUT65), .ZN(n300) );
  XOR2_X1 U342 ( .A(KEYINPUT69), .B(KEYINPUT9), .Z(n299) );
  NAND2_X1 U343 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XOR2_X1 U344 ( .A(G29GAT), .B(G43GAT), .Z(n304) );
  XNOR2_X1 U345 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n315) );
  XOR2_X1 U347 ( .A(G85GAT), .B(G92GAT), .Z(n306) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G106GAT), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n306), .B(n305), .ZN(n332) );
  XNOR2_X1 U350 ( .A(n315), .B(n332), .ZN(n307) );
  XNOR2_X1 U351 ( .A(n308), .B(n307), .ZN(n557) );
  XNOR2_X1 U352 ( .A(n309), .B(n557), .ZN(n542) );
  XOR2_X1 U353 ( .A(KEYINPUT75), .B(G113GAT), .Z(n311) );
  XNOR2_X1 U354 ( .A(G36GAT), .B(G50GAT), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U356 ( .A(n312), .B(G197GAT), .Z(n314) );
  XOR2_X1 U357 ( .A(G141GAT), .B(G22GAT), .Z(n423) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(n423), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n319) );
  XOR2_X1 U360 ( .A(n315), .B(KEYINPUT70), .Z(n317) );
  NAND2_X1 U361 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U363 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U364 ( .A(KEYINPUT73), .B(G15GAT), .Z(n321) );
  XNOR2_X1 U365 ( .A(G8GAT), .B(G1GAT), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT74), .B(n322), .Z(n358) );
  XOR2_X1 U368 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n324) );
  XNOR2_X1 U369 ( .A(KEYINPUT72), .B(KEYINPUT29), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U371 ( .A(n358), .B(n325), .ZN(n326) );
  XOR2_X1 U372 ( .A(n327), .B(n326), .Z(n498) );
  INV_X1 U373 ( .A(n498), .ZN(n570) );
  XOR2_X1 U374 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XOR2_X1 U375 ( .A(KEYINPUT13), .B(G57GAT), .Z(n344) );
  XNOR2_X1 U376 ( .A(n437), .B(n344), .ZN(n339) );
  XOR2_X1 U377 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n329) );
  NAND2_X1 U378 ( .A1(G230GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U380 ( .A(n330), .B(KEYINPUT76), .Z(n334) );
  XNOR2_X1 U381 ( .A(G78GAT), .B(KEYINPUT77), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n331), .B(G148GAT), .ZN(n426) );
  XNOR2_X1 U383 ( .A(n426), .B(n332), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U385 ( .A(G176GAT), .B(G64GAT), .Z(n375) );
  XOR2_X1 U386 ( .A(n335), .B(n375), .Z(n337) );
  XNOR2_X1 U387 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U389 ( .A(n339), .B(n338), .Z(n574) );
  XOR2_X1 U390 ( .A(KEYINPUT41), .B(n574), .Z(n497) );
  NOR2_X1 U391 ( .A1(n570), .A2(n497), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n340), .B(KEYINPUT46), .ZN(n341) );
  NOR2_X1 U393 ( .A1(n557), .A2(n341), .ZN(n361) );
  XOR2_X1 U394 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n343) );
  XNOR2_X1 U395 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U397 ( .A(KEYINPUT12), .B(n344), .Z(n346) );
  XNOR2_X1 U398 ( .A(G22GAT), .B(G211GAT), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U400 ( .A(n348), .B(n347), .Z(n350) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U403 ( .A(G78GAT), .B(G155GAT), .Z(n352) );
  XNOR2_X1 U404 ( .A(G183GAT), .B(G71GAT), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U406 ( .A(n354), .B(n353), .Z(n360) );
  XOR2_X1 U407 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n356) );
  XNOR2_X1 U408 ( .A(G127GAT), .B(G64GAT), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U411 ( .A(n360), .B(n359), .Z(n467) );
  INV_X1 U412 ( .A(n467), .ZN(n579) );
  NAND2_X1 U413 ( .A1(n361), .A2(n579), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n362), .B(KEYINPUT113), .ZN(n363) );
  XNOR2_X1 U415 ( .A(KEYINPUT47), .B(n363), .ZN(n372) );
  XNOR2_X1 U416 ( .A(KEYINPUT36), .B(n542), .ZN(n482) );
  NOR2_X1 U417 ( .A1(n579), .A2(n482), .ZN(n366) );
  INV_X1 U418 ( .A(KEYINPUT45), .ZN(n364) );
  INV_X1 U419 ( .A(n574), .ZN(n471) );
  NOR2_X1 U420 ( .A1(n471), .A2(n498), .ZN(n367) );
  AND2_X1 U421 ( .A1(n368), .A2(n367), .ZN(n370) );
  XNOR2_X1 U422 ( .A(n370), .B(n369), .ZN(n371) );
  NAND2_X1 U423 ( .A1(n372), .A2(n371), .ZN(n374) );
  XNOR2_X1 U424 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n529) );
  XOR2_X1 U426 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U427 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U428 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U429 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n380) );
  XNOR2_X1 U430 ( .A(G8GAT), .B(G92GAT), .ZN(n379) );
  XNOR2_X1 U431 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U432 ( .A(n382), .B(n381), .Z(n392) );
  XNOR2_X1 U433 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n383) );
  XNOR2_X1 U434 ( .A(n383), .B(KEYINPUT18), .ZN(n384) );
  XOR2_X1 U435 ( .A(n384), .B(KEYINPUT17), .Z(n386) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(G183GAT), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n386), .B(n385), .ZN(n447) );
  XNOR2_X1 U438 ( .A(G211GAT), .B(KEYINPUT88), .ZN(n387) );
  XNOR2_X1 U439 ( .A(n387), .B(KEYINPUT87), .ZN(n388) );
  XOR2_X1 U440 ( .A(n388), .B(KEYINPUT21), .Z(n390) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G204GAT), .ZN(n389) );
  XNOR2_X1 U442 ( .A(n390), .B(n389), .ZN(n433) );
  XNOR2_X1 U443 ( .A(n447), .B(n433), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n517) );
  NAND2_X1 U445 ( .A1(n529), .A2(n517), .ZN(n394) );
  XOR2_X1 U446 ( .A(KEYINPUT54), .B(KEYINPUT123), .Z(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n419) );
  XOR2_X1 U448 ( .A(KEYINPUT0), .B(G134GAT), .Z(n396) );
  XNOR2_X1 U449 ( .A(KEYINPUT85), .B(G127GAT), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U451 ( .A(G113GAT), .B(n397), .ZN(n448) );
  XOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT94), .Z(n399) );
  XNOR2_X1 U453 ( .A(KEYINPUT93), .B(KEYINPUT95), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U455 ( .A(G148GAT), .B(G162GAT), .Z(n401) );
  XNOR2_X1 U456 ( .A(G141GAT), .B(G120GAT), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U458 ( .A(n403), .B(n402), .Z(n411) );
  XOR2_X1 U459 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n405) );
  XNOR2_X1 U460 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U462 ( .A(KEYINPUT2), .B(n406), .Z(n432) );
  XOR2_X1 U463 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n408) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(G57GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n432), .B(n409), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U468 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n413) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U471 ( .A(n415), .B(n414), .Z(n417) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(G85GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U474 ( .A(n448), .B(n418), .Z(n525) );
  NOR2_X2 U475 ( .A1(n419), .A2(n525), .ZN(n569) );
  XOR2_X1 U476 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n421) );
  XNOR2_X1 U477 ( .A(KEYINPUT91), .B(KEYINPUT23), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U479 ( .A(n422), .B(G106GAT), .Z(n425) );
  XNOR2_X1 U480 ( .A(n423), .B(G218GAT), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U482 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n459) );
  NAND2_X1 U488 ( .A1(n569), .A2(n459), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n436), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U490 ( .A(n437), .B(G176GAT), .Z(n439) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U493 ( .A(n440), .B(G99GAT), .Z(n445) );
  XOR2_X1 U494 ( .A(KEYINPUT66), .B(KEYINPUT20), .Z(n442) );
  INV_X1 U495 ( .A(G190GAT), .ZN(n452) );
  XNOR2_X1 U496 ( .A(G15GAT), .B(G190GAT), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U501 ( .A(n449), .B(n448), .Z(n532) );
  INV_X1 U502 ( .A(n532), .ZN(n519) );
  NAND2_X1 U503 ( .A1(n450), .A2(n519), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n451), .B(KEYINPUT124), .ZN(n566) );
  NOR2_X1 U505 ( .A1(n542), .A2(n566), .ZN(n454) );
  XOR2_X1 U506 ( .A(n459), .B(KEYINPUT28), .Z(n531) );
  XOR2_X1 U507 ( .A(n517), .B(KEYINPUT27), .Z(n527) );
  NOR2_X1 U508 ( .A1(n531), .A2(n527), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n532), .A2(n455), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n525), .A2(n456), .ZN(n466) );
  NAND2_X1 U511 ( .A1(n517), .A2(n519), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n459), .A2(n457), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT25), .B(n458), .Z(n464) );
  NOR2_X1 U514 ( .A1(n459), .A2(n519), .ZN(n461) );
  XNOR2_X1 U515 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n460) );
  XOR2_X1 U516 ( .A(n461), .B(n460), .Z(n548) );
  NOR2_X1 U517 ( .A1(n527), .A2(n548), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n462), .A2(n525), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n466), .A2(n465), .ZN(n483) );
  NAND2_X1 U521 ( .A1(n542), .A2(n467), .ZN(n468) );
  XNOR2_X1 U522 ( .A(KEYINPUT16), .B(n468), .ZN(n469) );
  NOR2_X1 U523 ( .A1(n483), .A2(n469), .ZN(n470) );
  XOR2_X1 U524 ( .A(KEYINPUT99), .B(n470), .Z(n499) );
  NOR2_X1 U525 ( .A1(n570), .A2(n471), .ZN(n486) );
  NAND2_X1 U526 ( .A1(n499), .A2(n486), .ZN(n472) );
  XOR2_X1 U527 ( .A(KEYINPUT100), .B(n472), .Z(n479) );
  NAND2_X1 U528 ( .A1(n479), .A2(n525), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n473), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n479), .A2(n517), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n475), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n477) );
  NAND2_X1 U534 ( .A1(n479), .A2(n519), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U536 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NAND2_X1 U537 ( .A1(n479), .A2(n531), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT102), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n489) );
  NOR2_X1 U541 ( .A1(n482), .A2(n483), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n484), .A2(n579), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n485), .B(KEYINPUT37), .ZN(n512) );
  NAND2_X1 U544 ( .A1(n512), .A2(n486), .ZN(n487) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(n487), .Z(n495) );
  NAND2_X1 U546 ( .A1(n495), .A2(n525), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U548 ( .A(G29GAT), .B(n490), .Z(G1328GAT) );
  NAND2_X1 U549 ( .A1(n495), .A2(n517), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n493) );
  NAND2_X1 U552 ( .A1(n495), .A2(n519), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U554 ( .A(G43GAT), .B(n494), .Z(G1330GAT) );
  NAND2_X1 U555 ( .A1(n495), .A2(n531), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  BUF_X1 U557 ( .A(n497), .Z(n562) );
  NOR2_X1 U558 ( .A1(n498), .A2(n562), .ZN(n513) );
  NAND2_X1 U559 ( .A1(n513), .A2(n499), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n500), .B(KEYINPUT105), .ZN(n508) );
  NAND2_X1 U561 ( .A1(n525), .A2(n508), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(KEYINPUT107), .ZN(n502) );
  XOR2_X1 U563 ( .A(n502), .B(KEYINPUT106), .Z(n504) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n508), .A2(n517), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n519), .A2(n508), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(KEYINPUT108), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U572 ( .A1(n508), .A2(n531), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  XOR2_X1 U575 ( .A(G85GAT), .B(KEYINPUT111), .Z(n516) );
  NAND2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U577 ( .A(KEYINPUT110), .B(n514), .Z(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n525), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n521), .A2(n519), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n523) );
  NAND2_X1 U585 ( .A1(n531), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  INV_X1 U588 ( .A(n525), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n528) );
  AND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT115), .B(n530), .Z(n549) );
  NOR2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n549), .A2(n533), .ZN(n541) );
  NOR2_X1 U594 ( .A1(n570), .A2(n541), .ZN(n534) );
  XOR2_X1 U595 ( .A(G113GAT), .B(n534), .Z(n535) );
  XNOR2_X1 U596 ( .A(KEYINPUT116), .B(n535), .ZN(G1340GAT) );
  NOR2_X1 U597 ( .A1(n562), .A2(n541), .ZN(n537) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NOR2_X1 U600 ( .A1(n579), .A2(n541), .ZN(n539) );
  XNOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  NOR2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n544) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(KEYINPUT118), .B(n545), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  INV_X1 U610 ( .A(n548), .ZN(n568) );
  NAND2_X1 U611 ( .A1(n568), .A2(n549), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT121), .B(n550), .Z(n558) );
  NOR2_X1 U613 ( .A1(n570), .A2(n558), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT122), .B(n551), .Z(n552) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  NOR2_X1 U616 ( .A1(n562), .A2(n558), .ZN(n554) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n579), .A2(n558), .ZN(n556) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  INV_X1 U622 ( .A(n557), .ZN(n559) );
  NOR2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NOR2_X1 U625 ( .A1(n570), .A2(n566), .ZN(n561) );
  XOR2_X1 U626 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  NOR2_X1 U627 ( .A1(n566), .A2(n562), .ZN(n564) );
  XNOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(n565), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n579), .A2(n566), .ZN(n567) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n582) );
  NOR2_X1 U634 ( .A1(n570), .A2(n582), .ZN(n572) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n582), .A2(n574), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n582), .ZN(n581) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n482), .A2(n582), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

