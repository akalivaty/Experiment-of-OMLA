//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n529, new_n530, new_n531, new_n532, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n589, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g037(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n459), .A2(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(KEYINPUT3), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n471), .A2(G137), .A3(new_n465), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n470), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G101), .A3(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n466), .A2(new_n477), .ZN(G160));
  AND2_X1   g053(.A1(new_n471), .A2(new_n473), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n471), .A2(new_n465), .A3(new_n473), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(G136), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT70), .ZN(G162));
  NAND2_X1  g062(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n473), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n465), .A3(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n465), .A2(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n471), .A2(new_n473), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n494), .B2(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n471), .A2(G126), .A3(G2105), .A4(new_n473), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n495), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT71), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(G543), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n514), .A2(new_n501), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n506), .A2(new_n507), .A3(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n510), .A2(new_n515), .A3(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  XNOR2_X1  g094(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n522), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n509), .A2(G51), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n516), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND2_X1  g103(.A1(new_n509), .A2(G52), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(new_n501), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(G90), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND2_X1  g109(.A1(new_n509), .A2(G43), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n501), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n516), .A2(G81), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  AOI22_X1  g120(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n501), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(G91), .B2(new_n516), .ZN(new_n548));
  NAND2_X1  g123(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n509), .A2(G53), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT73), .B(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n508), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(KEYINPUT74), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n550), .B2(new_n553), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n548), .B1(new_n555), .B2(new_n557), .ZN(G299));
  NAND4_X1  g133(.A1(new_n506), .A2(G49), .A3(G543), .A4(new_n507), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n506), .A2(G87), .A3(new_n507), .A4(new_n513), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(G288));
  INV_X1    g137(.A(G61), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n511), .B2(new_n512), .ZN(new_n564));
  AND2_X1   g139(.A1(G73), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n506), .A2(G48), .A3(G543), .A4(new_n507), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n506), .A2(G86), .A3(new_n507), .A4(new_n513), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G305));
  NAND2_X1  g147(.A1(new_n509), .A2(G47), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n516), .A2(G85), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n573), .B(new_n574), .C1(new_n501), .C2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n516), .A2(G92), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT10), .Z(new_n579));
  NAND2_X1  g154(.A1(new_n513), .A2(G66), .ZN(new_n580));
  NAND2_X1  g155(.A1(G79), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n501), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(G54), .B2(new_n509), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G284));
  OAI21_X1  g161(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G321));
  NAND2_X1  g162(.A1(G286), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(G299), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(G868), .ZN(G297));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(G868), .ZN(G280));
  XNOR2_X1  g166(.A(KEYINPUT76), .B(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(G860), .B2(new_n592), .ZN(G148));
  NAND2_X1  g168(.A1(new_n585), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g172(.A1(new_n475), .A2(new_n465), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n489), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT12), .Z(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT13), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(G2100), .ZN(new_n602));
  INV_X1    g177(.A(G2096), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n485), .A2(G135), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT77), .Z(new_n605));
  INV_X1    g180(.A(new_n480), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n465), .A2(G111), .ZN(new_n607));
  OAI21_X1  g182(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n606), .A2(G123), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n603), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n603), .B2(new_n612), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT78), .ZN(G156));
  XNOR2_X1  g190(.A(G2451), .B(G2454), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT16), .ZN(new_n617));
  XOR2_X1   g192(.A(G2443), .B(G2446), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G1341), .B(G1348), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT81), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT80), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n619), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT79), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2430), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n623), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(G14), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(G401));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  AND2_X1   g210(.A1(new_n635), .A2(KEYINPUT83), .ZN(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NOR3_X1   g213(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(KEYINPUT83), .B2(new_n635), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n635), .A2(KEYINPUT17), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(KEYINPUT17), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n641), .B(new_n642), .C1(new_n637), .C2(new_n638), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n638), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n635), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1971), .B(G1976), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n656), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT20), .Z(new_n660));
  AOI211_X1 g235(.A(new_n658), .B(new_n660), .C1(new_n653), .C2(new_n657), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G229));
  XOR2_X1   g242(.A(KEYINPUT85), .B(G16), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n669), .A2(G22), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(G166), .B2(new_n669), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT86), .Z(new_n672));
  OR2_X1    g247(.A1(new_n672), .A2(G1971), .ZN(new_n673));
  NOR2_X1   g248(.A1(G6), .A2(G16), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n571), .B2(G16), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT32), .B(G1981), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n672), .A2(G1971), .ZN(new_n684));
  NAND4_X1  g259(.A1(new_n673), .A2(new_n677), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n685), .A2(KEYINPUT34), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(KEYINPUT34), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n485), .A2(G131), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n465), .A2(G107), .ZN(new_n689));
  OAI21_X1  g264(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n690));
  INV_X1    g265(.A(G119), .ZN(new_n691));
  OAI221_X1 g266(.A(new_n688), .B1(new_n689), .B2(new_n690), .C1(new_n480), .C2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G25), .B(new_n692), .S(G29), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT35), .B(G1991), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT84), .ZN(new_n696));
  MUX2_X1   g271(.A(G24), .B(G290), .S(new_n669), .Z(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G1986), .Z(new_n698));
  NAND4_X1  g273(.A1(new_n686), .A2(new_n687), .A3(new_n696), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT36), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n669), .A2(G19), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n540), .B2(new_n669), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(G1341), .Z(new_n703));
  INV_X1    g278(.A(new_n598), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n704), .A2(G105), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n485), .A2(G141), .ZN(new_n710));
  INV_X1    g285(.A(G129), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n480), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G29), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G32), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n703), .B1(new_n717), .B2(KEYINPUT90), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n678), .A2(G4), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n585), .B2(new_n678), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1348), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n485), .A2(G139), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT87), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n723), .B(new_n726), .C1(new_n465), .C2(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G33), .B(new_n728), .S(G29), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT88), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n718), .B(new_n721), .C1(new_n731), .C2(G2072), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n668), .A2(G20), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT23), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n589), .B2(new_n678), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT97), .B(G1956), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n716), .B1(new_n713), .B2(new_n715), .ZN(new_n738));
  NOR2_X1   g313(.A1(G171), .A2(new_n678), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G5), .B2(new_n678), .ZN(new_n740));
  INV_X1    g315(.A(G1961), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n485), .A2(G140), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n465), .A2(G116), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n745));
  INV_X1    g320(.A(G128), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n743), .B1(new_n744), .B2(new_n745), .C1(new_n480), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n714), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2067), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(new_n714), .ZN(new_n756));
  INV_X1    g331(.A(G160), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n714), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2084), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n717), .A2(KEYINPUT90), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n742), .A2(new_n753), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n714), .A2(G27), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G164), .B2(new_n714), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT96), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT95), .B(G2078), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n737), .A2(new_n761), .A3(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n732), .B(new_n768), .C1(G2072), .C2(new_n731), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n678), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n678), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT92), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n740), .A2(new_n741), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(G1966), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n714), .B1(new_n777), .B2(G28), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(KEYINPUT91), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n777), .B2(G28), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(KEYINPUT91), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n775), .B(new_n782), .C1(new_n714), .C2(new_n611), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n773), .A2(new_n774), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(KEYINPUT93), .ZN(new_n785));
  NOR2_X1   g360(.A1(G29), .A2(G35), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G162), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT29), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n785), .B1(new_n788), .B2(G2090), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G2090), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(KEYINPUT93), .B2(new_n784), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n769), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n700), .A2(new_n792), .ZN(G150));
  INV_X1    g368(.A(G150), .ZN(G311));
  NAND2_X1  g369(.A1(new_n509), .A2(G55), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n516), .A2(G93), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n795), .B(new_n796), .C1(new_n501), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G860), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n585), .A2(G559), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n540), .B(new_n798), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT99), .ZN(new_n808));
  INV_X1    g383(.A(G860), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT100), .Z(new_n812));
  OAI21_X1  g387(.A(new_n801), .B1(new_n810), .B2(new_n812), .ZN(G145));
  INV_X1    g388(.A(KEYINPUT102), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n728), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n747), .B(G164), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n712), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n712), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n728), .A2(new_n814), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  XOR2_X1   g395(.A(new_n692), .B(KEYINPUT105), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n600), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n606), .A2(G130), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT103), .Z(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n825));
  INV_X1    g400(.A(G118), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n825), .A2(KEYINPUT104), .B1(new_n826), .B2(G2105), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(KEYINPUT104), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n485), .A2(G142), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n824), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n822), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n820), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n831), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n818), .B(new_n819), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n611), .B(new_n757), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G162), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  INV_X1    g415(.A(new_n838), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n832), .A2(new_n841), .A3(new_n835), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g419(.A(G868), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n571), .B(G290), .ZN(new_n846));
  XNOR2_X1  g421(.A(G303), .B(G288), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n848), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n850), .A2(KEYINPUT108), .B1(KEYINPUT42), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(KEYINPUT108), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n589), .A2(new_n585), .ZN(new_n854));
  NAND2_X1  g429(.A1(G299), .A2(new_n584), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(KEYINPUT41), .B2(new_n856), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n594), .B(new_n805), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n856), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n845), .B1(new_n853), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n853), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(KEYINPUT109), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT109), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n798), .B2(new_n845), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n865), .B1(new_n864), .B2(new_n867), .ZN(G295));
  AOI21_X1  g443(.A(new_n865), .B1(new_n864), .B2(new_n867), .ZN(G331));
  XNOR2_X1  g444(.A(G171), .B(G286), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(new_n805), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n805), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(KEYINPUT111), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT111), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n805), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n856), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n872), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n859), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n851), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n880));
  AOI21_X1  g455(.A(G37), .B1(new_n878), .B2(new_n851), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n856), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n857), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n875), .A3(new_n873), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(KEYINPUT41), .ZN(new_n886));
  OAI22_X1  g461(.A1(new_n885), .A2(new_n886), .B1(new_n856), .B2(new_n877), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n848), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g464(.A(KEYINPUT44), .B(new_n882), .C1(new_n889), .C2(new_n880), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n881), .A2(new_n880), .A3(new_n888), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n894));
  OAI21_X1  g469(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(G397));
  INV_X1    g470(.A(G1384), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n495), .B2(new_n499), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G40), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n473), .A2(new_n488), .A3(G125), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n462), .A2(new_n463), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n903), .B2(G2105), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n904), .A2(KEYINPUT112), .A3(new_n476), .A4(new_n474), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT112), .ZN(new_n906));
  OAI21_X1  g481(.A(G40), .B1(new_n464), .B2(new_n465), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(new_n477), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n899), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n712), .B(G1996), .Z(new_n911));
  XNOR2_X1  g486(.A(new_n747), .B(new_n752), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT113), .Z(new_n914));
  XOR2_X1   g489(.A(new_n692), .B(new_n694), .Z(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G290), .B(G1986), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n908), .A2(new_n905), .ZN(new_n919));
  OAI211_X1 g494(.A(KEYINPUT45), .B(new_n896), .C1(new_n495), .C2(new_n499), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n899), .A3(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(KEYINPUT56), .B(G2072), .Z(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n897), .A2(KEYINPUT50), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT50), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n925), .B(new_n896), .C1(new_n495), .C2(new_n499), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n919), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT122), .ZN(new_n928));
  INV_X1    g503(.A(G1956), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n927), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT57), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n554), .A2(new_n548), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(G299), .B2(KEYINPUT57), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n936), .B(new_n923), .C1(new_n930), .C2(new_n931), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1348), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n927), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n897), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n919), .A2(new_n943), .A3(new_n752), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n585), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n939), .B(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT59), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n919), .A2(new_n943), .ZN(new_n952));
  XOR2_X1   g527(.A(KEYINPUT58), .B(G1341), .Z(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n921), .A2(G1996), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n540), .B(new_n951), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT60), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n585), .A2(new_n942), .A3(new_n958), .A4(new_n944), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n921), .A2(G1996), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n539), .B1(new_n960), .B2(new_n954), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n962));
  OAI211_X1 g537(.A(new_n957), .B(new_n959), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n942), .A2(new_n584), .A3(new_n944), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n946), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n947), .B1(new_n949), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G2078), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n919), .A2(new_n899), .A3(new_n968), .A4(new_n920), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n927), .A2(new_n741), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(G2078), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n919), .A2(new_n899), .A3(new_n920), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(G301), .B(KEYINPUT54), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n969), .A2(new_n970), .B1(new_n927), .B2(new_n741), .ZN(new_n978));
  INV_X1    g553(.A(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(G40), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n465), .B1(new_n903), .B2(KEYINPUT124), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n980), .B(new_n477), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n899), .A3(new_n920), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1966), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n921), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2084), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n919), .A2(new_n924), .A3(new_n989), .A4(new_n926), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(G168), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G8), .ZN(new_n992));
  AOI21_X1  g567(.A(G168), .B1(new_n988), .B2(new_n990), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT51), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n995), .A3(G8), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n986), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1971), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n921), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G2090), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n919), .A2(new_n924), .A3(new_n1000), .A4(new_n926), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G303), .A2(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(G8), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT114), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n999), .B2(new_n1001), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n1005), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G288), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1012), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n952), .A2(new_n1014), .A3(G8), .A4(new_n1015), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1008), .B(new_n1013), .C1(new_n919), .C2(new_n943), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1008), .B1(new_n919), .B2(new_n943), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n569), .A2(G1981), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n1022));
  INV_X1    g597(.A(G1981), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n569), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1020), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT118), .B1(new_n1019), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1030), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(new_n1020), .A3(new_n1028), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1020), .A2(new_n1014), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT52), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .A4(new_n1016), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1007), .A2(new_n1011), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n1009), .B2(new_n1005), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1003), .B(KEYINPUT55), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n919), .A2(new_n924), .A3(new_n926), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1043), .A2(new_n1000), .B1(new_n921), .B2(new_n998), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1041), .B(new_n1042), .C1(new_n1044), .C2(new_n1008), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n997), .A2(new_n1039), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n967), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT125), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n994), .A2(new_n996), .A3(KEYINPUT62), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT62), .B1(new_n994), .B2(new_n996), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(G301), .B1(new_n978), .B2(new_n974), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1039), .A2(new_n1046), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1049), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1057));
  AND4_X1   g632(.A1(new_n1046), .A2(new_n1056), .A3(new_n1057), .A4(new_n1053), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(KEYINPUT125), .C1(new_n1051), .C2(new_n1050), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1048), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n680), .A2(new_n1012), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1024), .B1(new_n1031), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1020), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1034), .A2(new_n1036), .A3(new_n1016), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1063), .B(KEYINPUT116), .C1(new_n1056), .C2(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1042), .B1(new_n1044), .B2(new_n1008), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1043), .A2(new_n989), .B1(new_n921), .B2(new_n987), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G168), .A2(G8), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT119), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n988), .A2(new_n990), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(G8), .A4(G168), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1064), .A2(new_n1078), .ZN(new_n1079));
  AND4_X1   g654(.A1(new_n1070), .A2(new_n1056), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1056), .A2(new_n1057), .A3(new_n1046), .A4(new_n1077), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1078), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1082), .B2(KEYINPUT120), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1084), .A3(new_n1078), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1069), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1060), .B1(new_n1086), .B2(KEYINPUT121), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1088), .B(new_n1069), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n918), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n910), .A2(G1986), .A3(G290), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT48), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n916), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n692), .A2(new_n694), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT126), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n914), .A2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n747), .A2(G2067), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n910), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n912), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1099), .A2(new_n712), .ZN(new_n1100));
  OR3_X1    g675(.A1(new_n910), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT46), .B1(new_n910), .B2(G1996), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1100), .A2(new_n909), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT47), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1093), .A2(new_n1098), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1090), .A2(new_n1105), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g681(.A(G319), .ZN(new_n1108));
  OR2_X1    g682(.A1(G227), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g683(.A(G401), .B1(new_n1109), .B2(KEYINPUT127), .ZN(new_n1110));
  OAI21_X1  g684(.A(new_n1110), .B1(KEYINPUT127), .B2(new_n1109), .ZN(new_n1111));
  NOR2_X1   g685(.A1(G229), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g686(.A(new_n1112), .B(new_n843), .C1(new_n892), .C2(new_n891), .ZN(G225));
  INV_X1    g687(.A(G225), .ZN(G308));
endmodule


