//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n213), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G226), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G150), .ZN(new_n244));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  OAI22_X1  g0046(.A1(new_n244), .A2(new_n246), .B1(new_n201), .B2(new_n207), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT67), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT65), .A2(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT65), .A2(G20), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n247), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n214), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n207), .A3(G1), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n258), .B1(new_n206), .B2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n265), .B2(G50), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G223), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G222), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n271), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n273), .B1(new_n202), .B2(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g0083(.A(KEYINPUT66), .B(G41), .Z(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n206), .A2(G274), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n289), .B2(new_n285), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n288), .B1(G226), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G179), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n267), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n267), .A2(KEYINPUT9), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n260), .B2(new_n266), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n283), .B2(new_n292), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n294), .B2(G190), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n307), .A3(new_n304), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n297), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G68), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n245), .A2(G50), .B1(G20), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n254), .B2(new_n202), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n258), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT11), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n264), .A2(G68), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT70), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n261), .A2(G1), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(G20), .A3(new_n310), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT12), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n314), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(KEYINPUT14), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(KEYINPUT14), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n286), .A2(new_n287), .B1(new_n291), .B2(G238), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n278), .A2(G226), .A3(new_n271), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n278), .A2(G232), .A3(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n327), .A2(new_n328), .A3(new_n333), .A4(new_n329), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n282), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n325), .B(new_n326), .C1(new_n332), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(new_n282), .A3(new_n334), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n325), .B1(new_n338), .B2(new_n326), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n323), .B(new_n324), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n326), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT13), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G179), .A3(new_n336), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n336), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n324), .B1(new_n345), .B2(new_n323), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n320), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n302), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n342), .A2(new_n349), .A3(new_n336), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n320), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n213), .A2(G77), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  OAI221_X1 g0155(.A(new_n354), .B1(new_n246), .B2(new_n248), .C1(new_n254), .C2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n356), .A2(new_n258), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n262), .A2(new_n202), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n265), .B2(new_n202), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n272), .A2(G238), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n270), .A2(G107), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n363), .C1(new_n231), .C2(new_n280), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n282), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n288), .B1(G244), .B2(new_n291), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT68), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT68), .B1(new_n365), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n349), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n365), .A2(new_n366), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT68), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT68), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n302), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n361), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(G179), .B1(new_n367), .B2(new_n368), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(G169), .A3(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n360), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n309), .A2(new_n347), .A3(new_n353), .A4(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n253), .A2(new_n270), .A3(KEYINPUT7), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n276), .A2(new_n207), .A3(new_n277), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G68), .ZN(new_n386));
  INV_X1    g0186(.A(G58), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n310), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G58), .A2(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n245), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n259), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT72), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n383), .B1(new_n278), .B2(new_n213), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n392), .B1(new_n400), .B2(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n253), .B2(new_n270), .ZN(new_n403));
  NOR4_X1   g0203(.A1(new_n268), .A2(new_n269), .A3(new_n383), .A4(G20), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n405), .A2(new_n397), .A3(KEYINPUT16), .A4(new_n393), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n396), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n250), .A2(new_n262), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n265), .B2(new_n250), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n278), .A2(G223), .A3(new_n271), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  OAI211_X1 g0213(.A(G226), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n282), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT73), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n286), .A2(new_n287), .B1(new_n291), .B2(G232), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(KEYINPUT73), .A3(new_n282), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n418), .A2(new_n349), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n416), .A2(new_n419), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n302), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n408), .A2(new_n411), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n393), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT72), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n406), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n410), .B1(new_n430), .B2(new_n396), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT17), .A3(new_n424), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n408), .A2(new_n411), .ZN(new_n435));
  INV_X1    g0235(.A(new_n420), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT73), .B1(new_n415), .B2(new_n282), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G179), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n419), .A2(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n438), .A2(new_n440), .B1(new_n321), .B2(new_n422), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n434), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n418), .A3(new_n420), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n422), .A2(new_n321), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n431), .A2(KEYINPUT18), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT74), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT18), .B1(new_n431), .B2(new_n445), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT74), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n392), .B1(new_n385), .B2(G68), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n258), .B1(new_n450), .B2(KEYINPUT16), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n406), .B2(new_n429), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n441), .B(new_n434), .C1(new_n452), .C2(new_n410), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n433), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n380), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n272), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n278), .A2(G244), .A3(new_n271), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT77), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT4), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n459), .B2(new_n460), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n282), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT78), .ZN(new_n466));
  INV_X1    g0266(.A(new_n464), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n462), .A3(new_n458), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT78), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n282), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n206), .B(G45), .C1(new_n471), .C2(G41), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT66), .B(G41), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n471), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n282), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(G257), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(G274), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n466), .A2(new_n470), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G200), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n262), .B1(new_n206), .B2(G33), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(KEYINPUT76), .A3(new_n259), .ZN(new_n484));
  INV_X1    g0284(.A(new_n262), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n206), .A2(G33), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n259), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT76), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G97), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(G97), .B2(new_n262), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n465), .A2(new_n480), .A3(G190), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(new_n213), .B1(G77), .B2(new_n245), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n385), .A2(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n259), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT75), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n504), .A2(KEYINPUT75), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n492), .B(new_n493), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(G169), .B1(new_n465), .B2(new_n480), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n504), .B(KEYINPUT75), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n492), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n466), .A2(new_n439), .A3(new_n470), .A4(new_n480), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n482), .A2(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n278), .A2(G264), .A3(G1698), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n278), .A2(G257), .A3(new_n271), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n270), .A2(G303), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n282), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n474), .A2(new_n282), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G270), .ZN(new_n521));
  AND4_X1   g0321(.A1(G179), .A2(new_n519), .A3(new_n521), .A4(new_n478), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n519), .A2(new_n521), .A3(new_n478), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(KEYINPUT21), .A3(G169), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT81), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n253), .B(new_n528), .C1(G33), .C2(new_n495), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G20), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n259), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT20), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n527), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n529), .A2(new_n533), .A3(KEYINPUT81), .A4(KEYINPUT20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n535), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT80), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n487), .B2(new_n530), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n483), .A2(KEYINPUT80), .A3(G116), .A4(new_n259), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n541), .A2(new_n542), .B1(new_n317), .B2(new_n532), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n526), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n539), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n524), .A2(G169), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n519), .A2(new_n521), .A3(new_n478), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n349), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n524), .A2(new_n302), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n544), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n278), .A2(G250), .A3(new_n271), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n278), .A2(G257), .A3(G1698), .ZN(new_n557));
  XNOR2_X1  g0357(.A(KEYINPUT84), .B(G294), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n556), .B(new_n557), .C1(new_n275), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n282), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n520), .A2(G264), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n478), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n302), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(G190), .B2(new_n563), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n278), .A2(new_n253), .A3(G87), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT22), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT23), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n213), .A2(new_n570), .A3(new_n496), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G116), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n570), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n207), .B1(KEYINPUT23), .B2(G107), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n571), .A2(KEYINPUT83), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT83), .B1(new_n571), .B2(new_n574), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n568), .B(new_n569), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  XOR2_X1   g0377(.A(KEYINPUT82), .B(KEYINPUT24), .Z(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n566), .B(KEYINPUT22), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n578), .C1(new_n576), .C2(new_n575), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n582), .A3(new_n258), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n490), .A2(new_n496), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n262), .A2(new_n496), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n585), .B(KEYINPUT25), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n565), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n563), .A2(new_n439), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n563), .A2(G169), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n583), .A2(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n254), .B2(new_n495), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n278), .A2(new_n253), .A3(G68), .ZN(new_n594));
  INV_X1    g0394(.A(G87), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n495), .A3(new_n496), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n329), .A2(new_n592), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n213), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n258), .ZN(new_n600));
  INV_X1    g0400(.A(new_n355), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n484), .A2(new_n489), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n355), .A2(new_n262), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n287), .A2(G45), .ZN(new_n605));
  OAI21_X1  g0405(.A(G250), .B1(new_n285), .B2(G1), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n282), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n278), .A2(G238), .A3(new_n271), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n278), .A2(G244), .A3(G1698), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n572), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n607), .B1(new_n610), .B2(new_n282), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n321), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n439), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n604), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n611), .A2(KEYINPUT79), .A3(G190), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT79), .B1(new_n611), .B2(G190), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n599), .A2(new_n258), .B1(new_n262), .B2(new_n355), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n484), .A2(new_n489), .A3(G87), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n302), .C2(new_n611), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n615), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n588), .A2(new_n591), .A3(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n457), .A2(new_n514), .A3(new_n555), .A4(new_n623), .ZN(G372));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n448), .A2(new_n625), .A3(new_n453), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n448), .B2(new_n453), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n323), .B1(new_n337), .B2(new_n339), .ZN(new_n629));
  INV_X1    g0429(.A(new_n324), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n340), .A3(new_n343), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n378), .B1(new_n632), .B2(new_n320), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n427), .A2(new_n432), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n353), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n628), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n306), .A2(new_n308), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n297), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n380), .A2(new_n456), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n619), .A2(new_n602), .B1(new_n439), .B2(new_n611), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n641));
  OR3_X1    g0441(.A1(new_n611), .A2(KEYINPUT85), .A3(G169), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n612), .A2(G200), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n611), .A2(G190), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n644), .A2(new_n619), .A3(new_n620), .A4(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n565), .A2(new_n583), .A3(new_n587), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n647), .B(new_n648), .C1(new_n550), .C2(new_n591), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n509), .A2(new_n482), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n511), .A2(new_n492), .ZN(new_n651));
  INV_X1    g0451(.A(new_n510), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n513), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n643), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n651), .A2(new_n513), .A3(new_n652), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n647), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n653), .B2(new_n622), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n638), .B1(new_n639), .B2(new_n661), .ZN(G369));
  INV_X1    g0462(.A(new_n548), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT21), .B1(new_n663), .B2(new_n544), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n544), .B2(new_n526), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n253), .A2(new_n317), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G343), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n665), .A2(new_n544), .A3(new_n672), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n550), .A2(new_n554), .B1(new_n547), .B2(new_n671), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n583), .A2(new_n587), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n672), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n648), .ZN(new_n678));
  INV_X1    g0478(.A(new_n591), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n679), .B2(new_n672), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT87), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n675), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n665), .A2(new_n672), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n686), .A2(new_n680), .B1(new_n591), .B2(new_n671), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(KEYINPUT89), .ZN(new_n689));
  INV_X1    g0489(.A(new_n210), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n473), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n210), .A2(KEYINPUT89), .A3(new_n284), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n595), .A2(new_n495), .A3(new_n496), .A4(new_n530), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT88), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n206), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n216), .B2(new_n693), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  AND4_X1   g0500(.A1(new_n439), .A2(new_n563), .A3(new_n524), .A4(new_n612), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n481), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n479), .B1(new_n468), .B2(new_n282), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n611), .A2(new_n562), .A3(new_n561), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n522), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g0505(.A(KEYINPUT90), .B(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n481), .A2(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT91), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n703), .A2(new_n704), .A3(new_n522), .A4(KEYINPUT30), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n671), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n702), .A2(new_n707), .A3(new_n713), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n672), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n714), .A2(new_n716), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n514), .A2(new_n623), .A3(new_n555), .A4(new_n671), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n700), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n657), .B1(new_n653), .B2(new_n622), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT92), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT92), .B(new_n657), .C1(new_n653), .C2(new_n622), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n647), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n643), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n648), .A2(new_n643), .A3(new_n646), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n665), .B2(new_n679), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(new_n730), .B2(new_n514), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n672), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n671), .B1(new_n655), .B2(new_n660), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n721), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n699), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(new_n693), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n213), .A2(new_n261), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n206), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n673), .A2(new_n674), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n213), .A2(G179), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT94), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n349), .A2(new_n302), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n349), .A2(G179), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n253), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(G326), .B1(new_n558), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT97), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(KEYINPUT97), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n753), .A2(new_n349), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n253), .A2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n278), .B1(new_n770), .B2(G329), .ZN(new_n771));
  INV_X1    g0571(.A(G283), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n302), .A2(G179), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n767), .ZN(new_n775));
  INV_X1    g0575(.A(G303), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n207), .A2(new_n349), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n771), .B1(new_n772), .B2(new_n775), .C1(new_n776), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n349), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n753), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n779), .B1(G322), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n761), .A2(new_n762), .A3(new_n766), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n753), .A2(new_n349), .A3(new_n302), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT95), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n789), .A2(new_n202), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n770), .A2(G159), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  INV_X1    g0594(.A(new_n775), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G107), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n270), .B1(new_n758), .B2(G97), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(new_n595), .C2(new_n778), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G58), .A2(new_n782), .B1(new_n755), .B2(G50), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(new_n310), .C2(new_n763), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n784), .A2(new_n791), .B1(new_n792), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n214), .B1(G20), .B2(new_n321), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n748), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(G355), .B(KEYINPUT93), .Z(new_n805));
  NOR2_X1   g0605(.A1(new_n690), .A2(new_n270), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n690), .A2(new_n278), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n217), .A2(G45), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n239), .B2(G45), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n807), .B1(G116), .B2(new_n210), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n744), .B1(new_n750), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n745), .B(G330), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n744), .B2(new_n815), .ZN(G396));
  NOR2_X1   g0616(.A1(new_n803), .A2(new_n746), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n744), .B1(new_n202), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n378), .A2(new_n671), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n360), .A2(new_n671), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n369), .A2(new_n374), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n821), .B2(new_n360), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n819), .B1(new_n822), .B2(new_n378), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n270), .B1(new_n495), .B2(new_n757), .C1(new_n778), .C2(new_n496), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n775), .A2(new_n595), .B1(new_n769), .B2(new_n790), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(G303), .C2(new_n755), .ZN(new_n827));
  INV_X1    g0627(.A(G294), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n772), .B2(new_n763), .C1(new_n828), .C2(new_n781), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G116), .B2(new_n788), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G143), .A2(new_n782), .B1(new_n755), .B2(G137), .ZN(new_n831));
  INV_X1    g0631(.A(G159), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n244), .B2(new_n763), .C1(new_n789), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT34), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n775), .A2(new_n310), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n278), .B1(new_n387), .B2(new_n757), .C1(new_n769), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n778), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n835), .B(new_n837), .C1(G50), .C2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n830), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n803), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n818), .B1(new_n747), .B2(new_n824), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n734), .B(new_n824), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT98), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n721), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n744), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n843), .B2(new_n721), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT99), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n843), .A2(new_n721), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n848), .A2(KEYINPUT99), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n842), .B1(new_n851), .B2(new_n852), .ZN(G384));
  OAI21_X1  g0653(.A(new_n441), .B1(new_n452), .B2(new_n410), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n670), .B1(new_n452), .B2(new_n410), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n425), .A4(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n425), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT101), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n405), .B2(new_n393), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n860), .B2(new_n259), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT101), .B(new_n258), .C1(new_n401), .C2(KEYINPUT16), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n430), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n445), .B1(new_n863), .B2(new_n411), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n669), .B1(new_n863), .B2(new_n411), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n858), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n857), .B1(new_n866), .B2(new_n856), .ZN(new_n867));
  INV_X1    g0667(.A(new_n865), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT38), .B(new_n867), .C1(new_n455), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT103), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n626), .A2(new_n627), .A3(new_n433), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n855), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT86), .B1(new_n442), .B2(new_n446), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n448), .A2(new_n625), .A3(new_n453), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n634), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n855), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(KEYINPUT103), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n854), .A2(new_n855), .A3(new_n425), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT102), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT102), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n882), .A3(KEYINPUT37), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n857), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n873), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n870), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n671), .B1(new_n710), .B2(new_n713), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT104), .B1(new_n888), .B2(KEYINPUT31), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(KEYINPUT31), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n718), .A2(new_n891), .A3(new_n715), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n720), .A2(new_n889), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n320), .B1(new_n348), .B2(new_n350), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n320), .B(new_n672), .C1(new_n632), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n320), .A2(new_n672), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n347), .A2(new_n353), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n823), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n893), .A2(new_n898), .A3(KEYINPUT40), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT105), .B1(new_n887), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n878), .A2(new_n884), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT103), .B1(new_n876), .B2(new_n877), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n886), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n869), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT105), .ZN(new_n905));
  INV_X1    g0705(.A(new_n899), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n867), .B1(new_n455), .B2(new_n868), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n886), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n869), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n893), .A3(new_n898), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n900), .A2(new_n907), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n457), .A2(new_n893), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n915), .A2(new_n916), .A3(new_n700), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n669), .B1(new_n626), .B2(new_n627), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n819), .B1(new_n734), .B2(new_n823), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n895), .A2(new_n897), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n911), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n910), .B2(new_n869), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n887), .B2(new_n924), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n632), .A2(new_n320), .A3(new_n671), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n923), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n733), .A2(new_n457), .A3(new_n736), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n638), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n917), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n917), .A2(new_n933), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(new_n206), .C2(new_n740), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n501), .A2(KEYINPUT35), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n253), .A2(new_n214), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n501), .A2(KEYINPUT35), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n937), .A2(G116), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT36), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(KEYINPUT36), .ZN(new_n943));
  OAI21_X1  g0743(.A(G77), .B1(new_n387), .B2(new_n310), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n944), .A2(new_n216), .B1(G50), .B2(new_n310), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(G1), .A3(new_n261), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT100), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n936), .A2(new_n948), .ZN(G367));
  AND2_X1   g0749(.A1(new_n808), .A2(new_n235), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n804), .B1(new_n210), .B2(new_n355), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n775), .A2(new_n202), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n278), .B1(new_n310), .B2(new_n757), .C1(new_n778), .C2(new_n387), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(G137), .C2(new_n770), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n244), .B2(new_n781), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G143), .B2(new_n755), .ZN(new_n956));
  INV_X1    g0756(.A(G50), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n956), .B1(new_n957), .B2(new_n789), .C1(new_n832), .C2(new_n763), .ZN(new_n958));
  INV_X1    g0758(.A(new_n755), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n959), .A2(new_n790), .B1(new_n776), .B2(new_n781), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n775), .A2(new_n495), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n778), .A2(new_n530), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT46), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n278), .B1(new_n758), .B2(G107), .ZN(new_n964));
  INV_X1    g0764(.A(G317), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n964), .B1(new_n965), .B2(new_n769), .ZN(new_n966));
  NOR4_X1   g0766(.A1(new_n960), .A2(new_n961), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n559), .B2(new_n763), .C1(new_n772), .C2(new_n789), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n958), .A2(KEYINPUT47), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n803), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT47), .B1(new_n958), .B2(new_n968), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n743), .B1(new_n950), .B2(new_n951), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT111), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n671), .B1(new_n619), .B2(new_n620), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n643), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n647), .B2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n748), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  NOR4_X1   g0780(.A1(new_n678), .A2(new_n665), .A3(new_n591), .A4(new_n672), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n651), .A2(new_n672), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n650), .A2(new_n653), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n656), .A2(new_n672), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n650), .A2(new_n591), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n672), .B1(new_n988), .B2(new_n653), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n986), .B2(KEYINPUT42), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n978), .B(KEYINPUT43), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n991), .A2(KEYINPUT107), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT107), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT108), .ZN(new_n996));
  INV_X1    g0796(.A(new_n685), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n985), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT43), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n978), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n987), .A2(new_n990), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT106), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT106), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n987), .A2(new_n990), .A3(new_n1004), .A4(new_n1001), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n995), .A2(new_n996), .A3(new_n999), .A4(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n999), .C1(new_n994), .C2(new_n993), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n993), .A2(new_n994), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1006), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n998), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1007), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n687), .A2(new_n985), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n1017));
  OR3_X1    g0817(.A1(new_n687), .A2(new_n985), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n687), .B2(new_n985), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(KEYINPUT110), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT110), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n1017), .C1(new_n687), .C2(new_n985), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n997), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1016), .A2(new_n1020), .A3(new_n685), .A4(new_n1022), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n681), .B(new_n686), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(new_n675), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n737), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n737), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n693), .B(KEYINPUT41), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n742), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n980), .B1(new_n1013), .B2(new_n1032), .ZN(G387));
  OAI21_X1  g0833(.A(new_n270), .B1(new_n775), .B2(new_n530), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT113), .B(G322), .Z(new_n1035));
  AOI22_X1  g0835(.A1(G317), .A2(new_n782), .B1(new_n755), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n790), .B2(new_n763), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G303), .B2(new_n788), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT48), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(KEYINPUT48), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n838), .A2(new_n558), .B1(G283), .B2(new_n758), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1034), .B(new_n1044), .C1(G326), .C2(new_n770), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n778), .A2(new_n202), .B1(new_n769), .B2(new_n244), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n757), .A2(new_n355), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n1046), .A2(new_n961), .A3(new_n270), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n764), .A2(new_n250), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n755), .A2(G159), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n782), .A2(G50), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G68), .B2(new_n788), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n803), .B1(new_n1045), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n806), .A2(new_n695), .B1(new_n496), .B2(new_n690), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT112), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n232), .A2(G45), .ZN(new_n1057));
  AOI211_X1 g0857(.A(G45), .B(new_n695), .C1(G68), .C2(G77), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n248), .A2(G50), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n809), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1056), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n804), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n743), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n681), .B2(new_n748), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1054), .A2(new_n1065), .B1(new_n742), .B2(new_n1027), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n737), .A2(new_n1027), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n739), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n737), .A2(new_n1027), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(G393));
  NAND2_X1  g0870(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n1067), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n739), .A3(new_n1028), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n804), .B1(new_n495), .B2(new_n210), .C1(new_n809), .C2(new_n242), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n743), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n985), .A2(new_n749), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n959), .A2(new_n965), .B1(new_n790), .B2(new_n781), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n778), .A2(new_n772), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n278), .B1(new_n758), .B2(G116), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n796), .A2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(new_n770), .C2(new_n1035), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1078), .B(new_n1082), .C1(new_n776), .C2(new_n763), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n789), .A2(new_n828), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G159), .A2(new_n782), .B1(new_n755), .B2(G150), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n838), .A2(G68), .B1(new_n770), .B2(G143), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n270), .B1(new_n758), .B2(G77), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n595), .C2(new_n775), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G50), .B2(new_n764), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n789), .B2(new_n248), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1083), .A2(new_n1084), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1075), .B(new_n1076), .C1(new_n803), .C2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n742), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1073), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT115), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1073), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n921), .A2(new_n928), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n903), .A2(new_n924), .A3(new_n869), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n925), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n920), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n376), .A2(new_n377), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n361), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n375), .B2(new_n820), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n732), .A2(new_n1108), .B1(new_n378), .B2(new_n671), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n904), .B(new_n928), .C1(new_n1105), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n721), .A2(new_n898), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1104), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n887), .A2(new_n929), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n732), .A2(new_n1108), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n819), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n920), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n926), .A2(new_n1101), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n893), .A2(new_n898), .A3(G330), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1112), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n893), .A2(G330), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT116), .B1(new_n639), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT116), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n457), .A2(new_n1123), .A3(G330), .A4(new_n893), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n931), .A2(new_n1122), .A3(new_n1124), .A4(new_n638), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n920), .B1(new_n721), .B2(new_n824), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n919), .B1(new_n1126), .B2(new_n1118), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1105), .B1(new_n1121), .B2(new_n823), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1109), .A2(new_n1128), .A3(new_n1111), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1125), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1120), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1112), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n739), .A3(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1120), .A2(new_n741), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n817), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n743), .B1(new_n250), .B2(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n775), .A2(new_n310), .B1(new_n769), .B2(new_n828), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n270), .B1(new_n202), .B2(new_n757), .C1(new_n778), .C2(new_n595), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(new_n782), .C2(G116), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n496), .B2(new_n763), .C1(new_n772), .C2(new_n959), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n789), .A2(new_n495), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n838), .A2(G150), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT53), .Z(new_n1144));
  AOI22_X1  g0944(.A1(G132), .A2(new_n782), .B1(new_n755), .B2(G128), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n764), .A2(G137), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n278), .B1(new_n832), .B2(new_n757), .C1(new_n769), .C2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G50), .B2(new_n795), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n789), .A2(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1141), .A2(new_n1142), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1137), .B1(new_n1153), .B2(new_n803), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n927), .B2(new_n747), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT117), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1134), .A2(new_n1135), .A3(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(new_n309), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n267), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n670), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n309), .B1(new_n267), .B2(new_n669), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n746), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n743), .B1(G50), .B2(new_n1136), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n957), .B1(G33), .B2(G41), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n284), .B2(new_n270), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n795), .A2(G58), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n310), .B2(new_n757), .C1(new_n772), .C2(new_n769), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G107), .B2(new_n782), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n270), .B(new_n284), .C1(new_n778), .C2(new_n202), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT118), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n755), .A2(G116), .B1(KEYINPUT118), .B2(new_n1174), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n764), .A2(G97), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n601), .B2(new_n788), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1170), .B1(new_n1179), .B2(KEYINPUT58), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n782), .A2(G128), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1151), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n838), .A2(new_n1182), .B1(G150), .B2(new_n758), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n1147), .B2(new_n959), .C1(new_n836), .C2(new_n763), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G137), .B2(new_n788), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G33), .B(G41), .C1(new_n795), .C2(G159), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT119), .B(G124), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1188), .B(new_n1189), .C1(new_n769), .C2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1180), .B1(KEYINPUT58), .B2(new_n1179), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1168), .B1(new_n1193), .B2(new_n803), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1167), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n918), .B1(new_n922), .B2(new_n921), .C1(new_n926), .C2(new_n928), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n893), .A2(new_n898), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n869), .B2(new_n910), .ZN(new_n1199));
  OAI21_X1  g0999(.A(G330), .B1(new_n1199), .B2(KEYINPUT40), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1166), .B(new_n1200), .C1(new_n907), .C2(new_n900), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1166), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n900), .A2(new_n907), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n700), .B1(new_n912), .B2(new_n908), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1197), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(new_n1207));
  AOI211_X1 g1007(.A(KEYINPUT105), .B(new_n899), .C1(new_n903), .C2(new_n869), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1204), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1166), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1203), .A2(new_n1204), .A3(new_n1202), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n930), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1206), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1196), .B1(new_n1213), .B2(new_n742), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1125), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1133), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT57), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT120), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1210), .A2(new_n1218), .A3(new_n930), .A4(new_n1211), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1206), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1212), .A2(KEYINPUT120), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1217), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1206), .A2(new_n1212), .B1(new_n1215), .B2(new_n1133), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n739), .B1(new_n1223), .B2(KEYINPUT57), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1214), .B1(new_n1222), .B2(new_n1224), .ZN(G375));
  AND2_X1   g1025(.A1(new_n1129), .A2(new_n1127), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1125), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT121), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT121), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1229), .A3(new_n1125), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1228), .A2(new_n1131), .A3(new_n1031), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1226), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1105), .A2(new_n746), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n743), .B1(G68), .B2(new_n1136), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n778), .A2(new_n495), .B1(new_n769), .B2(new_n776), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n952), .A2(new_n278), .A3(new_n1047), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(G283), .C2(new_n782), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(new_n530), .B2(new_n763), .C1(new_n828), .C2(new_n959), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n789), .A2(new_n496), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n789), .A2(new_n244), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n778), .A2(new_n832), .B1(new_n957), .B2(new_n757), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT122), .B1(new_n1171), .B2(new_n278), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G128), .C2(new_n770), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1171), .A2(KEYINPUT122), .A3(new_n278), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G137), .A2(new_n782), .B1(new_n755), .B2(G132), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n764), .A2(new_n1182), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1238), .A2(new_n1239), .B1(new_n1240), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1234), .B1(new_n1248), .B2(new_n803), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1232), .A2(new_n742), .B1(new_n1233), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1231), .A2(new_n1250), .ZN(G381));
  NOR2_X1   g1051(.A1(G375), .A2(G378), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1099), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1098), .B1(new_n1073), .B2(new_n1095), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(G387), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(G381), .A2(G384), .A3(G396), .A4(G393), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1255), .A3(new_n1256), .ZN(G407));
  INV_X1    g1057(.A(new_n1252), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G407), .B(G213), .C1(G343), .C2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT123), .ZN(G409));
  OR2_X1    g1060(.A1(new_n1013), .A2(new_n1032), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1261), .A2(new_n980), .A3(new_n1099), .A4(new_n1097), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G390), .A2(G387), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G393), .B(G396), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1265), .A2(new_n1266), .A3(KEYINPUT126), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1264), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1261), .A2(new_n980), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n1255), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1268), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT127), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT126), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1271), .A2(new_n1268), .A3(new_n1272), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G213), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(G343), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(G2897), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1228), .B(new_n1230), .C1(new_n1284), .C2(new_n1130), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1227), .A2(new_n1284), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1286), .A2(new_n693), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(G384), .A3(new_n1250), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1288), .B2(new_n1250), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1283), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1250), .ZN(new_n1293));
  INV_X1    g1093(.A(G384), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1289), .A3(new_n1282), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1196), .B1(new_n1223), .B2(new_n1031), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1212), .A2(KEYINPUT120), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1206), .A2(new_n1219), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n742), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G378), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1213), .A2(new_n742), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1195), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1201), .A2(new_n1205), .A3(new_n1197), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n930), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1216), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT57), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n693), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(KEYINPUT57), .B(new_n1216), .C1(new_n1299), .C2(new_n1300), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1304), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1302), .B1(new_n1311), .B2(G378), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1297), .B1(new_n1312), .B2(new_n1281), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G378), .B(new_n1214), .C1(new_n1222), .C2(new_n1224), .ZN(new_n1315));
  INV_X1    g1115(.A(G378), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n741), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1216), .B(new_n1031), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1195), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1316), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1315), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1281), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1295), .A2(new_n1289), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .A4(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1313), .A2(new_n1314), .A3(new_n1326), .ZN(new_n1327));
  AOI211_X1 g1127(.A(new_n1281), .B(new_n1324), .C1(new_n1315), .C2(new_n1320), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1328), .A2(new_n1322), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1279), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1281), .B1(new_n1315), .B2(new_n1320), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1314), .B(new_n1331), .C1(new_n1332), .C2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT124), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1328), .B2(KEYINPUT63), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1332), .A2(new_n1325), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT63), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1338), .A2(KEYINPUT124), .A3(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1335), .A2(new_n1337), .A3(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1321), .A2(KEYINPUT63), .A3(new_n1323), .A4(new_n1325), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(KEYINPUT125), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1330), .B1(new_n1341), .B2(new_n1343), .ZN(G405));
  OAI21_X1  g1144(.A(new_n1325), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1275), .A2(new_n1276), .A3(new_n1324), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1311), .B(new_n1316), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1347), .B(new_n1348), .ZN(G402));
endmodule


