//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G128), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n195), .B1(G143), .B2(new_n189), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n195), .A3(G128), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT0), .B(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT0), .A4(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT64), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n198), .A2(new_n207), .A3(KEYINPUT0), .A4(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n202), .B1(new_n201), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G224), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G953), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n210), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G101), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT67), .A2(G119), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT67), .A2(G119), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(G116), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G119), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n226), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n233), .B1(new_n226), .B2(new_n228), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n223), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n221), .A2(G101), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n216), .A2(new_n219), .A3(new_n238), .A4(new_n220), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT82), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n226), .A2(KEYINPUT5), .A3(new_n228), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n242), .B(G113), .C1(KEYINPUT5), .C2(new_n226), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n226), .A2(new_n228), .A3(new_n233), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n215), .A2(G107), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n218), .A2(G104), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n243), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n226), .A2(new_n228), .ZN(new_n250));
  INV_X1    g064(.A(new_n233), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n244), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT82), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .A4(new_n223), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n241), .A2(new_n249), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G122), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n256), .A2(new_n249), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n262), .A2(KEYINPUT83), .A3(new_n259), .A4(new_n241), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n241), .A2(new_n259), .A3(new_n249), .A4(new_n256), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n258), .B1(new_n257), .B2(new_n260), .ZN(new_n268));
  AOI211_X1 g082(.A(new_n214), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT7), .B(new_n213), .C1(new_n210), .C2(KEYINPUT84), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n209), .A2(new_n201), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n213), .A2(KEYINPUT7), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n271), .A2(new_n202), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n243), .A2(new_n244), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n239), .A2(new_n247), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n249), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n259), .B(KEYINPUT8), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n270), .A2(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n267), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n188), .B1(new_n269), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n267), .A2(new_n268), .ZN(new_n285));
  INV_X1    g099(.A(new_n261), .ZN(new_n286));
  INV_X1    g100(.A(new_n214), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n267), .B2(new_n280), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n187), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(G475), .A2(G902), .ZN(new_n292));
  XNOR2_X1  g106(.A(G113), .B(G122), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(new_n215), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT85), .ZN(new_n295));
  INV_X1    g109(.A(G237), .ZN(new_n296));
  INV_X1    g110(.A(G953), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(G214), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(new_n191), .ZN(new_n299));
  NOR2_X1   g113(.A1(G237), .A2(G953), .ZN(new_n300));
  AOI21_X1  g114(.A(G143), .B1(new_n300), .B2(G214), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n299), .A2(new_n301), .A3(G131), .ZN(new_n302));
  INV_X1    g116(.A(G131), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n191), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(G143), .A3(G214), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n295), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G125), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n201), .A2(G140), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n201), .A2(KEYINPUT71), .A3(G140), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT16), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G146), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT19), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n312), .B2(new_n313), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(KEYINPUT19), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n189), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G131), .B1(new_n299), .B2(new_n301), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n304), .A2(new_n303), .A3(new_n305), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(KEYINPUT85), .A3(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n307), .A2(new_n318), .A3(new_n323), .A4(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n312), .A2(G146), .A3(new_n313), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n189), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n304), .A2(new_n305), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(KEYINPUT18), .B(G131), .C1(new_n299), .C2(new_n301), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n294), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT86), .ZN(new_n336));
  INV_X1    g150(.A(new_n334), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT17), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n324), .A2(new_n338), .A3(new_n325), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n306), .A2(KEYINPUT17), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n314), .A2(new_n189), .A3(new_n316), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n189), .B1(new_n314), .B2(new_n316), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n337), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n294), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n335), .A2(KEYINPUT86), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n292), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT20), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n335), .A2(KEYINPUT86), .B1(new_n345), .B2(new_n294), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n327), .A2(new_n334), .ZN(new_n352));
  INV_X1    g166(.A(new_n294), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT86), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT20), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n292), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n345), .B(new_n294), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n282), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n350), .A2(new_n359), .B1(G475), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n227), .A2(G122), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n227), .A2(G122), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(KEYINPUT14), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(KEYINPUT14), .ZN(new_n367));
  INV_X1    g181(.A(new_n364), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT89), .B1(new_n364), .B2(KEYINPUT14), .ZN(new_n370));
  OAI211_X1 g184(.A(G107), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n368), .A2(new_n365), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n218), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n194), .A2(G143), .ZN(new_n376));
  INV_X1    g190(.A(G134), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n191), .A2(G128), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT88), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n377), .B1(new_n376), .B2(new_n378), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n382), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT88), .B1(new_n384), .B2(new_n379), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n375), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT9), .B(G234), .ZN(new_n387));
  INV_X1    g201(.A(G217), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n387), .A2(new_n388), .A3(G953), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT90), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT13), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n376), .B1(new_n391), .B2(new_n378), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT13), .B1(new_n191), .B2(G128), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT87), .ZN(new_n394));
  OAI21_X1  g208(.A(G134), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n372), .B(new_n218), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n379), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n390), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n390), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n384), .A2(KEYINPUT88), .A3(new_n379), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n374), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n397), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n404), .A3(new_n282), .ZN(new_n405));
  INV_X1    g219(.A(G478), .ZN(new_n406));
  NOR2_X1   g220(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n410), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n398), .A2(new_n404), .A3(new_n282), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n362), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT92), .B(G952), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(G953), .ZN(new_n418));
  NAND2_X1  g232(.A1(G234), .A2(G237), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(G898), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(G902), .A3(G953), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G214), .B1(G237), .B2(G902), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT81), .ZN(new_n427));
  NOR4_X1   g241(.A1(new_n291), .A2(new_n416), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n377), .B2(G137), .ZN(new_n430));
  INV_X1    g244(.A(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT11), .A3(G134), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n377), .A2(G137), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(new_n432), .A3(new_n303), .A4(new_n433), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(KEYINPUT65), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT65), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n438), .A3(G131), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n209), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n197), .A2(new_n199), .ZN(new_n442));
  INV_X1    g256(.A(new_n433), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n377), .A2(G137), .ZN(new_n444));
  OAI21_X1  g258(.A(G131), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n436), .A3(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n440), .A2(new_n441), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n441), .B1(new_n440), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n253), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n253), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n450), .A3(new_n446), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n300), .A2(G210), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT27), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT26), .B(G101), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n449), .A2(KEYINPUT68), .A3(new_n451), .A4(new_n455), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT31), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n455), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n440), .A2(new_n446), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n253), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n464), .B2(new_n451), .ZN(new_n465));
  INV_X1    g279(.A(new_n451), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(KEYINPUT28), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n461), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT31), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n449), .A2(new_n469), .A3(new_n451), .A4(new_n455), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n460), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(G472), .A2(G902), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT32), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G472), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n465), .A2(new_n467), .A3(new_n461), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT29), .ZN(new_n479));
  INV_X1    g293(.A(new_n449), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n461), .B1(new_n480), .B2(new_n466), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n478), .B2(KEYINPUT29), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n473), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n460), .B2(new_n471), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n476), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G234), .ZN(new_n490));
  OAI21_X1  g304(.A(G217), .B1(new_n490), .B2(G902), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT69), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT73), .ZN(new_n494));
  INV_X1    g308(.A(G110), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n224), .A2(G128), .A3(new_n225), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT70), .B1(new_n496), .B2(KEYINPUT23), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n224), .A2(new_n225), .ZN(new_n499));
  INV_X1    g313(.A(G128), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(KEYINPUT70), .A3(KEYINPUT23), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n495), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(KEYINPUT66), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G128), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n508), .A3(G119), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n496), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT24), .B(G110), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n342), .A2(new_n343), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n318), .A2(new_n329), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n502), .A2(new_n501), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n495), .B(new_n504), .C1(new_n515), .C2(new_n497), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT72), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n510), .A2(new_n517), .A3(new_n511), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n510), .B2(new_n511), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n514), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n494), .B1(new_n513), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n516), .ZN(new_n523));
  INV_X1    g337(.A(new_n514), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n504), .B1(new_n515), .B2(new_n497), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G110), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n510), .A2(new_n511), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n314), .A2(new_n189), .A3(new_n316), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n318), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(KEYINPUT73), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT22), .B(G137), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n297), .A2(G221), .A3(G234), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n522), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n523), .A2(new_n524), .B1(new_n527), .B2(new_n530), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT74), .A3(new_n535), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT74), .B1(new_n538), .B2(new_n535), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n537), .B(new_n282), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n535), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n539), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n548), .A2(KEYINPUT25), .A3(new_n282), .A4(new_n537), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n493), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n548), .ZN(new_n551));
  INV_X1    g365(.A(new_n537), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n492), .A2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G221), .B1(new_n387), .B2(G902), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n209), .A2(new_n254), .A3(new_n223), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT76), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n200), .A2(new_n562), .A3(new_n276), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT77), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n190), .A2(new_n192), .A3(G128), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G128), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n565), .A2(new_n195), .B1(new_n567), .B2(new_n193), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n564), .B1(new_n568), .B2(new_n276), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n193), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n199), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n248), .A2(new_n571), .A3(KEYINPUT77), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n563), .B1(new_n573), .B2(new_n562), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n561), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n437), .A2(new_n439), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(G110), .B(G140), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n297), .A2(G227), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n581), .B(new_n582), .Z(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n561), .A2(new_n574), .A3(new_n578), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n574), .A2(new_n576), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n200), .A2(new_n276), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n573), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(KEYINPUT78), .A3(new_n593), .A4(new_n577), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n593), .B1(new_n576), .B2(KEYINPUT78), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n569), .A2(new_n572), .B1(new_n200), .B2(new_n276), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(new_n576), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n583), .B1(new_n590), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n586), .A2(new_n599), .A3(G469), .ZN(new_n600));
  NAND2_X1  g414(.A1(G469), .A2(G902), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n594), .A2(new_n597), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT80), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n584), .A4(new_n589), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n589), .A2(new_n584), .A3(new_n597), .A4(new_n594), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT80), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n561), .A2(new_n574), .A3(new_n578), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n578), .B1(new_n561), .B2(new_n574), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n583), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n605), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G469), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n282), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n558), .B1(new_n602), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n428), .A2(new_n489), .A3(new_n556), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  OR2_X1    g430(.A1(new_n550), .A2(new_n555), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n460), .B2(new_n471), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n474), .B1(new_n477), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n614), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n288), .A2(KEYINPUT93), .A3(new_n289), .A4(new_n187), .ZN(new_n623));
  INV_X1    g437(.A(new_n427), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT93), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n284), .A2(new_n626), .A3(new_n290), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n398), .A2(new_n404), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n402), .B2(new_n403), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT33), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n398), .A2(new_n404), .A3(new_n631), .A4(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n406), .A2(G902), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n635), .A2(new_n636), .B1(new_n406), .B2(new_n405), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n361), .A2(G475), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n358), .B1(new_n357), .B2(new_n292), .ZN(new_n640));
  INV_X1    g454(.A(new_n292), .ZN(new_n641));
  AOI211_X1 g455(.A(KEYINPUT20), .B(new_n641), .C1(new_n351), .C2(new_n356), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n639), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n628), .A2(new_n425), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n623), .A2(new_n624), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n288), .A2(new_n289), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT93), .B1(new_n650), .B2(new_n188), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n649), .B1(new_n651), .B2(new_n290), .ZN(new_n652));
  INV_X1    g466(.A(new_n425), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n414), .B(new_n639), .C1(new_n640), .C2(new_n642), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT95), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n652), .A2(new_n658), .A3(new_n653), .A4(new_n655), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n621), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NAND2_X1  g476(.A1(new_n522), .A2(new_n532), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT36), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n535), .ZN(new_n665));
  AOI211_X1 g479(.A(KEYINPUT36), .B(new_n536), .C1(new_n522), .C2(new_n532), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n665), .A2(new_n666), .A3(new_n554), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n544), .A2(new_n549), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(new_n492), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n619), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n428), .A2(new_n614), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT96), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  NOR2_X1   g488(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n475), .B(new_n486), .C1(new_n460), .C2(new_n471), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n669), .B1(new_n677), .B2(new_n485), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n421), .B1(new_n679), .B2(new_n424), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n654), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n625), .A2(new_n627), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT97), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n625), .A2(new_n627), .A3(new_n681), .A4(KEYINPUT97), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n678), .A2(new_n684), .A3(new_n614), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT98), .B(G128), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G30));
  XOR2_X1   g502(.A(new_n291), .B(KEYINPUT38), .Z(new_n689));
  NOR2_X1   g503(.A1(new_n362), .A2(new_n415), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n689), .A2(new_n624), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n680), .B(KEYINPUT39), .Z(new_n692));
  AND2_X1   g506(.A1(new_n614), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n458), .A2(new_n459), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n455), .B1(new_n464), .B2(new_n451), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n282), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G472), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n476), .A2(new_n488), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n669), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n691), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NOR3_X1   g517(.A1(new_n362), .A2(new_n637), .A3(new_n680), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n704), .A2(new_n627), .A3(new_n625), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n678), .A2(new_n614), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  AOI21_X1  g521(.A(new_n617), .B1(new_n677), .B2(new_n485), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n611), .A2(new_n282), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT99), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n613), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n709), .A2(KEYINPUT99), .A3(G469), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n558), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n708), .A2(new_n645), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT41), .B(G113), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT100), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n715), .B(new_n717), .ZN(G15));
  NAND2_X1  g532(.A1(new_n712), .A2(new_n713), .ZN(new_n719));
  INV_X1    g533(.A(new_n558), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n489), .A3(new_n556), .A4(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n659), .B2(new_n657), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n227), .ZN(G18));
  NOR2_X1   g537(.A1(new_n416), .A2(new_n425), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n678), .A2(new_n714), .A3(new_n724), .A4(new_n652), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NOR3_X1   g540(.A1(new_n362), .A2(new_n425), .A3(new_n415), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n714), .A2(new_n620), .A3(new_n652), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NAND2_X1  g543(.A1(new_n668), .A2(new_n492), .ZN(new_n730));
  INV_X1    g544(.A(new_n667), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n618), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n487), .B1(new_n733), .B2(G472), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT101), .B1(new_n619), .B2(new_n669), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n704), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n719), .A2(new_n720), .A3(new_n652), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n201), .ZN(G27));
  NAND3_X1  g555(.A1(new_n284), .A2(new_n624), .A3(new_n290), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n284), .A2(KEYINPUT103), .A3(new_n624), .A4(new_n290), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n599), .A2(KEYINPUT102), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n583), .C1(new_n590), .C2(new_n598), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(G469), .A3(new_n586), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n613), .A2(new_n601), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n720), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT104), .B1(new_n746), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n750), .A2(new_n601), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n558), .B1(new_n754), .B2(new_n613), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n756), .A3(new_n744), .A4(new_n745), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n474), .A2(KEYINPUT106), .A3(new_n475), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n487), .B2(KEYINPUT32), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n488), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n484), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n759), .A2(new_n761), .A3(new_n763), .A4(new_n488), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n617), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n758), .A2(new_n767), .A3(new_n704), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n489), .A2(new_n556), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n753), .B2(new_n757), .ZN(new_n770));
  INV_X1    g584(.A(new_n704), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT42), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n768), .A2(KEYINPUT42), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  INV_X1    g589(.A(new_n681), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n769), .B(new_n776), .C1(new_n753), .C2(new_n757), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n377), .ZN(G36));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n586), .B2(new_n599), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n779), .A2(new_n780), .A3(new_n612), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n747), .A2(KEYINPUT45), .A3(new_n586), .A4(new_n749), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n779), .B2(new_n612), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n601), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n601), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n787), .A2(new_n613), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n558), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n638), .A2(new_n362), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n792), .A3(KEYINPUT43), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n643), .B2(new_n637), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n619), .A3(new_n732), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n790), .A2(new_n692), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n797), .A2(KEYINPUT44), .A3(new_n619), .A4(new_n732), .ZN(new_n802));
  INV_X1    g616(.A(new_n746), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT109), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  NOR4_X1   g621(.A1(new_n746), .A2(new_n489), .A3(new_n771), .A4(new_n556), .ZN(new_n808));
  INV_X1    g622(.A(new_n613), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n785), .B2(new_n786), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n788), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT47), .B1(new_n811), .B2(new_n720), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n813), .B(new_n558), .C1(new_n810), .C2(new_n788), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n808), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT110), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n817), .B(new_n808), .C1(new_n812), .C2(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  INV_X1    g634(.A(new_n620), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n793), .A2(new_n421), .A3(new_n796), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT113), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n793), .A2(new_n796), .A3(new_n824), .A4(new_n421), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n803), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n812), .A2(new_n814), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n719), .A2(new_n558), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n719), .A2(new_n720), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n746), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n699), .A2(new_n617), .A3(new_n420), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n638), .A2(new_n643), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n803), .A2(new_n714), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n823), .B2(new_n825), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n736), .A2(new_n737), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n834), .A2(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n689), .A2(new_n831), .A3(new_n624), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n826), .A3(KEYINPUT50), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT50), .B1(new_n840), .B2(new_n826), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT51), .B1(new_n830), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n813), .B1(new_n789), .B2(new_n558), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n811), .A2(KEYINPUT47), .A3(new_n720), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n829), .ZN(new_n848));
  INV_X1    g662(.A(new_n827), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  INV_X1    g665(.A(new_n843), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n841), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n850), .A2(new_n851), .A3(new_n853), .A4(new_n839), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n837), .A2(new_n767), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT48), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n832), .A2(new_n833), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n418), .B1(new_n858), .B2(new_n644), .ZN(new_n859));
  INV_X1    g673(.A(new_n739), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n826), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT114), .B1(new_n855), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n865), .B(new_n862), .C1(new_n845), .C2(new_n854), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n685), .A2(new_n489), .A3(new_n614), .A4(new_n732), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT97), .B1(new_n652), .B2(new_n681), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n738), .A2(new_n739), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n680), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n751), .A2(new_n720), .A3(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n625), .A2(new_n690), .A3(new_n627), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n669), .A4(new_n699), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(KEYINPUT52), .A3(new_n706), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n686), .B(new_n706), .C1(new_n739), .C2(new_n738), .ZN(new_n879));
  INV_X1    g693(.A(new_n876), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n738), .B1(new_n757), .B2(new_n753), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n489), .A2(new_n614), .A3(new_n732), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n362), .A2(new_n415), .A3(new_n873), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n746), .A3(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n777), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n715), .A2(new_n725), .A3(new_n728), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n654), .B1(new_n362), .B2(new_n637), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n427), .B1(new_n284), .B2(new_n290), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n653), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n620), .A2(new_n614), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n615), .A2(new_n892), .A3(new_n671), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n888), .A2(new_n722), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n887), .A2(new_n774), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n868), .B1(new_n882), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n768), .A2(KEYINPUT42), .ZN(new_n898));
  INV_X1    g712(.A(new_n777), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n770), .A2(new_n773), .ZN(new_n900));
  INV_X1    g714(.A(new_n738), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n886), .B1(new_n758), .B2(new_n901), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n879), .B2(new_n880), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n706), .A2(new_n876), .A3(KEYINPUT52), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n872), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n706), .A2(new_n876), .A3(KEYINPUT52), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT111), .B1(new_n871), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n905), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n903), .A2(new_n911), .A3(KEYINPUT53), .A4(new_n894), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n896), .A2(new_n897), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n905), .A2(new_n908), .A3(new_n910), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n868), .B1(new_n914), .B2(new_n895), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n877), .A2(new_n881), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n903), .A2(KEYINPUT53), .A3(new_n916), .A4(new_n894), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n897), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n867), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(G952), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n297), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n689), .ZN(new_n924));
  NOR4_X1   g738(.A1(new_n617), .A2(new_n791), .A3(new_n558), .A4(new_n427), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n677), .A3(new_n698), .A4(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT49), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n719), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n719), .A2(new_n927), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n923), .A2(KEYINPUT115), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT115), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n867), .A2(new_n919), .B1(new_n921), .B2(new_n297), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n931), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(G75));
  NAND2_X1  g751(.A1(new_n921), .A2(G953), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT117), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n282), .B1(new_n896), .B2(new_n912), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n940), .B2(G210), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n287), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n269), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT55), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n939), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n941), .A2(new_n945), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(KEYINPUT116), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(KEYINPUT116), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G51));
  INV_X1    g764(.A(new_n939), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n896), .A2(new_n912), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT54), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n896), .A2(new_n897), .A3(new_n912), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n601), .B(KEYINPUT57), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n611), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n940), .A2(new_n781), .A3(new_n782), .A4(new_n783), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(G54));
  NAND3_X1  g774(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(new_n357), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n951), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT59), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n913), .B2(new_n918), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n635), .B(KEYINPUT118), .Z(new_n968));
  AOI21_X1  g782(.A(new_n951), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n965), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT119), .B1(new_n955), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n897), .B1(new_n896), .B2(new_n912), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT119), .B(new_n970), .C1(new_n913), .C2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n969), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT120), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n969), .B(KEYINPUT120), .C1(new_n971), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(G63));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT121), .Z(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT60), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n896), .B2(new_n912), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n551), .A2(new_n552), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n939), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n665), .A2(new_n666), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n983), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT61), .ZN(G66));
  OR2_X1    g802(.A1(new_n894), .A2(G953), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n422), .A2(new_n211), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n989), .B(KEYINPUT122), .C1(new_n297), .C2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(KEYINPUT122), .B2(new_n989), .ZN(new_n992));
  INV_X1    g806(.A(G898), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n942), .B1(new_n993), .B2(G953), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT123), .Z(new_n995));
  XNOR2_X1  g809(.A(new_n992), .B(new_n995), .ZN(G69));
  AOI21_X1  g810(.A(new_n297), .B1(G227), .B2(G900), .ZN(new_n997));
  INV_X1    g811(.A(new_n879), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n790), .A2(new_n692), .A3(new_n767), .A4(new_n875), .ZN(new_n999));
  AND4_X1   g813(.A1(new_n899), .A2(new_n806), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n1000), .A2(new_n297), .A3(new_n774), .A4(new_n819), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n447), .A2(new_n448), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n320), .A2(new_n322), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1002), .B(new_n1003), .Z(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(G900), .B2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(KEYINPUT127), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1001), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  INV_X1    g825(.A(new_n702), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(new_n879), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n998), .A2(new_n702), .A3(KEYINPUT62), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n708), .A2(new_n803), .A3(new_n693), .A4(new_n889), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT124), .Z(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n801), .B2(new_n805), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n819), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT125), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n819), .A2(new_n1015), .A3(KEYINPUT125), .A4(new_n1018), .ZN(new_n1022));
  AOI21_X1  g836(.A(G953), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1004), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n997), .B1(new_n1010), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT126), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1025), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n997), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n1029), .B(new_n1027), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1026), .B1(new_n1030), .B2(new_n1032), .ZN(G72));
  NOR2_X1   g847(.A1(new_n480), .A2(new_n466), .ZN(new_n1034));
  AND4_X1   g848(.A1(new_n774), .A2(new_n1000), .A3(new_n819), .A4(new_n894), .ZN(new_n1035));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n1034), .B(new_n461), .C1(new_n1035), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n915), .A2(new_n917), .ZN(new_n1040));
  INV_X1    g854(.A(new_n481), .ZN(new_n1041));
  OAI211_X1 g855(.A(new_n1040), .B(new_n1037), .C1(new_n695), .C2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1039), .A2(new_n939), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1021), .A2(new_n894), .A3(new_n1022), .ZN(new_n1044));
  AOI211_X1 g858(.A(new_n1034), .B(new_n461), .C1(new_n1044), .C2(new_n1037), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1043), .A2(new_n1045), .ZN(G57));
endmodule


