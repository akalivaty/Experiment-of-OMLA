

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  BUF_X1 U552 ( .A(n637), .Z(n516) );
  XNOR2_X1 U553 ( .A(n532), .B(n531), .ZN(n906) );
  XNOR2_X2 U554 ( .A(n524), .B(n712), .ZN(n717) );
  AND2_X2 U555 ( .A1(n523), .A2(n522), .ZN(n524) );
  AND2_X2 U556 ( .A1(n546), .A2(n545), .ZN(G164) );
  XNOR2_X1 U557 ( .A(KEYINPUT1), .B(n557), .ZN(n637) );
  BUF_X4 U558 ( .A(n906), .Z(n517) );
  NOR2_X1 U559 ( .A1(n633), .A2(n632), .ZN(n635) );
  NOR2_X1 U560 ( .A1(n623), .A2(n622), .ZN(n660) );
  NAND2_X1 U561 ( .A1(n635), .A2(n634), .ZN(n978) );
  BUF_X1 U562 ( .A(n645), .Z(n683) );
  AND2_X1 U563 ( .A1(n526), .A2(n525), .ZN(G160) );
  AND2_X2 U564 ( .A1(G2104), .A2(G2105), .ZN(n910) );
  AND2_X1 U565 ( .A1(G160), .A2(G40), .ZN(n718) );
  XNOR2_X1 U566 ( .A(n621), .B(KEYINPUT27), .ZN(n623) );
  NOR2_X1 U567 ( .A1(n675), .A2(n605), .ZN(n607) );
  INV_X1 U568 ( .A(KEYINPUT100), .ZN(n672) );
  NOR2_X1 U569 ( .A1(n711), .A2(n520), .ZN(n522) );
  INV_X1 U570 ( .A(KEYINPUT108), .ZN(n712) );
  INV_X1 U571 ( .A(KEYINPUT109), .ZN(n748) );
  AND2_X1 U572 ( .A1(G125), .A2(n912), .ZN(n518) );
  AND2_X1 U573 ( .A1(n710), .A2(n528), .ZN(n519) );
  AND2_X1 U574 ( .A1(n710), .A2(KEYINPUT33), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n521), .A2(n993), .ZN(n698) );
  NAND2_X1 U576 ( .A1(n694), .A2(n695), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n521), .A2(n702), .ZN(n703) );
  NAND2_X1 U578 ( .A1(n700), .A2(n519), .ZN(n523) );
  NOR2_X1 U579 ( .A1(n538), .A2(n518), .ZN(n525) );
  XNOR2_X1 U580 ( .A(n527), .B(KEYINPUT67), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n534), .A2(n535), .ZN(n527) );
  AND2_X1 U582 ( .A1(n536), .A2(G2104), .ZN(n904) );
  NOR2_X1 U583 ( .A1(G2104), .A2(n536), .ZN(n912) );
  AND2_X1 U584 ( .A1(n680), .A2(n677), .ZN(n678) );
  NOR2_X1 U585 ( .A1(n681), .A2(n699), .ZN(n528) );
  XOR2_X1 U586 ( .A(KEYINPUT74), .B(n640), .Z(n529) );
  AND2_X1 U587 ( .A1(G8), .A2(n675), .ZN(n530) );
  NOR2_X1 U588 ( .A1(n676), .A2(n530), .ZN(n677) );
  XNOR2_X1 U589 ( .A(n691), .B(KEYINPUT103), .ZN(n692) );
  INV_X1 U590 ( .A(KEYINPUT105), .ZN(n697) );
  NAND2_X1 U591 ( .A1(G8), .A2(n645), .ZN(n681) );
  AND2_X1 U592 ( .A1(n555), .A2(G651), .ZN(n556) );
  INV_X1 U593 ( .A(G651), .ZN(n548) );
  INV_X1 U594 ( .A(KEYINPUT17), .ZN(n531) );
  NOR2_X2 U595 ( .A1(n582), .A2(n548), .ZN(n811) );
  XOR2_X1 U596 ( .A(KEYINPUT70), .B(n571), .Z(G301) );
  NAND2_X1 U597 ( .A1(n906), .A2(G137), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n910), .A2(G113), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT66), .ZN(n534) );
  INV_X1 U600 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U601 ( .A1(G101), .A2(n904), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT23), .B(n537), .ZN(n538) );
  NAND2_X1 U603 ( .A1(G138), .A2(n517), .ZN(n540) );
  NAND2_X1 U604 ( .A1(G102), .A2(n904), .ZN(n539) );
  NAND2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n541), .B(KEYINPUT91), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G126), .A2(n912), .ZN(n544) );
  NAND2_X1 U608 ( .A1(G114), .A2(n910), .ZN(n542) );
  XNOR2_X1 U609 ( .A(KEYINPUT90), .B(n542), .ZN(n543) );
  AND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U611 ( .A1(G651), .A2(G543), .ZN(n810) );
  NAND2_X1 U612 ( .A1(n810), .A2(G89), .ZN(n547) );
  XNOR2_X1 U613 ( .A(KEYINPUT4), .B(n547), .ZN(n551) );
  XOR2_X1 U614 ( .A(G543), .B(KEYINPUT0), .Z(n582) );
  NAND2_X1 U615 ( .A1(n811), .A2(G76), .ZN(n549) );
  XOR2_X1 U616 ( .A(KEYINPUT75), .B(n549), .Z(n550) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(KEYINPUT5), .ZN(n562) );
  NOR2_X1 U619 ( .A1(G651), .A2(n582), .ZN(n553) );
  XOR2_X2 U620 ( .A(KEYINPUT65), .B(n553), .Z(n807) );
  NAND2_X1 U621 ( .A1(n807), .A2(G51), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n554), .B(KEYINPUT76), .ZN(n559) );
  INV_X1 U623 ( .A(G543), .ZN(n555) );
  XOR2_X1 U624 ( .A(KEYINPUT68), .B(n556), .Z(n557) );
  NAND2_X1 U625 ( .A1(G63), .A2(n516), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT6), .B(n560), .Z(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U630 ( .A1(n807), .A2(G52), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G64), .A2(n516), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G90), .A2(n810), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G77), .A2(n811), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U638 ( .A(G301), .ZN(G171) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G88), .A2(n810), .ZN(n573) );
  NAND2_X1 U641 ( .A1(G75), .A2(n811), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G62), .A2(n516), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT84), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G50), .A2(n807), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U647 ( .A1(n578), .A2(n577), .ZN(G166) );
  INV_X1 U648 ( .A(G166), .ZN(G303) );
  NAND2_X1 U649 ( .A1(G49), .A2(n807), .ZN(n580) );
  NAND2_X1 U650 ( .A1(G74), .A2(G651), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U652 ( .A(KEYINPUT80), .B(n581), .Z(n586) );
  NAND2_X1 U653 ( .A1(G87), .A2(n582), .ZN(n583) );
  XNOR2_X1 U654 ( .A(KEYINPUT81), .B(n583), .ZN(n584) );
  NOR2_X1 U655 ( .A1(n516), .A2(n584), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U657 ( .A1(G73), .A2(n811), .ZN(n587) );
  XOR2_X1 U658 ( .A(KEYINPUT2), .B(n587), .Z(n593) );
  NAND2_X1 U659 ( .A1(n810), .A2(G86), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n588), .B(KEYINPUT82), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G61), .A2(n516), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U663 ( .A(KEYINPUT83), .B(n591), .Z(n592) );
  NOR2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n807), .A2(G48), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(G305) );
  NAND2_X1 U667 ( .A1(G85), .A2(n810), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G72), .A2(n811), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G60), .A2(n516), .ZN(n598) );
  XNOR2_X1 U671 ( .A(KEYINPUT69), .B(n598), .ZN(n599) );
  NOR2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n807), .A2(G47), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n602), .A2(n601), .ZN(G290) );
  NOR2_X2 U675 ( .A1(G164), .A2(G1384), .ZN(n720) );
  NAND2_X2 U676 ( .A1(n718), .A2(n720), .ZN(n645) );
  NOR2_X1 U677 ( .A1(G2084), .A2(n683), .ZN(n675) );
  NOR2_X1 U678 ( .A1(G1966), .A2(n681), .ZN(n604) );
  INV_X1 U679 ( .A(KEYINPUT96), .ZN(n603) );
  XNOR2_X1 U680 ( .A(n604), .B(n603), .ZN(n674) );
  NAND2_X1 U681 ( .A1(n674), .A2(G8), .ZN(n605) );
  XNOR2_X1 U682 ( .A(KEYINPUT99), .B(KEYINPUT30), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n607), .B(n606), .ZN(n608) );
  NOR2_X1 U684 ( .A1(G168), .A2(n608), .ZN(n612) );
  XNOR2_X1 U685 ( .A(G2078), .B(KEYINPUT25), .ZN(n959) );
  NOR2_X1 U686 ( .A1(n683), .A2(n959), .ZN(n610) );
  AND2_X1 U687 ( .A1(n683), .A2(G1961), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n666) );
  NOR2_X1 U689 ( .A1(n666), .A2(G171), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U691 ( .A(KEYINPUT31), .B(n613), .ZN(n671) );
  NAND2_X1 U692 ( .A1(n807), .A2(G53), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G65), .A2(n516), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G91), .A2(n810), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G78), .A2(n811), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n982) );
  INV_X1 U699 ( .A(n645), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n620), .A2(G2072), .ZN(n621) );
  AND2_X1 U701 ( .A1(G1956), .A2(n683), .ZN(n622) );
  NOR2_X1 U702 ( .A1(n982), .A2(n660), .ZN(n625) );
  XNOR2_X1 U703 ( .A(KEYINPUT97), .B(KEYINPUT28), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n625), .B(n624), .ZN(n664) );
  XNOR2_X1 U705 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n651) );
  NOR2_X1 U706 ( .A1(G1996), .A2(n651), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n810), .A2(G81), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n626), .B(KEYINPUT12), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G68), .A2(n811), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U711 ( .A(KEYINPUT13), .B(n629), .Z(n633) );
  NAND2_X1 U712 ( .A1(n637), .A2(G56), .ZN(n630) );
  XNOR2_X1 U713 ( .A(n630), .B(KEYINPUT73), .ZN(n631) );
  XNOR2_X1 U714 ( .A(n631), .B(KEYINPUT14), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n807), .A2(G43), .ZN(n634) );
  NOR2_X1 U716 ( .A1(n636), .A2(n978), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n807), .A2(G54), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n810), .A2(G92), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G66), .A2(n516), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n811), .A2(G79), .ZN(n640) );
  NOR2_X1 U722 ( .A1(n641), .A2(n529), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U724 ( .A(KEYINPUT15), .B(n644), .Z(n782) );
  NAND2_X1 U725 ( .A1(G1348), .A2(n645), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G2067), .A2(n620), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n782), .A2(n657), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n656) );
  INV_X1 U730 ( .A(G1341), .ZN(n979) );
  NAND2_X1 U731 ( .A1(n979), .A2(n651), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n650), .A2(n683), .ZN(n654) );
  AND2_X1 U733 ( .A1(G1996), .A2(n620), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U736 ( .A1(n656), .A2(n655), .ZN(n659) );
  NOR2_X1 U737 ( .A1(n657), .A2(n782), .ZN(n658) );
  NOR2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U739 ( .A1(n982), .A2(n660), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n665), .B(KEYINPUT29), .ZN(n668) );
  AND2_X1 U743 ( .A1(n666), .A2(G171), .ZN(n667) );
  NOR2_X1 U744 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n669), .B(KEYINPUT98), .ZN(n670) );
  NOR2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n673) );
  XNOR2_X1 U747 ( .A(n673), .B(n672), .ZN(n680) );
  INV_X1 U748 ( .A(n674), .ZN(n676) );
  XNOR2_X1 U749 ( .A(n678), .B(KEYINPUT101), .ZN(n695) );
  AND2_X1 U750 ( .A1(G286), .A2(G8), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n690) );
  INV_X1 U752 ( .A(G8), .ZN(n688) );
  NOR2_X1 U753 ( .A1(G1971), .A2(n681), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n682), .B(KEYINPUT102), .ZN(n685) );
  NOR2_X1 U755 ( .A1(n683), .A2(G2090), .ZN(n684) );
  NOR2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U757 ( .A1(n686), .A2(G303), .ZN(n687) );
  OR2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n693) );
  XNOR2_X1 U760 ( .A(KEYINPUT32), .B(KEYINPUT104), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(G1976), .A2(G288), .ZN(n704) );
  NOR2_X1 U763 ( .A1(G1971), .A2(G303), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n704), .A2(n696), .ZN(n993) );
  XNOR2_X1 U765 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U766 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U767 ( .A(n980), .ZN(n699) );
  NOR2_X1 U768 ( .A1(G2090), .A2(G303), .ZN(n701) );
  NAND2_X1 U769 ( .A1(G8), .A2(n701), .ZN(n702) );
  AND2_X1 U770 ( .A1(n703), .A2(n681), .ZN(n711) );
  NAND2_X1 U771 ( .A1(KEYINPUT33), .A2(n704), .ZN(n705) );
  XNOR2_X1 U772 ( .A(KEYINPUT106), .B(n705), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n681), .A2(n706), .ZN(n707) );
  XOR2_X1 U774 ( .A(KEYINPUT107), .B(n707), .Z(n709) );
  XOR2_X1 U775 ( .A(G1981), .B(G305), .Z(n997) );
  INV_X1 U776 ( .A(n997), .ZN(n708) );
  NOR2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U778 ( .A1(G1981), .A2(G305), .ZN(n713) );
  XNOR2_X1 U779 ( .A(n713), .B(KEYINPUT95), .ZN(n714) );
  XNOR2_X1 U780 ( .A(n714), .B(KEYINPUT24), .ZN(n715) );
  NOR2_X1 U781 ( .A1(n681), .A2(n715), .ZN(n716) );
  NOR2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n747) );
  INV_X1 U783 ( .A(n718), .ZN(n719) );
  NOR2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n762) );
  XNOR2_X1 U785 ( .A(G2067), .B(KEYINPUT37), .ZN(n760) );
  NAND2_X1 U786 ( .A1(n904), .A2(G104), .ZN(n721) );
  XNOR2_X1 U787 ( .A(n721), .B(KEYINPUT92), .ZN(n723) );
  NAND2_X1 U788 ( .A1(G140), .A2(n517), .ZN(n722) );
  NAND2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U790 ( .A(KEYINPUT34), .B(n724), .ZN(n729) );
  NAND2_X1 U791 ( .A1(G116), .A2(n910), .ZN(n726) );
  NAND2_X1 U792 ( .A1(G128), .A2(n912), .ZN(n725) );
  NAND2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U794 ( .A(KEYINPUT35), .B(n727), .Z(n728) );
  NOR2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U796 ( .A(KEYINPUT36), .B(n730), .ZN(n900) );
  NOR2_X1 U797 ( .A1(n760), .A2(n900), .ZN(n942) );
  NAND2_X1 U798 ( .A1(n762), .A2(n942), .ZN(n758) );
  NAND2_X1 U799 ( .A1(G141), .A2(n517), .ZN(n732) );
  NAND2_X1 U800 ( .A1(G117), .A2(n910), .ZN(n731) );
  NAND2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n735) );
  NAND2_X1 U802 ( .A1(n904), .A2(G105), .ZN(n733) );
  XOR2_X1 U803 ( .A(KEYINPUT38), .B(n733), .Z(n734) );
  NOR2_X1 U804 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U805 ( .A1(n912), .A2(G129), .ZN(n736) );
  NAND2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n888) );
  AND2_X1 U807 ( .A1(n888), .A2(G1996), .ZN(n938) );
  NAND2_X1 U808 ( .A1(G131), .A2(n517), .ZN(n739) );
  NAND2_X1 U809 ( .A1(G95), .A2(n904), .ZN(n738) );
  NAND2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n743) );
  NAND2_X1 U811 ( .A1(G107), .A2(n910), .ZN(n741) );
  NAND2_X1 U812 ( .A1(G119), .A2(n912), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U814 ( .A1(n743), .A2(n742), .ZN(n884) );
  XNOR2_X1 U815 ( .A(KEYINPUT93), .B(G1991), .ZN(n960) );
  NOR2_X1 U816 ( .A1(n884), .A2(n960), .ZN(n932) );
  OR2_X1 U817 ( .A1(n938), .A2(n932), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n744), .A2(n762), .ZN(n752) );
  NAND2_X1 U819 ( .A1(n758), .A2(n752), .ZN(n745) );
  XNOR2_X1 U820 ( .A(KEYINPUT94), .B(n745), .ZN(n746) );
  NOR2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U822 ( .A(n749), .B(n748), .ZN(n751) );
  XNOR2_X1 U823 ( .A(G1986), .B(G290), .ZN(n986) );
  NAND2_X1 U824 ( .A1(n986), .A2(n762), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n765) );
  NOR2_X1 U826 ( .A1(G1996), .A2(n888), .ZN(n929) );
  INV_X1 U827 ( .A(n752), .ZN(n755) );
  AND2_X1 U828 ( .A1(n960), .A2(n884), .ZN(n934) );
  NOR2_X1 U829 ( .A1(G1986), .A2(G290), .ZN(n753) );
  NOR2_X1 U830 ( .A1(n934), .A2(n753), .ZN(n754) );
  NOR2_X1 U831 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U832 ( .A1(n929), .A2(n756), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n757), .B(KEYINPUT39), .ZN(n759) );
  NAND2_X1 U834 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U835 ( .A1(n760), .A2(n900), .ZN(n943) );
  NAND2_X1 U836 ( .A1(n761), .A2(n943), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U838 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n766), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U840 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n768) );
  XNOR2_X1 U841 ( .A(G2446), .B(G2451), .ZN(n767) );
  XNOR2_X1 U842 ( .A(n768), .B(n767), .ZN(n772) );
  XOR2_X1 U843 ( .A(G2435), .B(G2438), .Z(n770) );
  XNOR2_X1 U844 ( .A(G2454), .B(KEYINPUT110), .ZN(n769) );
  XNOR2_X1 U845 ( .A(n770), .B(n769), .ZN(n771) );
  XOR2_X1 U846 ( .A(n772), .B(n771), .Z(n774) );
  XNOR2_X1 U847 ( .A(G2443), .B(G2427), .ZN(n773) );
  XNOR2_X1 U848 ( .A(n774), .B(n773), .ZN(n777) );
  XNOR2_X1 U849 ( .A(G1348), .B(G2430), .ZN(n775) );
  XNOR2_X1 U850 ( .A(n775), .B(n979), .ZN(n776) );
  XOR2_X1 U851 ( .A(n777), .B(n776), .Z(n778) );
  AND2_X1 U852 ( .A1(G14), .A2(n778), .ZN(G401) );
  AND2_X1 U853 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  INV_X1 U855 ( .A(G132), .ZN(G219) );
  NAND2_X1 U856 ( .A1(G7), .A2(G661), .ZN(n779) );
  XNOR2_X1 U857 ( .A(n779), .B(KEYINPUT72), .ZN(n780) );
  XNOR2_X1 U858 ( .A(KEYINPUT10), .B(n780), .ZN(G223) );
  INV_X1 U859 ( .A(G223), .ZN(n846) );
  NAND2_X1 U860 ( .A1(n846), .A2(G567), .ZN(n781) );
  XOR2_X1 U861 ( .A(KEYINPUT11), .B(n781), .Z(G234) );
  INV_X1 U862 ( .A(G860), .ZN(n788) );
  OR2_X1 U863 ( .A1(n978), .A2(n788), .ZN(G153) );
  NAND2_X1 U864 ( .A1(G301), .A2(G868), .ZN(n784) );
  INV_X1 U865 ( .A(n782), .ZN(n805) );
  INV_X1 U866 ( .A(n805), .ZN(n987) );
  INV_X1 U867 ( .A(G868), .ZN(n827) );
  NAND2_X1 U868 ( .A1(n987), .A2(n827), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(G284) );
  NAND2_X1 U870 ( .A1(n982), .A2(n827), .ZN(n785) );
  XNOR2_X1 U871 ( .A(n785), .B(KEYINPUT77), .ZN(n787) );
  NOR2_X1 U872 ( .A1(n827), .A2(G286), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(G297) );
  NAND2_X1 U874 ( .A1(n788), .A2(G559), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n789), .A2(n805), .ZN(n790) );
  XNOR2_X1 U876 ( .A(n790), .B(KEYINPUT78), .ZN(n791) );
  XNOR2_X1 U877 ( .A(KEYINPUT16), .B(n791), .ZN(G148) );
  NOR2_X1 U878 ( .A1(G868), .A2(n978), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G868), .A2(n805), .ZN(n792) );
  NOR2_X1 U880 ( .A1(G559), .A2(n792), .ZN(n793) );
  NOR2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U882 ( .A(KEYINPUT79), .B(n795), .Z(G282) );
  NAND2_X1 U883 ( .A1(G123), .A2(n912), .ZN(n796) );
  XNOR2_X1 U884 ( .A(n796), .B(KEYINPUT18), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n910), .A2(G111), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U887 ( .A1(G135), .A2(n517), .ZN(n800) );
  NAND2_X1 U888 ( .A1(G99), .A2(n904), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n931) );
  XNOR2_X1 U891 ( .A(G2096), .B(n931), .ZN(n804) );
  INV_X1 U892 ( .A(G2100), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n804), .A2(n803), .ZN(G156) );
  NAND2_X1 U894 ( .A1(n805), .A2(G559), .ZN(n824) );
  XNOR2_X1 U895 ( .A(n978), .B(n824), .ZN(n806) );
  NOR2_X1 U896 ( .A1(n806), .A2(G860), .ZN(n816) );
  NAND2_X1 U897 ( .A1(n807), .A2(G55), .ZN(n809) );
  NAND2_X1 U898 ( .A1(G67), .A2(n516), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G93), .A2(n810), .ZN(n813) );
  NAND2_X1 U901 ( .A1(G80), .A2(n811), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n826) );
  XNOR2_X1 U904 ( .A(n816), .B(n826), .ZN(G145) );
  XOR2_X1 U905 ( .A(G290), .B(n978), .Z(n817) );
  XNOR2_X1 U906 ( .A(G288), .B(n817), .ZN(n821) );
  XNOR2_X1 U907 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n819) );
  XNOR2_X1 U908 ( .A(G305), .B(n982), .ZN(n818) );
  XNOR2_X1 U909 ( .A(n819), .B(n818), .ZN(n820) );
  XOR2_X1 U910 ( .A(n821), .B(n820), .Z(n823) );
  XNOR2_X1 U911 ( .A(G166), .B(n826), .ZN(n822) );
  XNOR2_X1 U912 ( .A(n823), .B(n822), .ZN(n853) );
  XNOR2_X1 U913 ( .A(n824), .B(n853), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n825), .A2(G868), .ZN(n829) );
  NAND2_X1 U915 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U916 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U917 ( .A(KEYINPUT86), .B(n830), .Z(G295) );
  NAND2_X1 U918 ( .A1(G2084), .A2(G2078), .ZN(n831) );
  XOR2_X1 U919 ( .A(KEYINPUT20), .B(n831), .Z(n832) );
  NAND2_X1 U920 ( .A1(G2090), .A2(n832), .ZN(n833) );
  XNOR2_X1 U921 ( .A(KEYINPUT21), .B(n833), .ZN(n834) );
  NAND2_X1 U922 ( .A1(n834), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U923 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  XNOR2_X1 U924 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U925 ( .A1(G219), .A2(G220), .ZN(n836) );
  XNOR2_X1 U926 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n835) );
  XNOR2_X1 U927 ( .A(n836), .B(n835), .ZN(n837) );
  NOR2_X1 U928 ( .A1(n837), .A2(G218), .ZN(n838) );
  NAND2_X1 U929 ( .A1(G96), .A2(n838), .ZN(n839) );
  XNOR2_X1 U930 ( .A(KEYINPUT88), .B(n839), .ZN(n852) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n852), .ZN(n844) );
  NAND2_X1 U932 ( .A1(G120), .A2(G108), .ZN(n840) );
  NOR2_X1 U933 ( .A1(G237), .A2(n840), .ZN(n841) );
  NAND2_X1 U934 ( .A1(G69), .A2(n841), .ZN(n851) );
  NAND2_X1 U935 ( .A1(G567), .A2(n851), .ZN(n842) );
  XOR2_X1 U936 ( .A(KEYINPUT89), .B(n842), .Z(n843) );
  NAND2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n927) );
  NAND2_X1 U938 ( .A1(G661), .A2(G483), .ZN(n845) );
  NOR2_X1 U939 ( .A1(n927), .A2(n845), .ZN(n850) );
  NAND2_X1 U940 ( .A1(n850), .A2(G36), .ZN(G176) );
  NAND2_X1 U941 ( .A1(G2106), .A2(n846), .ZN(G217) );
  AND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U943 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n848) );
  XOR2_X1 U945 ( .A(KEYINPUT113), .B(n848), .Z(n849) );
  NAND2_X1 U946 ( .A1(n850), .A2(n849), .ZN(G188) );
  XNOR2_X1 U947 ( .A(G108), .B(KEYINPUT123), .ZN(G238) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  NOR2_X1 U951 ( .A1(n852), .A2(n851), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U953 ( .A(n987), .B(n853), .ZN(n855) );
  XNOR2_X1 U954 ( .A(G286), .B(G301), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  NOR2_X1 U956 ( .A1(G37), .A2(n856), .ZN(G397) );
  XOR2_X1 U957 ( .A(KEYINPUT116), .B(G2678), .Z(n858) );
  XNOR2_X1 U958 ( .A(KEYINPUT43), .B(G2096), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n859), .B(KEYINPUT115), .Z(n861) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2084), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U963 ( .A(G2100), .B(G2072), .Z(n863) );
  XNOR2_X1 U964 ( .A(G2090), .B(G2078), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U966 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U967 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(G227) );
  XOR2_X1 U969 ( .A(G1976), .B(G1956), .Z(n869) );
  XNOR2_X1 U970 ( .A(G1986), .B(G1971), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U972 ( .A(n870), .B(G2474), .Z(n872) );
  XNOR2_X1 U973 ( .A(G1996), .B(G1991), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U975 ( .A(KEYINPUT41), .B(G1961), .Z(n874) );
  XNOR2_X1 U976 ( .A(G1981), .B(G1966), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(G229) );
  NAND2_X1 U979 ( .A1(G124), .A2(n912), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n877), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n910), .A2(G112), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G136), .A2(n517), .ZN(n881) );
  NAND2_X1 U984 ( .A1(G100), .A2(n904), .ZN(n880) );
  NAND2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U986 ( .A1(n883), .A2(n882), .ZN(G162) );
  XOR2_X1 U987 ( .A(KEYINPUT48), .B(KEYINPUT121), .Z(n886) );
  XNOR2_X1 U988 ( .A(n884), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U990 ( .A(n887), .B(n931), .Z(n890) );
  XOR2_X1 U991 ( .A(n888), .B(G162), .Z(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U993 ( .A(G164), .B(n891), .ZN(n903) );
  NAND2_X1 U994 ( .A1(G118), .A2(n910), .ZN(n893) );
  NAND2_X1 U995 ( .A1(G130), .A2(n912), .ZN(n892) );
  NAND2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n899) );
  NAND2_X1 U997 ( .A1(n517), .A2(G142), .ZN(n894) );
  XOR2_X1 U998 ( .A(KEYINPUT117), .B(n894), .Z(n896) );
  NAND2_X1 U999 ( .A1(n904), .A2(G106), .ZN(n895) );
  NAND2_X1 U1000 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U1001 ( .A(n897), .B(KEYINPUT45), .Z(n898) );
  NOR2_X1 U1002 ( .A1(n899), .A2(n898), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n919) );
  NAND2_X1 U1005 ( .A1(n904), .A2(G103), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n905), .B(KEYINPUT118), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(G139), .A2(n517), .ZN(n907) );
  NAND2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1009 ( .A(KEYINPUT119), .B(n909), .Z(n917) );
  NAND2_X1 U1010 ( .A1(n910), .A2(G115), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n911), .B(KEYINPUT120), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(G127), .A2(n912), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1014 ( .A(KEYINPUT47), .B(n915), .Z(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n947) );
  XOR2_X1 U1016 ( .A(n947), .B(G160), .Z(n918) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n920), .ZN(G395) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n927), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(G397), .A2(n922), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n925), .A2(G395), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n926), .B(KEYINPUT122), .ZN(G308) );
  INV_X1 U1026 ( .A(G308), .ZN(G225) );
  INV_X1 U1027 ( .A(n982), .ZN(G299) );
  INV_X1 U1028 ( .A(n927), .ZN(G319) );
  INV_X1 U1029 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n930), .Z(n940) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n936) );
  XOR2_X1 U1034 ( .A(G160), .B(G2084), .Z(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(KEYINPUT124), .B(n945), .ZN(n952) );
  XNOR2_X1 U1042 ( .A(G164), .B(G2078), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(KEYINPUT125), .ZN(n949) );
  XOR2_X1 U1044 ( .A(G2072), .B(n947), .Z(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1046 ( .A(KEYINPUT50), .B(n950), .Z(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n953), .ZN(n954) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n974) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n974), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n955), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1052 ( .A(G2090), .B(G35), .ZN(n969) );
  XOR2_X1 U1053 ( .A(G2067), .B(G26), .Z(n956) );
  NAND2_X1 U1054 ( .A1(n956), .A2(G28), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(G1996), .B(G32), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(G33), .B(G2072), .ZN(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n964) );
  XOR2_X1 U1058 ( .A(n959), .B(G27), .Z(n962) );
  XOR2_X1 U1059 ( .A(n960), .B(G25), .Z(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n967), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n970) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n970), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n974), .B(n973), .ZN(n976) );
  INV_X1 U1069 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n977), .ZN(n1030) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .ZN(n1003) );
  XNOR2_X1 U1073 ( .A(n979), .B(n978), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n995) );
  XNOR2_X1 U1075 ( .A(G1956), .B(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(G1971), .A2(G303), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n989) );
  XOR2_X1 U1079 ( .A(G1348), .B(n987), .Z(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G1961), .B(G301), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(KEYINPUT126), .B(n996), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G168), .B(G1966), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(KEYINPUT57), .B(n999), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1028) );
  INV_X1 U1091 ( .A(G16), .ZN(n1026) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G5), .B(G1961), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1016) );
  XNOR2_X1 U1095 ( .A(KEYINPUT59), .B(G1348), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G4), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G20), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(G1341), .B(G19), .ZN(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(KEYINPUT127), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1014), .Z(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(G1986), .B(G24), .Z(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

