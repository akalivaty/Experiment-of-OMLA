//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT34), .ZN(new_n205));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT69), .ZN(new_n208));
  XOR2_X1   g007(.A(G113gat), .B(G120gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(G169gat), .A3(G176gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n224), .A2(new_n226), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(G183gat), .B(G190gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT66), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n232), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G190gat), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n236), .B1(new_n241), .B2(KEYINPUT24), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n227), .A2(new_n229), .A3(new_n226), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .A4(new_n224), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n223), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT64), .B(G176gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n246), .B(new_n228), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n219), .B1(new_n249), .B2(new_n234), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n235), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n228), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n222), .B2(KEYINPUT26), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n222), .A2(KEYINPUT26), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n237), .A2(KEYINPUT27), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT27), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G183gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n239), .B1(new_n262), .B2(KEYINPUT28), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT68), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n265));
  AOI21_X1  g064(.A(G190gat), .B1(new_n265), .B2(KEYINPUT67), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n258), .A4(new_n260), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n270), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n257), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n218), .B1(new_n251), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n257), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n264), .A2(new_n272), .A3(new_n268), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n264), .B2(new_n268), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n235), .A2(new_n245), .A3(new_n250), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n280), .A3(new_n217), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G227gat), .ZN(new_n283));
  INV_X1    g082(.A(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n205), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  AOI211_X1 g086(.A(KEYINPUT34), .B(new_n285), .C1(new_n275), .C2(new_n281), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n275), .A2(new_n285), .A3(new_n281), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT32), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT33), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G71gat), .B(G99gat), .Z(new_n294));
  XNOR2_X1  g093(.A(G15gat), .B(G43gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n292), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n298), .B2(new_n296), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n290), .A2(KEYINPUT32), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n289), .A2(new_n297), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n287), .ZN(new_n303));
  INV_X1    g102(.A(new_n288), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n297), .A2(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n204), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n302), .A2(new_n305), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT36), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n310), .B(new_n204), .C1(new_n302), .C2(new_n305), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G226gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(new_n284), .ZN(new_n314));
  OAI22_X1  g113(.A1(new_n251), .A2(new_n274), .B1(KEYINPUT29), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n314), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n279), .A2(new_n280), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  AND2_X1   g117(.A1(G211gat), .A2(G218gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(KEYINPUT22), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G211gat), .B(G218gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n315), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n315), .A2(KEYINPUT75), .A3(new_n317), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n322), .B(KEYINPUT74), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n315), .B2(new_n317), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  NAND3_X1  g133(.A1(new_n328), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT30), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n334), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n336), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI211_X1 g139(.A(new_n340), .B(new_n330), .C1(new_n326), .C2(new_n327), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n328), .A2(new_n331), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n334), .B(KEYINPUT76), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT0), .ZN(new_n349));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(KEYINPUT77), .ZN(new_n359));
  INV_X1    g158(.A(G141gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(G148gat), .ZN(new_n361));
  INV_X1    g160(.A(G148gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(G141gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n357), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365));
  OAI22_X1  g164(.A1(new_n361), .A2(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n358), .A2(KEYINPUT77), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n370));
  INV_X1    g169(.A(G155gat), .ZN(new_n371));
  INV_X1    g170(.A(G162gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G162gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n371), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n370), .B1(new_n376), .B2(new_n365), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT80), .B(G162gat), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT81), .B(KEYINPUT2), .C1(new_n378), .C2(new_n371), .ZN(new_n379));
  OR2_X1    g178(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(G148gat), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n361), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n356), .A2(new_n385), .A3(new_n357), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT79), .B1(new_n364), .B2(new_n355), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n377), .A2(new_n379), .A3(new_n384), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT82), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n386), .A2(new_n387), .B1(new_n382), .B2(new_n383), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n377), .A3(new_n392), .A4(new_n379), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n369), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n218), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n369), .B(new_n217), .C1(new_n390), .C2(new_n393), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n354), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT5), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n217), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT3), .B(new_n369), .C1(new_n390), .C2(new_n393), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n353), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n396), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n394), .A2(new_n218), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT4), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n394), .A2(new_n404), .A3(new_n218), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n398), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n390), .A2(new_n393), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n368), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n218), .B1(new_n413), .B2(KEYINPUT3), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n399), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n354), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT5), .B1(new_n408), .B2(new_n409), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n352), .B1(new_n411), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n404), .B1(new_n394), .B2(new_n218), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT83), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n410), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n398), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n418), .A3(new_n351), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n351), .B1(new_n425), .B2(new_n418), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n347), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n322), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n399), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n413), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n433), .ZN(new_n440));
  INV_X1    g239(.A(new_n329), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n435), .ZN(new_n442));
  OAI21_X1  g241(.A(G22gat), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n444));
  INV_X1    g243(.A(new_n440), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n435), .A2(new_n441), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT29), .B1(new_n394), .B2(new_n399), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n438), .B1(new_n448), .B2(new_n323), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n432), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G78gat), .B(G106gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT31), .B(G50gat), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n453), .B(new_n454), .Z(new_n455));
  NAND4_X1  g254(.A1(new_n443), .A2(new_n444), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n458), .A2(new_n455), .B1(new_n443), .B2(new_n452), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n312), .B1(new_n431), .B2(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(new_n351), .B(KEYINPUT85), .Z(new_n462));
  AND3_X1   g261(.A1(new_n394), .A2(new_n404), .A3(new_n218), .ZN(new_n463));
  OAI22_X1  g262(.A1(new_n463), .A2(new_n421), .B1(new_n400), .B2(new_n401), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n354), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n408), .A2(new_n409), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n414), .A2(new_n415), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n353), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n395), .A2(new_n396), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT39), .B1(new_n470), .B2(new_n354), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n462), .B(new_n466), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n347), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n423), .A2(new_n424), .B1(new_n416), .B2(new_n417), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n472), .A2(new_n473), .B1(new_n476), .B2(new_n462), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT86), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n344), .B1(new_n328), .B2(new_n331), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n341), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n480), .A2(new_n337), .B1(new_n472), .B2(new_n473), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n472), .A2(new_n473), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n425), .A2(new_n418), .ZN(new_n484));
  INV_X1    g283(.A(new_n462), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n443), .A2(new_n452), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n445), .A2(new_n446), .B1(new_n449), .B2(new_n432), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n444), .B1(new_n490), .B2(new_n451), .ZN(new_n491));
  INV_X1    g290(.A(new_n455), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n456), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT6), .B1(new_n476), .B2(new_n351), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n495), .A2(new_n486), .B1(KEYINPUT6), .B2(new_n429), .ZN(new_n496));
  AOI211_X1 g295(.A(KEYINPUT37), .B(new_n330), .C1(new_n326), .C2(new_n327), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n344), .A2(KEYINPUT38), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n315), .A2(new_n317), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT37), .B1(new_n499), .B2(new_n329), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n322), .B1(new_n315), .B2(new_n317), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n335), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n334), .B1(new_n343), .B2(KEYINPUT37), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(KEYINPUT37), .B2(new_n343), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n505), .B2(KEYINPUT38), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n494), .B1(new_n496), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n461), .B1(new_n488), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n456), .A3(new_n308), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n431), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n347), .A2(KEYINPUT35), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n511), .A2(KEYINPUT35), .B1(new_n513), .B2(new_n510), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT87), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n488), .A2(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n428), .A2(new_n430), .ZN(new_n517));
  INV_X1    g316(.A(new_n347), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n297), .A2(new_n301), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n287), .B2(new_n288), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n289), .A2(new_n297), .A3(new_n301), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n203), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n523), .A2(new_n310), .B1(new_n308), .B2(KEYINPUT36), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n519), .A2(new_n494), .B1(new_n524), .B2(new_n307), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT35), .B1(new_n519), .B2(new_n509), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n510), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT16), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(G1gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(G1gat), .B2(new_n533), .ZN(new_n536));
  INV_X1    g335(.A(G8gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(G43gat), .A2(G50gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(G43gat), .A2(G50gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT15), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT89), .B(G43gat), .Z(new_n542));
  INV_X1    g341(.A(G50gat), .ZN(new_n543));
  AOI211_X1 g342(.A(KEYINPUT15), .B(new_n539), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(G29gat), .A2(G36gat), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(KEYINPUT14), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(KEYINPUT14), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT88), .B(G29gat), .ZN(new_n548));
  INV_X1    g347(.A(G36gat), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n541), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n550), .A2(new_n541), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT17), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n551), .A2(new_n552), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT90), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n553), .A2(new_n558), .A3(KEYINPUT17), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n538), .B(new_n554), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G229gat), .A2(G233gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n538), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n555), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT18), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n560), .A2(KEYINPUT18), .A3(new_n561), .A4(new_n563), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n553), .B2(new_n538), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n561), .B(KEYINPUT13), .Z(new_n571));
  NAND3_X1  g370(.A1(new_n562), .A2(new_n555), .A3(new_n568), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G197gat), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT11), .B(G169gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT12), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n566), .A2(new_n573), .A3(new_n581), .A4(new_n567), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n202), .B1(new_n532), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n583), .ZN(new_n586));
  AOI211_X1 g385(.A(KEYINPUT92), .B(new_n586), .C1(new_n515), .C2(new_n531), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n517), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n598), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n602), .B(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n608), .B2(new_n605), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n554), .B(new_n609), .C1(new_n557), .C2(new_n559), .ZN(new_n610));
  XOR2_X1   g409(.A(G190gat), .B(G218gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n609), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n613), .A2(new_n555), .B1(KEYINPUT41), .B2(new_n591), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n610), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n612), .B1(new_n610), .B2(new_n614), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n595), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n594), .A3(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(G71gat), .A2(G78gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G57gat), .B(G64gat), .Z(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n626), .B2(KEYINPUT93), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(KEYINPUT9), .B2(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI221_X1 g428(.A(new_n626), .B1(KEYINPUT9), .B2(new_n623), .C1(new_n625), .C2(KEYINPUT93), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(KEYINPUT21), .ZN(new_n632));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n562), .B1(KEYINPUT21), .B2(new_n631), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT95), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT94), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n636), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n631), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n609), .A2(KEYINPUT97), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT97), .B1(new_n609), .B2(new_n651), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n608), .A2(new_n631), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT98), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n608), .A2(new_n657), .A3(new_n631), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n656), .A2(new_n658), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n663), .B(new_n664), .C1(new_n652), .C2(new_n653), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n631), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n650), .B1(new_n661), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n660), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n670), .B(new_n649), .C1(new_n660), .C2(new_n659), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n646), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n589), .A2(new_n590), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g476(.A(new_n674), .B1(new_n585), .B2(new_n588), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n347), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n537), .B1(new_n678), .B2(new_n347), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n679), .B2(new_n681), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(G1325gat));
  XOR2_X1   g486(.A(new_n312), .B(KEYINPUT100), .Z(new_n688));
  NAND3_X1  g487(.A1(new_n678), .A2(G15gat), .A3(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n308), .B(new_n675), .C1(new_n584), .C2(new_n587), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT99), .ZN(new_n691));
  INV_X1    g490(.A(G15gat), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(new_n690), .B2(new_n692), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n689), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n689), .B(new_n697), .C1(new_n693), .C2(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1326gat));
  NAND3_X1  g498(.A1(new_n589), .A2(new_n494), .A3(new_n675), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NOR3_X1   g501(.A1(new_n672), .A2(new_n621), .A3(new_n644), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n589), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n590), .A2(new_n548), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n706), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n508), .A2(new_n514), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n621), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n532), .A2(KEYINPUT44), .A3(new_n622), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n644), .B(KEYINPUT102), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(new_n586), .A3(new_n672), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n517), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n709), .B(new_n710), .C1(new_n548), .C2(new_n719), .ZN(G1328gat));
  NAND4_X1  g519(.A1(new_n589), .A2(new_n549), .A3(new_n347), .A4(new_n703), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n721), .A2(KEYINPUT103), .A3(KEYINPUT46), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n713), .A2(new_n714), .A3(new_n347), .A4(new_n717), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n723), .A2(G36gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n721), .B1(new_n724), .B2(KEYINPUT46), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT103), .B1(new_n721), .B2(KEYINPUT46), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(G1329gat));
  INV_X1    g526(.A(new_n542), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT47), .B(new_n728), .C1(new_n718), .C2(new_n312), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n589), .A2(new_n542), .A3(new_n308), .A4(new_n703), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n713), .A2(new_n714), .A3(new_n688), .A4(new_n717), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n728), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n731), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n733), .A2(new_n738), .ZN(G1330gat));
  NAND4_X1  g538(.A1(new_n589), .A2(new_n543), .A3(new_n494), .A4(new_n703), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n713), .A2(new_n714), .A3(new_n494), .A4(new_n717), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G50gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1331gat));
  NAND3_X1  g544(.A1(new_n646), .A2(new_n586), .A3(new_n672), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n711), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n590), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g548(.A(new_n518), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT105), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1333gat));
  NAND2_X1  g553(.A1(new_n747), .A2(new_n688), .ZN(new_n755));
  INV_X1    g554(.A(new_n308), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(G71gat), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n755), .A2(G71gat), .B1(new_n747), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n747), .A2(new_n494), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT106), .B(G78gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1335gat));
  NOR3_X1   g561(.A1(new_n673), .A2(new_n583), .A3(new_n644), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n715), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n517), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n712), .A2(new_n586), .A3(new_n645), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT51), .Z(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n672), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n590), .A2(new_n599), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n673), .A2(new_n518), .A3(G92gat), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT108), .Z(new_n772));
  AND2_X1   g571(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n713), .A2(new_n714), .A3(new_n347), .A4(new_n763), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(KEYINPUT107), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT52), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n767), .A2(new_n778), .A3(new_n771), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n779), .B(new_n775), .C1(KEYINPUT107), .C2(new_n778), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1337gat));
  INV_X1    g580(.A(new_n688), .ZN(new_n782));
  OAI21_X1  g581(.A(G99gat), .B1(new_n764), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n756), .A2(G99gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n768), .B2(new_n784), .ZN(G1338gat));
  OR3_X1    g584(.A1(new_n460), .A2(new_n673), .A3(G106gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT110), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n767), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n713), .A2(new_n714), .A3(new_n494), .A4(new_n763), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n789), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT53), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n786), .A2(KEYINPUT53), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n767), .A2(new_n792), .B1(KEYINPUT109), .B2(KEYINPUT53), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(G106gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n665), .A2(new_n662), .A3(new_n666), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n670), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n649), .B1(new_n667), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n671), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n798), .B2(new_n800), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n561), .B1(new_n560), .B2(new_n563), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n571), .B1(new_n570), .B2(new_n572), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n578), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n582), .A2(new_n618), .A3(new_n620), .A4(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n802), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n801), .A2(new_n671), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n798), .A2(new_n800), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n811), .A2(new_n812), .B1(new_n580), .B2(new_n582), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n582), .A2(new_n806), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n810), .A2(new_n813), .B1(new_n672), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n809), .B1(new_n815), .B2(new_n622), .ZN(new_n816));
  INV_X1    g615(.A(new_n716), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n674), .A2(new_n583), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n509), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n590), .A2(new_n518), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n583), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n672), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G120gat), .ZN(G1341gat));
  AND3_X1   g628(.A1(new_n825), .A2(G127gat), .A3(new_n716), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n824), .A2(KEYINPUT111), .A3(new_n645), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(G127gat), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT111), .B1(new_n824), .B2(new_n645), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n825), .A2(new_n622), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G134gat), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(G134gat), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n838), .B2(KEYINPUT56), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n837), .A2(KEYINPUT112), .A3(new_n841), .ZN(new_n842));
  OAI221_X1 g641(.A(new_n836), .B1(KEYINPUT56), .B2(new_n838), .C1(new_n840), .C2(new_n842), .ZN(G1343gat));
  NAND2_X1  g642(.A1(new_n380), .A2(new_n381), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n312), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n460), .B1(new_n818), .B2(new_n820), .ZN(new_n847));
  XOR2_X1   g646(.A(KEYINPUT113), .B(KEYINPUT57), .Z(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n819), .B1(new_n816), .B2(new_n645), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n460), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n846), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n844), .B1(new_n854), .B2(new_n586), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n847), .A2(new_n782), .A3(new_n823), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n360), .A3(new_n583), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT114), .B(KEYINPUT58), .Z(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(G1344gat));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n362), .A3(new_n672), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n362), .A2(KEYINPUT59), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n854), .B2(new_n673), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT115), .Z(new_n864));
  XNOR2_X1  g663(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n494), .B1(new_n851), .B2(KEYINPUT118), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n672), .A2(new_n814), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n811), .A2(new_n812), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n583), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n869), .B2(new_n802), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n808), .B1(new_n870), .B2(new_n621), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n820), .B1(new_n871), .B2(new_n644), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n852), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n847), .A2(new_n849), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n673), .B1(new_n845), .B2(KEYINPUT117), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n877), .B(new_n878), .C1(KEYINPUT117), .C2(new_n845), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n865), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n880), .ZN(G1345gat));
  AOI21_X1  g680(.A(G155gat), .B1(new_n856), .B2(new_n644), .ZN(new_n882));
  INV_X1    g681(.A(new_n854), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n716), .A2(G155gat), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT119), .Z(new_n885));
  AOI21_X1  g684(.A(new_n882), .B1(new_n883), .B2(new_n885), .ZN(G1346gat));
  NAND3_X1  g685(.A1(new_n856), .A2(new_n378), .A3(new_n622), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n854), .A2(new_n621), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n378), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n590), .A2(new_n518), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n821), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n586), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(new_n220), .ZN(G1348gat));
  AND2_X1   g692(.A1(new_n821), .A2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n672), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G176gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n247), .B2(new_n895), .ZN(G1349gat));
  AOI21_X1  g696(.A(new_n237), .B1(new_n894), .B2(new_n716), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n891), .A2(new_n261), .A3(new_n645), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT120), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g700(.A1(new_n894), .A2(new_n622), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT121), .B1(new_n902), .B2(G190gat), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(KEYINPUT121), .A3(G190gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(KEYINPUT122), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n908), .B(new_n239), .C1(new_n894), .C2(new_n622), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(KEYINPUT61), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n239), .A3(new_n622), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n911), .B(new_n912), .C1(KEYINPUT61), .C2(new_n910), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n688), .A2(new_n518), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n590), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n460), .B1(new_n872), .B2(new_n873), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n851), .A2(KEYINPUT118), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT57), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n847), .A2(new_n849), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n583), .B(new_n916), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n877), .A2(KEYINPUT124), .A3(new_n583), .A4(new_n916), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n924), .A3(G197gat), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n915), .B2(new_n460), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n914), .A2(KEYINPUT123), .A3(new_n494), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n590), .B1(new_n818), .B2(new_n820), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OR3_X1    g729(.A1(new_n930), .A2(G197gat), .A3(new_n586), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n925), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1352gat));
  NOR3_X1   g735(.A1(new_n930), .A2(G204gat), .A3(new_n673), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT62), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n877), .A2(new_n916), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n672), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G204gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(G1353gat));
  OR3_X1    g741(.A1(new_n930), .A2(G211gat), .A3(new_n645), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n939), .A2(new_n644), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1354gat));
  INV_X1    g746(.A(new_n930), .ZN(new_n948));
  AOI21_X1  g747(.A(G218gat), .B1(new_n948), .B2(new_n622), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n622), .A2(G218gat), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT127), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n952), .B1(new_n939), .B2(KEYINPUT126), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n949), .B1(new_n950), .B2(new_n953), .ZN(G1355gat));
endmodule


