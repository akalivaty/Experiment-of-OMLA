//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT69), .ZN(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  AOI21_X1  g048(.A(new_n465), .B1(new_n462), .B2(new_n463), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n465), .A2(G112), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(G136), .B2(new_n464), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g055(.A(G138), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n465), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n462), .B2(new_n463), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(KEYINPUT71), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n482), .B(KEYINPUT71), .C1(new_n484), .C2(new_n483), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n488), .B(new_n494), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(G543), .B1(KEYINPUT75), .B2(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n503), .A2(KEYINPUT75), .A3(KEYINPUT5), .A4(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT76), .Z(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT77), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n507), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT6), .B1(new_n514), .B2(new_n516), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n514), .B(KEYINPUT6), .C1(new_n515), .C2(new_n516), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n513), .A2(new_n519), .A3(G88), .A4(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n519), .A2(G50), .A3(G543), .A4(new_n520), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n524), .B(G651), .C1(new_n508), .C2(new_n510), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n512), .A2(new_n523), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n519), .A2(new_n520), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n506), .A2(new_n507), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n513), .A2(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n531), .A2(new_n534), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  XOR2_X1   g116(.A(KEYINPUT78), .B(G90), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n530), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n533), .A2(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n516), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR3_X1    g124(.A1(new_n549), .A2(KEYINPUT79), .A3(new_n516), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT79), .B1(new_n549), .B2(new_n516), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n513), .A2(new_n519), .A3(G81), .A4(new_n520), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n519), .A2(G43), .A3(G543), .A4(new_n520), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g133(.A(KEYINPUT80), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n530), .A2(G91), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n513), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT82), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n519), .A2(G543), .A3(new_n520), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n563), .A2(new_n567), .A3(new_n573), .A4(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  NAND2_X1  g151(.A1(new_n530), .A2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n533), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n513), .A2(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n516), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n513), .A2(new_n519), .A3(G86), .A4(new_n520), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n519), .A2(G48), .A3(G543), .A4(new_n520), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n584), .A2(new_n587), .A3(KEYINPUT83), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(KEYINPUT83), .B1(new_n584), .B2(new_n587), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(G305));
  XNOR2_X1  g166(.A(KEYINPUT84), .B(G85), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n530), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n533), .A2(G47), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n593), .B(new_n594), .C1(new_n516), .C2(new_n595), .ZN(G290));
  NAND4_X1  g171(.A1(new_n513), .A2(new_n519), .A3(G92), .A4(new_n520), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G79), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT85), .B1(new_n600), .B2(new_n532), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n600), .A2(new_n532), .A3(KEYINPUT85), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT86), .B(G66), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n529), .C2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n533), .B2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  AND4_X1   g186(.A1(new_n563), .A2(new_n567), .A3(new_n573), .A4(new_n574), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G297));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G280));
  INV_X1    g189(.A(new_n606), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n555), .A2(new_n607), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n606), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n469), .A2(new_n466), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XOR2_X1   g198(.A(KEYINPUT87), .B(KEYINPUT13), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n464), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n474), .A2(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n465), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2096), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n625), .B2(new_n626), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n628), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT90), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT89), .B(KEYINPUT14), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n644), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(G14), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT91), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n656), .A2(new_n657), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n661), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT92), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n670), .A2(new_n671), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(new_n673), .ZN(new_n679));
  MUX2_X1   g254(.A(new_n679), .B(new_n678), .S(new_n669), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  NOR2_X1   g262(.A1(G29), .A2(G35), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G162), .B2(G29), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT29), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(G2090), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n556), .A2(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G16), .B2(G19), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT95), .B(G1341), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G20), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT23), .Z(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G299), .B2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G1956), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n695), .A2(new_n696), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n697), .A2(G21), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G168), .B2(new_n697), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G1966), .ZN(new_n706));
  NOR2_X1   g281(.A1(G171), .A2(new_n697), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G5), .B2(new_n697), .ZN(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n709), .B2(new_n708), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n464), .A2(G139), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n714), .B(new_n715), .C1(new_n465), .C2(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G33), .B(new_n717), .S(G29), .Z(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT24), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G34), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n720), .B2(G34), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G160), .B2(G29), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n718), .A2(G2072), .B1(G2084), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(KEYINPUT31), .A2(G11), .ZN(new_n725));
  NAND2_X1  g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n633), .A2(new_n719), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT30), .B(G28), .ZN(new_n729));
  AOI211_X1 g304(.A(new_n727), .B(new_n728), .C1(new_n719), .C2(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n724), .B(new_n730), .C1(G2072), .C2(new_n718), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n719), .A2(G32), .ZN(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT26), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n474), .A2(G129), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n464), .A2(G141), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n466), .A2(G105), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n732), .B1(new_n740), .B2(new_n719), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT27), .B(G1996), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n743), .B1(G2084), .B2(new_n723), .C1(new_n705), .C2(G1966), .ZN(new_n744));
  NOR2_X1   g319(.A1(G27), .A2(G29), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G164), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2078), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n731), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n711), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n719), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT28), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n464), .A2(G140), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n474), .A2(G128), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n465), .A2(G116), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n751), .B1(new_n760), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  INV_X1    g337(.A(G1348), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n615), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G4), .B2(G16), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n763), .B2(new_n765), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n691), .A2(new_n703), .A3(new_n749), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n464), .A2(G131), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n474), .A2(G119), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n465), .A2(G107), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n769), .B(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  MUX2_X1   g348(.A(G25), .B(new_n773), .S(G29), .Z(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT93), .Z(new_n775));
  XOR2_X1   g350(.A(KEYINPUT35), .B(G1991), .Z(new_n776));
  AOI22_X1  g351(.A1(new_n775), .A2(new_n776), .B1(KEYINPUT94), .B2(KEYINPUT36), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  MUX2_X1   g353(.A(G24), .B(G290), .S(G16), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1986), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G166), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G16), .B2(G22), .ZN(new_n783));
  INV_X1    g358(.A(G1971), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n697), .A2(G23), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G288), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n785), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(G6), .A2(G16), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G305), .B2(new_n697), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT32), .B(G1981), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n791), .A2(KEYINPUT34), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(KEYINPUT34), .B1(new_n791), .B2(new_n795), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n781), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(KEYINPUT94), .B2(KEYINPUT36), .ZN(new_n799));
  NOR2_X1   g374(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(new_n781), .C1(new_n796), .C2(new_n797), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n768), .B1(new_n799), .B2(new_n801), .ZN(G311));
  XNOR2_X1  g377(.A(G311), .B(KEYINPUT98), .ZN(G150));
  NAND2_X1  g378(.A1(G80), .A2(G543), .ZN(new_n804));
  INV_X1    g379(.A(G67), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n529), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(KEYINPUT99), .B(new_n804), .C1(new_n529), .C2(new_n805), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n808), .A2(G651), .A3(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(G93), .A2(new_n530), .B1(new_n533), .B2(G55), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n615), .A2(G559), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT38), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n555), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n551), .A2(new_n554), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n818), .A2(new_n810), .A3(new_n550), .A4(new_n811), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n816), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT100), .Z(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n822), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n814), .B1(new_n824), .B2(new_n826), .ZN(G145));
  XOR2_X1   g402(.A(G160), .B(new_n633), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G162), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n760), .B(G164), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(new_n717), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n717), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n740), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n623), .B(new_n773), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n474), .A2(G130), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT101), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n464), .A2(G142), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n465), .A2(G118), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n836), .B(new_n842), .Z(new_n843));
  NAND3_X1  g418(.A1(new_n831), .A2(new_n740), .A3(new_n832), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n835), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n843), .B1(new_n835), .B2(new_n844), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n846), .A3(new_n845), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n829), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n849), .A2(new_n829), .A3(new_n845), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(G395));
  NAND2_X1  g433(.A1(new_n812), .A2(new_n607), .ZN(new_n859));
  NAND2_X1  g434(.A1(G290), .A2(G288), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(G290), .A2(G288), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT106), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(G290), .A2(G288), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT106), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT105), .B1(new_n589), .B2(new_n590), .ZN(new_n868));
  INV_X1    g443(.A(new_n590), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n870), .A3(new_n588), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G166), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n871), .A3(G303), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n867), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n866), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n873), .B2(new_n874), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT42), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n612), .A2(new_n606), .ZN(new_n881));
  NAND3_X1  g456(.A1(G299), .A2(new_n599), .A3(new_n605), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g460(.A(KEYINPUT104), .B(KEYINPUT41), .C1(new_n881), .C2(new_n882), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n820), .B(new_n619), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(KEYINPUT103), .A3(new_n882), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n615), .A2(new_n890), .A3(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n892), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n879), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n859), .B1(new_n897), .B2(new_n607), .ZN(G295));
  OAI21_X1  g473(.A(new_n859), .B1(new_n897), .B2(new_n607), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n817), .A2(new_n819), .A3(G301), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G301), .B1(new_n817), .B2(new_n819), .ZN(new_n903));
  OAI21_X1  g478(.A(G286), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n820), .A2(G171), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(G168), .A3(new_n901), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n887), .A2(new_n904), .A3(new_n893), .A4(new_n906), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n902), .A2(new_n903), .A3(G286), .ZN(new_n908));
  AOI21_X1  g483(.A(G168), .B1(new_n905), .B2(new_n901), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n892), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n875), .A2(new_n877), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n892), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT41), .A4(new_n883), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n878), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n854), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT107), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n911), .B2(new_n912), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(new_n917), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n900), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n878), .A2(new_n910), .A3(new_n907), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT43), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n900), .B1(new_n920), .B2(new_n924), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(G397));
  XNOR2_X1  g506(.A(KEYINPUT108), .B(G1384), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT45), .B1(new_n500), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G40), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n468), .A2(new_n472), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1996), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(new_n834), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT110), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n760), .A2(G2067), .ZN(new_n941));
  INV_X1    g516(.A(G2067), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n758), .A2(new_n942), .A3(new_n759), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n740), .A2(new_n937), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n936), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n776), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n773), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n773), .A2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n936), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NOR2_X1   g528(.A1(G290), .A2(G1986), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n936), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT109), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G8), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n489), .A2(new_n493), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT71), .B1(new_n469), .B2(new_n482), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n487), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n485), .A2(new_n486), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n964), .B2(new_n935), .ZN(new_n965));
  INV_X1    g540(.A(G1981), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n584), .A2(new_n587), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n585), .A2(new_n586), .ZN(new_n968));
  OAI21_X1  g543(.A(G1981), .B1(new_n583), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n967), .A2(KEYINPUT49), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT49), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n964), .A2(new_n935), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G8), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n974), .A2(G1976), .A3(G288), .ZN(new_n975));
  INV_X1    g550(.A(new_n967), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n965), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n962), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n488), .A2(new_n493), .A3(new_n489), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT45), .B(new_n932), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(new_n935), .C1(new_n964), .C2(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n784), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n964), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n470), .A2(new_n471), .ZN(new_n986));
  OAI211_X1 g561(.A(G40), .B(new_n467), .C1(new_n986), .C2(new_n465), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n964), .B2(new_n984), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n978), .B2(new_n979), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n982), .B1(new_n992), .B2(G2090), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g569(.A1(G303), .A2(G8), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  NAND4_X1  g573(.A1(G303), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(G8), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n993), .A2(new_n1000), .A3(G8), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT113), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n993), .A2(new_n1000), .A3(new_n1003), .A4(G8), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n577), .A2(new_n578), .A3(G1976), .A4(new_n579), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n965), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(new_n965), .A3(new_n1006), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(new_n974), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n977), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n500), .A2(new_n984), .A3(new_n989), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n984), .B1(new_n500), .B2(new_n989), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n935), .B(new_n1016), .C1(new_n1017), .C2(KEYINPUT111), .ZN(new_n1018));
  INV_X1    g593(.A(new_n991), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT120), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT120), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n985), .A2(new_n988), .A3(new_n1021), .A4(new_n991), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n709), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n987), .B1(new_n990), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G2078), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT124), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1025), .A2(KEYINPUT124), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(KEYINPUT53), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n981), .B2(G2078), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1023), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1035), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT125), .B1(new_n1035), .B2(G171), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1000), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n1017), .B2(new_n987), .ZN(new_n1041));
  OAI211_X1 g616(.A(KEYINPUT114), .B(new_n935), .C1(new_n964), .C2(new_n984), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1016), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  AOI21_X1  g619(.A(G2090), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1041), .A2(KEYINPUT115), .A3(new_n1042), .A4(new_n1016), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1045), .A2(new_n1046), .B1(new_n784), .B2(new_n981), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1039), .B1(new_n1047), .B2(new_n958), .ZN(new_n1048));
  OR3_X1    g623(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT116), .B1(new_n1012), .B2(new_n974), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(new_n1005), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1038), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n985), .A2(new_n988), .A3(new_n1056), .A4(new_n991), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n935), .B1(new_n964), .B2(KEYINPUT45), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n990), .A2(new_n1024), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1061), .A3(G168), .ZN(new_n1062));
  AND2_X1   g637(.A1(KEYINPUT123), .A2(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(KEYINPUT51), .A3(new_n1063), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(G8), .A3(G286), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n958), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(KEYINPUT122), .A3(G286), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1068), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1015), .B1(new_n1055), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n612), .B(KEYINPUT57), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1025), .A2(new_n980), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1043), .A2(new_n1084), .A3(new_n701), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1043), .B2(new_n701), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1081), .B(new_n1083), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1020), .A2(new_n763), .A3(new_n1022), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n964), .A2(new_n935), .A3(new_n942), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n615), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1081), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1088), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n606), .A4(new_n1090), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n990), .A2(new_n1024), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1099), .A2(new_n937), .A3(new_n935), .A4(new_n980), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n972), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n555), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1098), .B1(new_n1103), .B2(KEYINPUT121), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n981), .B2(G1996), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n556), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1107), .A3(new_n1098), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1097), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1091), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n615), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT61), .B1(new_n1095), .B2(new_n1087), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1087), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1096), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1002), .A2(new_n1004), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1074), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT122), .B1(new_n1073), .B2(G286), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1062), .A2(KEYINPUT51), .A3(new_n1063), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT51), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1122), .A2(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1121), .A2(new_n1126), .A3(new_n1048), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1033), .B1(KEYINPUT126), .B2(new_n1026), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(KEYINPUT126), .B2(new_n1026), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n933), .A2(new_n987), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n980), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1023), .A2(new_n1034), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G171), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(KEYINPUT54), .C1(G171), .C2(new_n1035), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1132), .A2(G171), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1036), .A2(new_n1037), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1127), .B(new_n1134), .C1(new_n1136), .C2(KEYINPUT54), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1080), .B1(new_n1120), .B2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1073), .A2(G168), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1121), .A2(new_n1048), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1005), .A2(KEYINPUT63), .A3(new_n1139), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n993), .A2(G8), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1013), .B1(new_n1146), .B2(new_n1000), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1147), .A2(KEYINPUT118), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(KEYINPUT118), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1143), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n957), .B1(new_n1138), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n936), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n947), .A2(new_n949), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n943), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT46), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n938), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT127), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n938), .A2(new_n1156), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n936), .B1(new_n944), .B2(new_n834), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT47), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n954), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT48), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n1155), .B(new_n1162), .C1(new_n952), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g741(.A1(new_n928), .A2(new_n929), .ZN(new_n1168));
  OR3_X1    g742(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1169));
  OR2_X1    g743(.A1(G229), .A2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g744(.A1(new_n856), .A2(new_n1168), .A3(new_n1170), .ZN(G308));
  OR3_X1    g745(.A1(new_n856), .A2(new_n1168), .A3(new_n1170), .ZN(G225));
endmodule


