

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  NAND2_X1 U321 ( .A1(n407), .A2(n406), .ZN(n486) );
  XNOR2_X1 U322 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U323 ( .A(KEYINPUT41), .B(n570), .Z(n559) );
  XNOR2_X1 U324 ( .A(KEYINPUT38), .B(n453), .ZN(n502) );
  XOR2_X1 U325 ( .A(KEYINPUT28), .B(n472), .Z(n534) );
  XOR2_X1 U326 ( .A(n392), .B(n371), .Z(n520) );
  XOR2_X1 U327 ( .A(n471), .B(KEYINPUT54), .Z(n289) );
  AND2_X1 U328 ( .A1(n556), .A2(n559), .ZN(n462) );
  NOR2_X1 U329 ( .A1(n459), .A2(n570), .ZN(n460) );
  XOR2_X1 U330 ( .A(G36GAT), .B(KEYINPUT78), .Z(n366) );
  XNOR2_X1 U331 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U332 ( .A(n367), .B(G8GAT), .ZN(n368) );
  XNOR2_X1 U333 ( .A(n426), .B(n425), .ZN(n431) );
  XNOR2_X1 U334 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U335 ( .A(n380), .B(n368), .ZN(n369) );
  XNOR2_X1 U336 ( .A(n321), .B(n320), .ZN(n329) );
  XOR2_X1 U337 ( .A(n393), .B(n392), .Z(n522) );
  INV_X1 U338 ( .A(G29GAT), .ZN(n454) );
  XNOR2_X1 U339 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U340 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U341 ( .A(n481), .B(n480), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n457), .B(n456), .ZN(G1328GAT) );
  XNOR2_X1 U343 ( .A(G127GAT), .B(G134GAT), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n290), .B(KEYINPUT84), .ZN(n291) );
  XOR2_X1 U345 ( .A(n291), .B(KEYINPUT0), .Z(n293) );
  XNOR2_X1 U346 ( .A(G113GAT), .B(G120GAT), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n391) );
  XOR2_X1 U348 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n295) );
  XNOR2_X1 U349 ( .A(KEYINPUT6), .B(KEYINPUT92), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U351 ( .A(KEYINPUT93), .B(KEYINPUT95), .Z(n297) );
  XNOR2_X1 U352 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U354 ( .A(n299), .B(n298), .Z(n308) );
  XOR2_X1 U355 ( .A(KEYINPUT3), .B(G162GAT), .Z(n301) );
  XNOR2_X1 U356 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(G141GAT), .B(n302), .Z(n384) );
  XOR2_X1 U359 ( .A(G29GAT), .B(G1GAT), .Z(n438) );
  XNOR2_X1 U360 ( .A(G148GAT), .B(G85GAT), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n303), .B(G57GAT), .ZN(n416) );
  XOR2_X1 U362 ( .A(n438), .B(n416), .Z(n305) );
  NAND2_X1 U363 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U364 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U365 ( .A(n384), .B(n306), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U367 ( .A(n391), .B(n309), .Z(n403) );
  XOR2_X1 U368 ( .A(KEYINPUT96), .B(n403), .Z(n517) );
  XOR2_X1 U369 ( .A(KEYINPUT73), .B(KEYINPUT77), .Z(n311) );
  XNOR2_X1 U370 ( .A(G106GAT), .B(G85GAT), .ZN(n310) );
  XOR2_X1 U371 ( .A(n311), .B(n310), .Z(n315) );
  XOR2_X1 U372 ( .A(n366), .B(G218GAT), .Z(n313) );
  XOR2_X1 U373 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n447) );
  XNOR2_X1 U374 ( .A(n447), .B(G134GAT), .ZN(n312) );
  XNOR2_X1 U375 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n321) );
  XOR2_X1 U377 ( .A(KEYINPUT64), .B(KEYINPUT65), .Z(n317) );
  XNOR2_X1 U378 ( .A(G29GAT), .B(G162GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n319) );
  AND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XOR2_X1 U381 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n323) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(G50GAT), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U384 ( .A(G92GAT), .B(KEYINPUT9), .Z(n325) );
  XNOR2_X1 U385 ( .A(G190GAT), .B(G99GAT), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n553) );
  XOR2_X1 U389 ( .A(n553), .B(KEYINPUT36), .Z(n578) );
  XOR2_X1 U390 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n331) );
  XNOR2_X1 U391 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n339) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XOR2_X1 U394 ( .A(G155GAT), .B(G183GAT), .Z(n333) );
  XNOR2_X1 U395 ( .A(G15GAT), .B(G22GAT), .ZN(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n335) );
  XOR2_X1 U397 ( .A(G127GAT), .B(G71GAT), .Z(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n351) );
  XOR2_X1 U401 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n341) );
  XNOR2_X1 U402 ( .A(G8GAT), .B(G64GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U404 ( .A(G57GAT), .B(G78GAT), .Z(n343) );
  XNOR2_X1 U405 ( .A(G1GAT), .B(G211GAT), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n349) );
  XNOR2_X1 U408 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n347) );
  XOR2_X1 U409 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n346) );
  XOR2_X1 U410 ( .A(KEYINPUT70), .B(n346), .Z(n427) );
  XOR2_X1 U411 ( .A(n347), .B(n427), .Z(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U413 ( .A(n351), .B(n350), .Z(n575) );
  INV_X1 U414 ( .A(n575), .ZN(n484) );
  XOR2_X1 U415 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n353) );
  XNOR2_X1 U416 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U418 ( .A(n354), .B(KEYINPUT88), .Z(n356) );
  XNOR2_X1 U419 ( .A(G190GAT), .B(G183GAT), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n356), .B(n355), .ZN(n358) );
  XOR2_X1 U421 ( .A(G169GAT), .B(G176GAT), .Z(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n392) );
  XNOR2_X1 U423 ( .A(G204GAT), .B(G92GAT), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n359), .B(G64GAT), .ZN(n428) );
  XOR2_X1 U425 ( .A(n428), .B(KEYINPUT98), .Z(n361) );
  NAND2_X1 U426 ( .A1(G226GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n370) );
  XNOR2_X1 U428 ( .A(G211GAT), .B(KEYINPUT91), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n362), .B(KEYINPUT90), .ZN(n363) );
  XOR2_X1 U430 ( .A(n363), .B(KEYINPUT21), .Z(n365) );
  XNOR2_X1 U431 ( .A(G197GAT), .B(G218GAT), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n380) );
  XOR2_X1 U433 ( .A(KEYINPUT97), .B(n366), .Z(n367) );
  XOR2_X1 U434 ( .A(n370), .B(n369), .Z(n371) );
  XOR2_X1 U435 ( .A(n520), .B(KEYINPUT99), .Z(n372) );
  XNOR2_X1 U436 ( .A(n372), .B(KEYINPUT27), .ZN(n398) );
  NAND2_X1 U437 ( .A1(n398), .A2(n517), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n373), .B(KEYINPUT100), .ZN(n528) );
  XOR2_X1 U439 ( .A(G106GAT), .B(G78GAT), .Z(n411) );
  XOR2_X1 U440 ( .A(n411), .B(G204GAT), .Z(n375) );
  NAND2_X1 U441 ( .A1(G228GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U443 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n377) );
  XNOR2_X1 U444 ( .A(G148GAT), .B(KEYINPUT22), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U446 ( .A(n379), .B(n378), .Z(n382) );
  XOR2_X1 U447 ( .A(G50GAT), .B(G22GAT), .Z(n439) );
  XNOR2_X1 U448 ( .A(n439), .B(n380), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n472) );
  NOR2_X1 U451 ( .A1(n528), .A2(n534), .ZN(n395) );
  XOR2_X1 U452 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n386) );
  NAND2_X1 U453 ( .A1(G227GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U455 ( .A(n387), .B(KEYINPUT86), .Z(n389) );
  XOR2_X1 U456 ( .A(G43GAT), .B(G15GAT), .Z(n442) );
  XOR2_X1 U457 ( .A(G99GAT), .B(G71GAT), .Z(n412) );
  XNOR2_X1 U458 ( .A(n442), .B(n412), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n391), .B(n390), .ZN(n393) );
  INV_X1 U461 ( .A(n522), .ZN(n531) );
  XOR2_X1 U462 ( .A(n531), .B(KEYINPUT89), .Z(n394) );
  NAND2_X1 U463 ( .A1(n395), .A2(n394), .ZN(n407) );
  NOR2_X1 U464 ( .A1(n522), .A2(n472), .ZN(n397) );
  XOR2_X1 U465 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n396) );
  XOR2_X1 U466 ( .A(n397), .B(n396), .Z(n547) );
  INV_X1 U467 ( .A(n547), .ZN(n564) );
  NAND2_X1 U468 ( .A1(n564), .A2(n398), .ZN(n402) );
  NAND2_X1 U469 ( .A1(n522), .A2(n520), .ZN(n399) );
  NAND2_X1 U470 ( .A1(n472), .A2(n399), .ZN(n400) );
  XOR2_X1 U471 ( .A(KEYINPUT25), .B(n400), .Z(n401) );
  NAND2_X1 U472 ( .A1(n402), .A2(n401), .ZN(n404) );
  NAND2_X1 U473 ( .A1(n404), .A2(n403), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n405), .B(KEYINPUT102), .ZN(n406) );
  NAND2_X1 U475 ( .A1(n484), .A2(n486), .ZN(n408) );
  NOR2_X1 U476 ( .A1(n578), .A2(n408), .ZN(n410) );
  XNOR2_X1 U477 ( .A(KEYINPUT106), .B(KEYINPUT37), .ZN(n409) );
  XNOR2_X1 U478 ( .A(n410), .B(n409), .ZN(n516) );
  XOR2_X1 U479 ( .A(KEYINPUT72), .B(n411), .Z(n414) );
  XNOR2_X1 U480 ( .A(G176GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n420) );
  INV_X1 U482 ( .A(KEYINPUT32), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n418) );
  NAND2_X1 U484 ( .A1(G230GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U486 ( .A(n420), .B(n419), .Z(n426) );
  XOR2_X1 U487 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n422) );
  XNOR2_X1 U488 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n421) );
  XOR2_X1 U489 ( .A(n422), .B(n421), .Z(n424) );
  XNOR2_X1 U490 ( .A(G120GAT), .B(KEYINPUT73), .ZN(n423) );
  INV_X1 U491 ( .A(n427), .ZN(n429) );
  XOR2_X1 U492 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n570) );
  XOR2_X1 U494 ( .A(G8GAT), .B(G197GAT), .Z(n433) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G141GAT), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U497 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n435) );
  XNOR2_X1 U498 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n451) );
  XOR2_X1 U501 ( .A(G113GAT), .B(G36GAT), .Z(n441) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U504 ( .A(n443), .B(n442), .Z(n449) );
  XOR2_X1 U505 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n445) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U510 ( .A(n451), .B(n450), .Z(n566) );
  NOR2_X1 U511 ( .A1(n570), .A2(n566), .ZN(n452) );
  XOR2_X1 U512 ( .A(KEYINPUT76), .B(n452), .Z(n488) );
  NOR2_X1 U513 ( .A1(n516), .A2(n488), .ZN(n453) );
  NAND2_X1 U514 ( .A1(n517), .A2(n502), .ZN(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n455) );
  INV_X1 U516 ( .A(n566), .ZN(n556) );
  NOR2_X1 U517 ( .A1(n484), .A2(n578), .ZN(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT45), .B(n458), .Z(n459) );
  XOR2_X1 U519 ( .A(KEYINPUT114), .B(n460), .Z(n461) );
  NOR2_X1 U520 ( .A1(n556), .A2(n461), .ZN(n468) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT46), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n553), .A2(n463), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n484), .ZN(n466) );
  XOR2_X1 U524 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n465) );
  XNOR2_X1 U525 ( .A(n466), .B(n465), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT48), .ZN(n529) );
  XOR2_X1 U528 ( .A(n520), .B(KEYINPUT120), .Z(n470) );
  NOR2_X1 U529 ( .A1(n529), .A2(n470), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n517), .A2(n289), .ZN(n565) );
  NAND2_X1 U531 ( .A1(n565), .A2(n472), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n474) );
  INV_X1 U533 ( .A(KEYINPUT55), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n531), .A2(n477), .ZN(n560) );
  NAND2_X1 U536 ( .A1(n560), .A2(n553), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n479) );
  XNOR2_X1 U538 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n478) );
  NAND2_X1 U539 ( .A1(n575), .A2(n560), .ZN(n483) );
  XNOR2_X1 U540 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(G1350GAT) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n490) );
  NOR2_X1 U543 ( .A1(n553), .A2(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(KEYINPUT16), .ZN(n487) );
  NAND2_X1 U545 ( .A1(n487), .A2(n486), .ZN(n504) );
  NOR2_X1 U546 ( .A1(n488), .A2(n504), .ZN(n495) );
  NAND2_X1 U547 ( .A1(n517), .A2(n495), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n520), .A2(n495), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n493) );
  NAND2_X1 U552 ( .A1(n495), .A2(n522), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U554 ( .A(G15GAT), .B(n494), .Z(G1326GAT) );
  NAND2_X1 U555 ( .A1(n534), .A2(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(KEYINPUT104), .ZN(n497) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n497), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G36GAT), .B(KEYINPUT107), .Z(n499) );
  NAND2_X1 U559 ( .A1(n502), .A2(n520), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n502), .A2(n522), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT40), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n502), .A2(n534), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n507) );
  NAND2_X1 U567 ( .A1(n559), .A2(n566), .ZN(n515) );
  NOR2_X1 U568 ( .A1(n504), .A2(n515), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT108), .ZN(n511) );
  NAND2_X1 U570 ( .A1(n517), .A2(n511), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n511), .A2(n520), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n511), .A2(n522), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U578 ( .A1(n511), .A2(n534), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT111), .Z(n519) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n524) );
  NAND2_X1 U583 ( .A1(n524), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n524), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n524), .A2(n522), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n526) );
  NAND2_X1 U590 ( .A1(n524), .A2(n534), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n527), .Z(G1339GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT115), .ZN(n546) );
  NOR2_X1 U595 ( .A1(n531), .A2(n546), .ZN(n532) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(n532), .Z(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n542), .A2(n556), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n537) );
  NAND2_X1 U601 ( .A1(n542), .A2(n559), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n540) );
  NAND2_X1 U605 ( .A1(n542), .A2(n575), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n553), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n556), .A2(n554), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U616 ( .A1(n554), .A2(n559), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n575), .A2(n554), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT123), .Z(n558) );
  NAND2_X1 U624 ( .A1(n560), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n577) );
  NOR2_X1 U631 ( .A1(n566), .A2(n577), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n572) );
  INV_X1 U636 ( .A(n577), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

