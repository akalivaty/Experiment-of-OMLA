//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n223), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n212), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n245), .A2(KEYINPUT68), .A3(new_n212), .ZN(new_n249));
  AND2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G68), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n252), .A2(G77), .B1(G20), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(new_n201), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g0058(.A(new_n258), .B(KEYINPUT11), .Z(new_n259));
  OR2_X1    g0059(.A1(new_n259), .A2(KEYINPUT75), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(KEYINPUT75), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n262), .A2(new_n213), .A3(G1), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n250), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n253), .B1(new_n265), .B2(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n263), .ZN(new_n267));
  OR3_X1    g0067(.A1(new_n267), .A2(KEYINPUT12), .A3(G68), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT12), .B1(new_n267), .B2(G68), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n264), .A2(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n260), .A2(new_n261), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT14), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G238), .ZN(new_n277));
  AND2_X1   g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  OAI21_X1  g0078(.A(G274), .B1(new_n278), .B2(new_n212), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n276), .A2(new_n277), .B1(new_n279), .B2(new_n275), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT65), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT65), .ZN(new_n288));
  INV_X1    g0088(.A(G226), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n285), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT73), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n285), .A2(KEYINPUT73), .A3(new_n288), .A4(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n285), .A2(G232), .A3(G1698), .A4(new_n288), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G97), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT74), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n274), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(new_n298), .A3(KEYINPUT74), .ZN(new_n302));
  AOI211_X1 g0102(.A(KEYINPUT13), .B(new_n280), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT13), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n300), .ZN(new_n305));
  INV_X1    g0105(.A(new_n274), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n280), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n272), .B(G169), .C1(new_n303), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n296), .A2(new_n297), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n293), .B2(new_n294), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n306), .B1(new_n312), .B2(KEYINPUT74), .ZN(new_n313));
  INV_X1    g0113(.A(new_n302), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n307), .A2(new_n304), .A3(new_n308), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n272), .B1(new_n320), .B2(G169), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n271), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT67), .B(G223), .Z(new_n323));
  INV_X1    g0123(.A(KEYINPUT66), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n285), .A2(new_n288), .ZN(new_n325));
  INV_X1    g0125(.A(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT65), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT65), .B1(new_n286), .B2(new_n287), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(KEYINPUT66), .A3(G1698), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n323), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(G222), .A3(new_n326), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n217), .B2(new_n330), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n306), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n279), .A2(new_n275), .ZN(new_n336));
  INV_X1    g0136(.A(new_n276), .ZN(new_n337));
  XOR2_X1   g0137(.A(KEYINPUT64), .B(G226), .Z(new_n338));
  AOI21_X1  g0138(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n265), .A2(G20), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G50), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n264), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n347));
  INV_X1    g0147(.A(G150), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT8), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n202), .B2(KEYINPUT69), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT69), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(KEYINPUT8), .A3(G58), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n252), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n347), .B1(new_n348), .B2(new_n256), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n250), .B1(new_n201), .B2(new_n263), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n346), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n342), .B(new_n357), .C1(G179), .C2(new_n340), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n346), .A2(new_n356), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT9), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n361), .ZN(new_n363));
  NAND2_X1  g0163(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n340), .A2(G200), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT10), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n335), .A2(G190), .A3(new_n339), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n358), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT71), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n277), .B1(new_n327), .B2(new_n331), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n330), .A2(G232), .A3(new_n326), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n219), .B2(new_n330), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n306), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n336), .B1(G244), .B2(new_n337), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n372), .B1(new_n378), .B2(G179), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n376), .A2(KEYINPUT71), .A3(new_n380), .A4(new_n377), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n341), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT8), .B(G58), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n256), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n250), .B1(new_n217), .B2(new_n263), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n264), .A2(G77), .A3(new_n343), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n379), .A2(new_n381), .A3(new_n382), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n378), .B2(G200), .ZN(new_n392));
  INV_X1    g0192(.A(G190), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n378), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n371), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G200), .B1(new_n303), .B2(new_n309), .ZN(new_n397));
  INV_X1    g0197(.A(new_n271), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n316), .A2(new_n317), .A3(G190), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n248), .A2(new_n249), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n202), .A2(new_n253), .ZN(new_n402));
  NOR2_X1   g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  OAI21_X1  g0203(.A(G20), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n255), .A2(G159), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT76), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT76), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n282), .A3(G33), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n409), .A3(new_n286), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n213), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n253), .B1(new_n411), .B2(KEYINPUT7), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT7), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n413), .A3(new_n213), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n406), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n401), .B1(new_n415), .B2(KEYINPUT16), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n413), .B(new_n213), .C1(new_n328), .C2(new_n329), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n213), .B1(new_n283), .B2(new_n284), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT7), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(G68), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n406), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT16), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n353), .B1(new_n265), .B2(G20), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n264), .A2(new_n425), .B1(new_n263), .B2(new_n353), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT77), .B1(new_n276), .B2(new_n223), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n274), .A2(new_n275), .A3(new_n428), .A4(G232), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n336), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n289), .A2(G1698), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G223), .B2(G1698), .ZN(new_n432));
  INV_X1    g0232(.A(G87), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n410), .A2(new_n432), .B1(new_n251), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n306), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n393), .ZN(new_n437));
  INV_X1    g0237(.A(G200), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n430), .B2(new_n435), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n424), .A2(new_n426), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n412), .A2(new_n414), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT16), .A3(new_n421), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n250), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n426), .B1(new_n446), .B2(new_n422), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(G169), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n380), .B2(new_n436), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT18), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(KEYINPUT18), .A3(new_n449), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(KEYINPUT78), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT78), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n447), .A2(new_n453), .A3(KEYINPUT18), .A4(new_n449), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n443), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  AND4_X1   g0255(.A1(new_n322), .A2(new_n396), .A3(new_n400), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n285), .A2(G250), .A3(G1698), .A4(new_n288), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT4), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n218), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n285), .A2(new_n326), .A3(new_n288), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n218), .A2(G1698), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n407), .A2(new_n409), .A3(new_n286), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n459), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n458), .A2(new_n461), .A3(new_n462), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n306), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n468), .A2(new_n274), .A3(G274), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n274), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n471), .B1(new_n475), .B2(new_n225), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n476), .B1(new_n466), .B2(new_n306), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(G190), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n438), .B1(new_n467), .B2(new_n477), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n224), .A2(KEYINPUT79), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT79), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G97), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(new_n219), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT79), .B(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n219), .A2(KEYINPUT6), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n224), .A2(new_n219), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n489), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n417), .A2(G107), .A3(new_n419), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n401), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n267), .A2(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n265), .A2(G33), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n401), .A2(new_n267), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(G97), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n484), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n481), .B1(new_n467), .B2(new_n477), .ZN(new_n509));
  AOI211_X1 g0309(.A(KEYINPUT81), .B(new_n476), .C1(new_n466), .C2(new_n306), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n341), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n498), .A2(G20), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n255), .A2(G77), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n500), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n250), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(new_n506), .B1(new_n380), .B2(new_n480), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n483), .A2(new_n508), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n218), .A2(G1698), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(G238), .B2(G1698), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n410), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT82), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(KEYINPUT82), .B(new_n518), .C1(new_n410), .C2(new_n520), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(new_n306), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n470), .A2(G250), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n306), .ZN(new_n527));
  INV_X1    g0327(.A(G274), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n470), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n393), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n438), .B1(new_n525), .B2(new_n530), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n491), .A2(new_n433), .A3(new_n219), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n213), .B1(new_n297), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n488), .A2(new_n252), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n407), .A2(new_n409), .A3(new_n213), .A4(new_n286), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n253), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n250), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n505), .A2(G87), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n383), .A2(new_n263), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n532), .A2(new_n533), .A3(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n536), .A2(new_n534), .B1(new_n538), .B2(new_n535), .ZN(new_n548));
  INV_X1    g0348(.A(new_n542), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n401), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n504), .A2(new_n383), .ZN(new_n551));
  INV_X1    g0351(.A(new_n545), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n525), .A2(G179), .A3(new_n530), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n274), .B1(new_n521), .B2(new_n522), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n524), .B1(new_n529), .B2(new_n527), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n341), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n553), .B1(new_n557), .B2(KEYINPUT83), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT83), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n554), .B(new_n559), .C1(new_n341), .C2(new_n556), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n547), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT23), .B1(new_n213), .B2(G107), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT85), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT85), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n564), .B(KEYINPUT23), .C1(new_n213), .C2(G107), .ZN(new_n565));
  OR3_X1    g0365(.A1(new_n213), .A2(KEYINPUT23), .A3(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n213), .A2(G33), .A3(G116), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n563), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT22), .B1(new_n541), .B2(new_n433), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n433), .A2(KEYINPUT22), .A3(G20), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n285), .A2(new_n288), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI211_X1 g0374(.A(KEYINPUT24), .B(new_n568), .C1(new_n569), .C2(new_n571), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n250), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n225), .A2(G1698), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G250), .B2(G1698), .ZN(new_n578));
  INV_X1    g0378(.A(G294), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n410), .A2(new_n578), .B1(new_n251), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n212), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n468), .A2(new_n470), .B1(new_n581), .B2(new_n273), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n580), .A2(new_n306), .B1(G264), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n393), .A3(new_n471), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n474), .A2(new_n279), .ZN(new_n585));
  AOI221_X4 g0385(.A(new_n585), .B1(new_n582), .B2(G264), .C1(new_n580), .C2(new_n306), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n586), .B2(G200), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n263), .A2(new_n219), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT25), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n505), .B2(G107), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n576), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT86), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT86), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n576), .A2(new_n587), .A3(new_n593), .A4(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT84), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n401), .A2(G116), .A3(new_n267), .A4(new_n503), .ZN(new_n598));
  INV_X1    g0398(.A(G116), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n263), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n245), .A2(new_n212), .B1(G20), .B2(new_n599), .ZN(new_n601));
  AOI21_X1  g0401(.A(G33), .B1(new_n485), .B2(new_n487), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n462), .A2(new_n213), .ZN(new_n603));
  OAI211_X1 g0403(.A(KEYINPUT20), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n603), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n491), .B2(G33), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT20), .B1(new_n607), .B2(new_n601), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n598), .B(new_n600), .C1(new_n605), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(G303), .B1(new_n328), .B2(new_n329), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n407), .A2(new_n409), .A3(new_n286), .ZN(new_n612));
  NOR2_X1   g0412(.A1(G257), .A2(G1698), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n220), .B2(G1698), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n274), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G270), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n471), .B1(new_n475), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(G169), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n597), .B1(new_n610), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(G303), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n285), .B2(new_n288), .ZN(new_n622));
  INV_X1    g0422(.A(new_n614), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(new_n410), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n306), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n618), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G190), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(G200), .B1(new_n616), .B2(new_n618), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n610), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(new_n626), .ZN(new_n630));
  INV_X1    g0430(.A(new_n597), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n630), .A2(new_n609), .A3(G169), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n616), .A2(new_n618), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n609), .A3(G179), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n620), .A2(new_n629), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n583), .A2(new_n380), .A3(new_n471), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n586), .B2(G169), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n576), .B2(new_n590), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n517), .A2(new_n561), .A3(new_n595), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n457), .A2(new_n640), .ZN(G372));
  NAND2_X1  g0441(.A1(new_n447), .A2(new_n449), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT18), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n451), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n322), .A2(new_n391), .ZN(new_n647));
  INV_X1    g0447(.A(new_n400), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n443), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n646), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n369), .A2(new_n370), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n358), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(KEYINPUT89), .B(new_n358), .C1(new_n650), .C2(new_n651), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n553), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n557), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n550), .A2(new_n552), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n659), .B(new_n544), .C1(new_n438), .C2(new_n556), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT87), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n532), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OR3_X1    g0462(.A1(new_n546), .A2(new_n533), .A3(new_n661), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n638), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n620), .A2(new_n634), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n632), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n664), .A2(new_n667), .A3(new_n595), .A4(new_n517), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n558), .A2(new_n560), .ZN(new_n669));
  INV_X1    g0469(.A(new_n547), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n511), .A2(new_n516), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT26), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT88), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n511), .A2(KEYINPUT88), .A3(new_n516), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n664), .A2(new_n675), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n658), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n668), .A2(new_n673), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n456), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n656), .A2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n666), .A2(new_n632), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n265), .A2(new_n213), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n610), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n635), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n638), .A2(new_n690), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n690), .B1(new_n576), .B2(new_n590), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n592), .B2(new_n594), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n695), .B1(new_n697), .B2(new_n638), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n683), .A2(new_n690), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n695), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n702), .A2(KEYINPUT90), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(KEYINPUT90), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(G399));
  NOR2_X1   g0505(.A1(new_n534), .A2(G116), .ZN(new_n706));
  INV_X1    g0506(.A(new_n207), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(new_n709), .A3(G1), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n210), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n664), .A2(new_n675), .A3(new_n677), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT26), .ZN(new_n715));
  INV_X1    g0515(.A(new_n672), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n561), .A2(new_n676), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n715), .A2(new_n717), .A3(new_n679), .A4(new_n668), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n713), .B1(new_n718), .B2(new_n690), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n680), .A2(new_n713), .A3(new_n690), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n517), .A2(new_n595), .A3(new_n639), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT91), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n561), .A4(new_n690), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT91), .B1(new_n640), .B2(new_n689), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n509), .A2(new_n510), .ZN(new_n728));
  AND4_X1   g0528(.A1(G179), .A2(new_n556), .A3(new_n583), .A4(new_n633), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NOR4_X1   g0531(.A1(new_n480), .A2(new_n633), .A3(new_n586), .A4(G179), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n730), .A2(new_n731), .B1(new_n531), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(KEYINPUT30), .A3(new_n729), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT31), .B1(new_n735), .B2(new_n689), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n737), .B(new_n690), .C1(new_n733), .C2(new_n734), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n722), .B1(new_n727), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n721), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n712), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n693), .A2(G330), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n262), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n265), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n708), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n746), .A2(new_n694), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n212), .B1(G20), .B2(new_n341), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n213), .A2(G179), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G190), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT32), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n213), .A2(new_n380), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n393), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n393), .A2(G200), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n213), .B1(new_n764), .B2(new_n380), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n759), .B1(new_n201), .B2(new_n763), .C1(new_n224), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n760), .A2(G190), .A3(new_n438), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n760), .A2(new_n755), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n330), .B1(new_n202), .B2(new_n767), .C1(new_n771), .C2(new_n217), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n754), .A2(G190), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n433), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n761), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n754), .A2(new_n393), .A3(G200), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n253), .B1(new_n777), .B2(new_n219), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n766), .A2(new_n772), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n325), .B1(new_n621), .B2(new_n773), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT94), .ZN(new_n781));
  INV_X1    g0581(.A(new_n768), .ZN(new_n782));
  INV_X1    g0582(.A(new_n756), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G311), .A2(new_n782), .B1(new_n783), .B2(G329), .ZN(new_n784));
  INV_X1    g0584(.A(G322), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n785), .B2(new_n767), .ZN(new_n786));
  INV_X1    g0586(.A(G326), .ZN(new_n787));
  INV_X1    g0587(.A(G283), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n763), .A2(new_n787), .B1(new_n777), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI22_X1  g0590(.A1(new_n776), .A2(new_n790), .B1(new_n579), .B2(new_n765), .ZN(new_n791));
  NOR4_X1   g0591(.A1(new_n781), .A2(new_n786), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n753), .B1(new_n779), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n753), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n612), .A2(new_n707), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n210), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n240), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n330), .A2(new_n207), .ZN(new_n801));
  INV_X1    g0601(.A(G355), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n802), .B1(G116), .B2(new_n207), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n797), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n793), .A2(new_n750), .A3(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT95), .Z(new_n806));
  INV_X1    g0606(.A(new_n796), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n693), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n752), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NAND2_X1  g0610(.A1(new_n680), .A2(new_n690), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n390), .A2(new_n689), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n391), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n391), .A2(new_n394), .A3(new_n812), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n680), .A2(new_n815), .A3(new_n690), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n741), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n750), .B1(new_n819), .B2(new_n741), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n816), .A2(new_n794), .ZN(new_n823));
  INV_X1    g0623(.A(new_n753), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n776), .A2(new_n348), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n763), .A2(new_n826), .B1(new_n827), .B2(new_n767), .ZN(new_n828));
  INV_X1    g0628(.A(new_n771), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n825), .B(new_n828), .C1(new_n829), .C2(G159), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT34), .Z(new_n831));
  AOI21_X1  g0631(.A(new_n410), .B1(new_n783), .B2(G132), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n765), .A2(new_n202), .B1(new_n773), .B2(new_n201), .ZN(new_n833));
  INV_X1    g0633(.A(new_n777), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(G68), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n765), .A2(new_n224), .B1(new_n767), .B2(new_n579), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT96), .Z(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n325), .B1(new_n839), .B2(new_n756), .C1(new_n771), .C2(new_n599), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n788), .A2(new_n776), .B1(new_n763), .B2(new_n621), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n433), .A2(new_n777), .B1(new_n773), .B2(new_n219), .ZN(new_n842));
  OR4_X1    g0642(.A1(new_n838), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n824), .B1(new_n836), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n753), .A2(new_n794), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n751), .B(new_n844), .C1(new_n217), .C2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  AOI21_X1  g0648(.A(new_n816), .B1(new_n727), .B2(new_n739), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n271), .A2(new_n689), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n322), .A2(new_n400), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(G169), .B1(new_n303), .B2(new_n309), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT14), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n318), .A3(new_n310), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n271), .B(new_n689), .C1(new_n854), .C2(new_n648), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  INV_X1    g0657(.A(new_n687), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n447), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n642), .A2(new_n859), .A3(new_n860), .A4(new_n441), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n426), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n415), .A2(KEYINPUT16), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n864), .B2(new_n416), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT97), .B1(new_n865), .B2(new_n687), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n415), .A2(KEYINPUT16), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n426), .B1(new_n446), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT97), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n858), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n449), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n866), .A2(new_n870), .A3(new_n441), .A4(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n862), .B1(KEYINPUT37), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n866), .A2(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n451), .A2(KEYINPUT78), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n454), .A3(new_n644), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n441), .B(KEYINPUT17), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n857), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n861), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n881), .B(KEYINPUT38), .C1(new_n455), .C2(new_n874), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n849), .A2(new_n856), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n884), .A2(KEYINPUT99), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT99), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n642), .A2(new_n859), .A3(new_n441), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(new_n860), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n859), .B1(new_n877), .B2(new_n645), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n857), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n849), .A2(new_n856), .A3(new_n893), .A4(KEYINPUT40), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n727), .A2(new_n739), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n456), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n895), .A2(new_n897), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n899), .A2(new_n722), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n879), .A2(new_n882), .A3(KEYINPUT39), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT39), .B1(new_n882), .B2(new_n892), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n854), .A2(new_n271), .A3(new_n690), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n646), .A2(new_n687), .ZN(new_n907));
  INV_X1    g0707(.A(new_n391), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n690), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n818), .A2(new_n909), .B1(new_n851), .B2(new_n855), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n883), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT98), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n721), .B2(new_n457), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n456), .B(KEYINPUT98), .C1(new_n719), .C2(new_n720), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n656), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n912), .B(new_n917), .Z(new_n918));
  OAI22_X1  g0718(.A1(new_n901), .A2(new_n918), .B1(new_n265), .B2(new_n747), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n918), .B2(new_n901), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(G116), .A3(new_n214), .A4(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT36), .Z(new_n924));
  OAI211_X1 g0724(.A(new_n211), .B(G77), .C1(new_n202), .C2(new_n253), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n201), .A2(G68), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n265), .B(G13), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  OR3_X1    g0727(.A1(new_n920), .A2(new_n924), .A3(new_n927), .ZN(G367));
  OAI21_X1  g0728(.A(new_n689), .B1(new_n501), .B2(new_n507), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n517), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n672), .B1(new_n930), .B2(new_n665), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(KEYINPUT100), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n689), .B1(new_n931), .B2(KEYINPUT100), .ZN(new_n933));
  INV_X1    g0733(.A(new_n698), .ZN(new_n934));
  INV_X1    g0734(.A(new_n701), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n716), .A2(new_n689), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n932), .A2(new_n933), .B1(new_n938), .B2(KEYINPUT42), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n546), .A2(new_n689), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n664), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n679), .B2(new_n941), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n939), .A2(new_n940), .B1(KEYINPUT43), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n699), .A2(new_n937), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n708), .B(KEYINPUT41), .Z(new_n949));
  NOR2_X1   g0749(.A1(new_n703), .A2(new_n704), .ZN(new_n950));
  INV_X1    g0750(.A(new_n937), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT45), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n703), .A2(new_n704), .A3(new_n937), .ZN(new_n955));
  XOR2_X1   g0755(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n956));
  OR2_X1    g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n950), .A2(new_n951), .A3(new_n956), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n699), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n698), .B(new_n935), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(new_n694), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n742), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n953), .A2(new_n700), .A3(new_n958), .A4(new_n957), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n949), .B1(new_n965), .B2(new_n743), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n948), .B1(new_n966), .B2(new_n749), .ZN(new_n967));
  INV_X1    g0767(.A(new_n798), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n797), .B1(new_n207), .B2(new_n383), .C1(new_n968), .C2(new_n236), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n750), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT102), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n827), .A2(new_n763), .B1(new_n776), .B2(new_n757), .ZN(new_n972));
  INV_X1    g0772(.A(new_n773), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n972), .B1(G58), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n829), .A2(G50), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n767), .A2(new_n348), .B1(new_n756), .B2(new_n826), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n325), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n765), .A2(new_n253), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G77), .B2(new_n834), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n975), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n579), .A2(new_n776), .B1(new_n763), .B2(new_n839), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n765), .A2(new_n219), .B1(new_n777), .B2(new_n491), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n773), .A2(new_n599), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n829), .B2(G283), .ZN(new_n986));
  INV_X1    g0786(.A(G317), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n410), .B1(new_n756), .B2(new_n987), .C1(new_n767), .C2(new_n621), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(KEYINPUT46), .B2(new_n984), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n983), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT47), .B1(new_n980), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n824), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n980), .A2(KEYINPUT47), .A3(new_n990), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n971), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n943), .B2(new_n807), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n967), .A2(new_n995), .ZN(G387));
  INV_X1    g0796(.A(new_n963), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n742), .A2(new_n962), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n708), .A3(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n801), .A2(new_n706), .B1(G107), .B2(new_n207), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n706), .B(new_n469), .C1(new_n253), .C2(new_n217), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT103), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n386), .A2(G50), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT50), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n968), .B1(new_n233), .B2(G45), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1000), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n797), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n750), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n767), .A2(new_n201), .B1(new_n768), .B2(new_n253), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G150), .B2(new_n783), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n765), .A2(new_n383), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G77), .B2(new_n973), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n353), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G159), .A2(new_n762), .B1(new_n775), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n410), .B1(new_n834), .B2(G97), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n839), .A2(new_n776), .B1(new_n763), .B2(new_n785), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT104), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n767), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n829), .A2(G303), .B1(G317), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(KEYINPUT104), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n765), .A2(new_n788), .B1(new_n773), .B2(new_n579), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n410), .B1(new_n756), .B2(new_n787), .C1(new_n599), .C2(new_n777), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT105), .Z(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT49), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1019), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT106), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n824), .B1(new_n1035), .B2(KEYINPUT106), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1011), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n934), .B2(new_n807), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT107), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n999), .B(new_n1040), .C1(new_n748), .C2(new_n962), .ZN(G393));
  NAND2_X1  g0841(.A1(new_n960), .A2(new_n964), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n997), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(new_n708), .A3(new_n965), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n960), .A2(new_n749), .A3(new_n964), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n797), .B1(new_n207), .B2(new_n491), .C1(new_n968), .C2(new_n243), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n750), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G150), .A2(new_n762), .B1(new_n1022), .B2(G159), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n612), .B1(new_n827), .B2(new_n756), .C1(new_n771), .C2(new_n386), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n776), .A2(new_n201), .B1(new_n777), .B2(new_n433), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n765), .A2(new_n217), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n253), .B2(new_n773), .ZN(new_n1054));
  OR4_X1    g0854(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G317), .A2(new_n762), .B1(new_n1022), .B2(G311), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT108), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT52), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G294), .A2(new_n782), .B1(new_n783), .B2(G322), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n776), .A2(new_n621), .B1(new_n773), .B2(new_n788), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n765), .A2(new_n599), .B1(new_n777), .B2(new_n219), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1058), .A2(new_n325), .A3(new_n1059), .A4(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1057), .A2(KEYINPUT52), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1055), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1047), .B1(new_n1065), .B2(new_n753), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n937), .B2(new_n807), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1045), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1044), .A2(new_n1068), .ZN(G390));
  OAI21_X1  g0869(.A(KEYINPUT110), .B1(new_n457), .B2(new_n741), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT110), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n456), .A2(new_n740), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n916), .A2(new_n1073), .A3(new_n656), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n896), .A2(G330), .A3(new_n815), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n856), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n909), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n717), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(KEYINPUT26), .B2(new_n714), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n668), .A2(new_n679), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n689), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1079), .B1(new_n1083), .B2(new_n815), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT109), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n856), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n851), .A2(new_n855), .A3(KEYINPUT109), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n1075), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1078), .A2(new_n1084), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n818), .A2(new_n909), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT111), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n856), .B1(new_n740), .B2(new_n815), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1075), .A2(KEYINPUT111), .A3(new_n1076), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1089), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n905), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n910), .A2(new_n1097), .B1(new_n902), .B2(new_n903), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1084), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n893), .A2(new_n905), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1077), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1098), .B(new_n1078), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1074), .A2(new_n1096), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1104), .A2(new_n708), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1074), .A2(new_n1096), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(KEYINPUT112), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT112), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1105), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n904), .A2(new_n794), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n774), .B1(G68), .B2(new_n834), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1022), .A2(G116), .B1(new_n783), .B2(G294), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n325), .A3(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1053), .B1(new_n763), .B2(new_n788), .C1(new_n219), .C2(new_n776), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n488), .C2(new_n829), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT53), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n773), .A2(new_n348), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n771), .A2(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1022), .A2(G132), .B1(new_n783), .B2(G125), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1120), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n330), .A3(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n776), .A2(new_n826), .B1(new_n777), .B2(new_n201), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n763), .A2(new_n1127), .B1(new_n757), .B2(new_n765), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1122), .A2(new_n1125), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n753), .B1(new_n1118), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n845), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n750), .C1(new_n1016), .C2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT113), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1113), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1107), .B2(new_n748), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1112), .A2(new_n1137), .ZN(G378));
  AND2_X1   g0938(.A1(new_n894), .A2(G330), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n886), .B2(new_n887), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT115), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(KEYINPUT115), .B(new_n1139), .C1(new_n886), .C2(new_n887), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n359), .A2(new_n687), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n371), .B(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1143), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n912), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n888), .A2(KEYINPUT115), .A3(new_n1139), .A4(new_n1147), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1104), .A2(new_n1074), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n912), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1104), .B2(new_n1074), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n708), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1156), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1147), .A2(new_n794), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n750), .B1(new_n1131), .B2(G50), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n612), .A2(G41), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1022), .A2(G107), .B1(new_n782), .B2(new_n384), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n788), .B2(new_n756), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n978), .B(new_n1171), .C1(G77), .C2(new_n973), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n834), .A2(G58), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G97), .A2(new_n775), .B1(new_n762), .B2(G116), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1167), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1169), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n775), .A2(G132), .B1(new_n782), .B2(G137), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT114), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n767), .A2(new_n1127), .B1(new_n773), .B2(new_n1119), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n762), .A2(G125), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n348), .B2(new_n765), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n834), .A2(G159), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1177), .B1(new_n1176), .B2(new_n1175), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1166), .B1(new_n1190), .B2(new_n753), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1154), .B2(new_n749), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1164), .A2(new_n1194), .ZN(G375));
  NAND3_X1  g0995(.A1(new_n1086), .A2(new_n794), .A3(new_n1087), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n829), .A2(G107), .B1(G116), .B2(new_n775), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT116), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n217), .A2(new_n777), .B1(new_n773), .B2(new_n224), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n325), .B1(new_n621), .B2(new_n756), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G294), .C2(new_n762), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1197), .A2(KEYINPUT116), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1014), .B1(G283), .B2(new_n1022), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT117), .Z(new_n1204));
  NAND4_X1  g1004(.A1(new_n1198), .A2(new_n1201), .A3(new_n1202), .A4(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n612), .B1(new_n826), .B2(new_n767), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1173), .B1(new_n776), .B2(new_n1119), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G132), .C2(new_n762), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n773), .A2(new_n757), .B1(new_n756), .B2(new_n1127), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT119), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n765), .A2(new_n201), .B1(new_n768), .B2(new_n348), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT118), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n824), .B1(new_n1205), .B2(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n751), .B(new_n1214), .C1(new_n253), .C2(new_n845), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1096), .A2(new_n749), .B1(new_n1196), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n949), .B1(new_n1074), .B2(new_n1096), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1074), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1096), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1217), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G381));
  INV_X1    g1023(.A(G390), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT120), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT120), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1228), .A2(G387), .A3(G381), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1112), .A2(new_n1137), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1194), .A4(new_n1164), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT121), .ZN(G407));
  INV_X1    g1032(.A(G213), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(G343), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT122), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G375), .C2(new_n1236), .ZN(G409));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G378), .B(new_n1194), .C1(new_n1156), .C2(new_n1163), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n949), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1158), .A2(new_n1240), .A3(new_n1155), .A4(new_n1159), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1158), .A2(new_n749), .A3(new_n1159), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n1192), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1230), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1234), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1106), .A2(new_n708), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1221), .A2(KEYINPUT60), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1074), .A2(new_n1096), .A3(KEYINPUT60), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1247), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n847), .B1(new_n1251), .B2(new_n1217), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(new_n1249), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G384), .B(new_n1216), .C1(new_n1255), .C2(new_n1247), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1245), .A2(new_n1246), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1235), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1259), .A2(new_n1260), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  XOR2_X1   g1063(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1252), .A2(new_n1256), .B1(G2897), .B2(new_n1235), .ZN(new_n1266));
  INV_X1    g1066(.A(G2897), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1246), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1266), .B1(new_n1258), .B2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1265), .B1(new_n1269), .B2(new_n1261), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1238), .B1(new_n1263), .B2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G390), .A2(new_n967), .A3(new_n995), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT123), .B1(G387), .B2(new_n1224), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G393), .B(new_n809), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1224), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1278), .B1(new_n1280), .B2(KEYINPUT123), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1272), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1277), .A2(new_n1281), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1234), .B(new_n1257), .C1(new_n1239), .C2(new_n1244), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1284), .B1(new_n1285), .B2(KEYINPUT62), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1235), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1245), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1266), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1268), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(new_n1257), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1264), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1286), .A2(KEYINPUT126), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1271), .A2(new_n1283), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1282), .A2(new_n1278), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1285), .A2(KEYINPUT63), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1261), .A2(KEYINPUT63), .A3(new_n1258), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1291), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1294), .A2(new_n1302), .ZN(G405));
  NAND2_X1  g1103(.A1(G375), .A2(new_n1230), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1239), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(KEYINPUT127), .A3(new_n1258), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1258), .A2(KEYINPUT127), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1239), .A3(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1283), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1283), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


