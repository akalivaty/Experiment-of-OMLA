

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n313), .B(G15GAT), .ZN(n322) );
  NOR2_X1 U325 ( .A1(n518), .A2(n528), .ZN(n424) );
  XNOR2_X1 U326 ( .A(n322), .B(n351), .ZN(n323) );
  NOR2_X1 U327 ( .A1(n532), .A2(n443), .ZN(n567) );
  XNOR2_X1 U328 ( .A(KEYINPUT91), .B(KEYINPUT25), .ZN(n450) );
  XNOR2_X1 U329 ( .A(n451), .B(n450), .ZN(n454) );
  NOR2_X1 U330 ( .A1(n568), .A2(n411), .ZN(n413) );
  XNOR2_X1 U331 ( .A(n401), .B(n400), .ZN(n402) );
  INV_X1 U332 ( .A(n556), .ZN(n465) );
  XNOR2_X1 U333 ( .A(n403), .B(n402), .ZN(n406) );
  NOR2_X1 U334 ( .A1(n587), .A2(n465), .ZN(n466) );
  NOR2_X1 U335 ( .A1(n460), .A2(n574), .ZN(n442) );
  XOR2_X1 U336 ( .A(KEYINPUT41), .B(n579), .Z(n552) );
  INV_X1 U337 ( .A(G183GAT), .ZN(n445) );
  XNOR2_X1 U338 ( .A(n445), .B(KEYINPUT122), .ZN(n446) );
  XNOR2_X1 U339 ( .A(n472), .B(G36GAT), .ZN(n473) );
  XNOR2_X1 U340 ( .A(n447), .B(n446), .ZN(G1350GAT) );
  XNOR2_X1 U341 ( .A(n474), .B(n473), .ZN(G1329GAT) );
  XOR2_X1 U342 ( .A(G1GAT), .B(G127GAT), .Z(n427) );
  XOR2_X1 U343 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n293) );
  XNOR2_X1 U344 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n296) );
  XOR2_X1 U346 ( .A(G22GAT), .B(G15GAT), .Z(n387) );
  XNOR2_X1 U347 ( .A(n387), .B(G155GAT), .ZN(n294) );
  XNOR2_X1 U348 ( .A(n294), .B(G64GAT), .ZN(n295) );
  XOR2_X1 U349 ( .A(n296), .B(n295), .Z(n302) );
  XOR2_X1 U350 ( .A(KEYINPUT75), .B(G211GAT), .Z(n298) );
  XNOR2_X1 U351 ( .A(G8GAT), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n352) );
  XOR2_X1 U353 ( .A(KEYINPUT13), .B(G57GAT), .Z(n300) );
  XNOR2_X1 U354 ( .A(G71GAT), .B(G78GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n404) );
  XNOR2_X1 U356 ( .A(n352), .B(n404), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U358 ( .A(n427), .B(n303), .Z(n305) );
  NAND2_X1 U359 ( .A1(G231GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n556) );
  XNOR2_X1 U361 ( .A(KEYINPUT112), .B(n556), .ZN(n540) );
  XOR2_X1 U362 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n307) );
  XNOR2_X1 U363 ( .A(G127GAT), .B(G176GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n328) );
  XOR2_X1 U365 ( .A(KEYINPUT78), .B(G183GAT), .Z(n309) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(G134GAT), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U368 ( .A(G190GAT), .B(G99GAT), .Z(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n324) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n312), .B(G120GAT), .ZN(n436) );
  XOR2_X1 U372 ( .A(G71GAT), .B(n436), .Z(n313) );
  XNOR2_X1 U373 ( .A(KEYINPUT80), .B(KEYINPUT17), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n314), .B(KEYINPUT19), .ZN(n317) );
  INV_X1 U375 ( .A(n317), .ZN(n315) );
  NAND2_X1 U376 ( .A1(n315), .A2(KEYINPUT79), .ZN(n319) );
  INV_X1 U377 ( .A(KEYINPUT79), .ZN(n316) );
  NAND2_X1 U378 ( .A1(n317), .A2(n316), .ZN(n318) );
  NAND2_X1 U379 ( .A1(n319), .A2(n318), .ZN(n321) );
  XNOR2_X1 U380 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n351) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n326) );
  NAND2_X1 U383 ( .A1(G227GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X2 U385 ( .A(n328), .B(n327), .Z(n532) );
  XOR2_X1 U386 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n330) );
  XNOR2_X1 U387 ( .A(KEYINPUT3), .B(KEYINPUT84), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(n331), .B(G155GAT), .Z(n333) );
  XNOR2_X1 U390 ( .A(G141GAT), .B(G148GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n440) );
  XOR2_X1 U392 ( .A(G197GAT), .B(KEYINPUT21), .Z(n356) );
  XOR2_X1 U393 ( .A(n356), .B(KEYINPUT82), .Z(n337) );
  XOR2_X1 U394 ( .A(G106GAT), .B(G162GAT), .Z(n335) );
  XNOR2_X1 U395 ( .A(G50GAT), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n363) );
  XNOR2_X1 U397 ( .A(n363), .B(KEYINPUT23), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U399 ( .A(G204GAT), .B(G78GAT), .Z(n339) );
  NAND2_X1 U400 ( .A1(G228GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U402 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U403 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n343) );
  XNOR2_X1 U404 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n342) );
  XNOR2_X1 U405 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n344), .B(G211GAT), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n440), .B(n347), .ZN(n460) );
  XOR2_X1 U409 ( .A(G92GAT), .B(G64GAT), .Z(n349) );
  XNOR2_X1 U410 ( .A(G204GAT), .B(KEYINPUT71), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U412 ( .A(G176GAT), .B(n350), .ZN(n407) );
  XOR2_X1 U413 ( .A(n351), .B(n407), .Z(n360) );
  XOR2_X1 U414 ( .A(G36GAT), .B(G190GAT), .Z(n364) );
  XOR2_X1 U415 ( .A(n352), .B(n364), .Z(n354) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U418 ( .A(n355), .B(KEYINPUT88), .Z(n358) );
  XNOR2_X1 U419 ( .A(G218GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n518) );
  XNOR2_X1 U422 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n361), .B(KEYINPUT7), .ZN(n391) );
  INV_X1 U424 ( .A(n391), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n377) );
  XOR2_X1 U426 ( .A(G99GAT), .B(G85GAT), .Z(n399) );
  XOR2_X1 U427 ( .A(n364), .B(n399), .Z(n366) );
  NAND2_X1 U428 ( .A1(G232GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U430 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n368) );
  XNOR2_X1 U431 ( .A(G92GAT), .B(KEYINPUT74), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U433 ( .A(n370), .B(n369), .Z(n375) );
  XOR2_X1 U434 ( .A(G29GAT), .B(G134GAT), .Z(n428) );
  XOR2_X1 U435 ( .A(KEYINPUT73), .B(KEYINPUT65), .Z(n372) );
  XNOR2_X1 U436 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n428), .B(n373), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n568) );
  XOR2_X1 U441 ( .A(G1GAT), .B(G113GAT), .Z(n379) );
  XNOR2_X1 U442 ( .A(G169GAT), .B(G141GAT), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U444 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n381) );
  XNOR2_X1 U445 ( .A(G8GAT), .B(KEYINPUT70), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n383), .B(n382), .ZN(n395) );
  XOR2_X1 U448 ( .A(G197GAT), .B(G50GAT), .Z(n385) );
  XNOR2_X1 U449 ( .A(G36GAT), .B(G29GAT), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U451 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U452 ( .A1(G229GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U454 ( .A(n390), .B(KEYINPUT69), .Z(n393) );
  XNOR2_X1 U455 ( .A(n391), .B(KEYINPUT29), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n576) );
  XOR2_X1 U458 ( .A(KEYINPUT31), .B(G106GAT), .Z(n397) );
  XNOR2_X1 U459 ( .A(G120GAT), .B(G148GAT), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U461 ( .A(n399), .B(n398), .Z(n403) );
  NAND2_X1 U462 ( .A1(G230GAT), .A2(G233GAT), .ZN(n401) );
  INV_X1 U463 ( .A(KEYINPUT32), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n404), .B(KEYINPUT33), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n579) );
  INV_X1 U467 ( .A(n552), .ZN(n562) );
  NAND2_X1 U468 ( .A1(n576), .A2(n562), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n409), .B(KEYINPUT46), .ZN(n410) );
  NAND2_X1 U470 ( .A1(n410), .A2(n540), .ZN(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n420) );
  XNOR2_X1 U473 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n416) );
  INV_X1 U474 ( .A(n568), .ZN(n559) );
  XNOR2_X1 U475 ( .A(n559), .B(KEYINPUT96), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n414), .B(KEYINPUT36), .ZN(n587) );
  NOR2_X1 U477 ( .A1(n556), .A2(n587), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n417) );
  NAND2_X1 U479 ( .A1(n579), .A2(n417), .ZN(n418) );
  NOR2_X1 U480 ( .A1(n576), .A2(n418), .ZN(n419) );
  NOR2_X1 U481 ( .A1(n420), .A2(n419), .ZN(n423) );
  XNOR2_X1 U482 ( .A(KEYINPUT64), .B(KEYINPUT114), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n421), .B(KEYINPUT48), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n528) );
  XNOR2_X1 U485 ( .A(n424), .B(KEYINPUT54), .ZN(n441) );
  XOR2_X1 U486 ( .A(KEYINPUT86), .B(KEYINPUT4), .Z(n426) );
  XNOR2_X1 U487 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U489 ( .A(G85GAT), .B(n427), .Z(n430) );
  XNOR2_X1 U490 ( .A(G162GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U492 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U493 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U495 ( .A(n435), .B(KEYINPUT1), .Z(n438) );
  XNOR2_X1 U496 ( .A(n436), .B(KEYINPUT5), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U498 ( .A(n440), .B(n439), .Z(n456) );
  XNOR2_X1 U499 ( .A(KEYINPUT87), .B(n456), .ZN(n514) );
  NAND2_X1 U500 ( .A1(n441), .A2(n514), .ZN(n574) );
  XNOR2_X1 U501 ( .A(n442), .B(KEYINPUT55), .ZN(n443) );
  INV_X1 U502 ( .A(n567), .ZN(n444) );
  NOR2_X1 U503 ( .A1(n540), .A2(n444), .ZN(n447) );
  NAND2_X1 U504 ( .A1(n579), .A2(n576), .ZN(n448) );
  XOR2_X1 U505 ( .A(KEYINPUT72), .B(n448), .Z(n480) );
  NOR2_X1 U506 ( .A1(n532), .A2(n518), .ZN(n449) );
  NOR2_X1 U507 ( .A1(n460), .A2(n449), .ZN(n451) );
  NAND2_X1 U508 ( .A1(n460), .A2(n532), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n452), .B(KEYINPUT26), .ZN(n575) );
  XNOR2_X1 U510 ( .A(n518), .B(KEYINPUT27), .ZN(n458) );
  NOR2_X1 U511 ( .A1(n575), .A2(n458), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT92), .ZN(n457) );
  NOR2_X1 U514 ( .A1(n457), .A2(n456), .ZN(n464) );
  NOR2_X1 U515 ( .A1(n458), .A2(n514), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT89), .ZN(n527) );
  XOR2_X1 U517 ( .A(KEYINPUT28), .B(n460), .Z(n530) );
  NAND2_X1 U518 ( .A1(n532), .A2(n530), .ZN(n461) );
  NOR2_X1 U519 ( .A1(n527), .A2(n461), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT90), .ZN(n463) );
  NOR2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n477) );
  INV_X1 U522 ( .A(n477), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(KEYINPUT37), .Z(n468) );
  XNOR2_X1 U525 ( .A(n469), .B(n468), .ZN(n513) );
  NAND2_X1 U526 ( .A1(n480), .A2(n513), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT98), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n471), .B(KEYINPUT38), .ZN(n496) );
  NOR2_X1 U529 ( .A1(n518), .A2(n496), .ZN(n474) );
  INV_X1 U530 ( .A(KEYINPUT100), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n476) );
  NAND2_X1 U532 ( .A1(n559), .A2(n465), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(n478) );
  NOR2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n479) );
  XOR2_X1 U535 ( .A(n479), .B(KEYINPUT93), .Z(n500) );
  NAND2_X1 U536 ( .A1(n500), .A2(n480), .ZN(n487) );
  NOR2_X1 U537 ( .A1(n514), .A2(n487), .ZN(n481) );
  XOR2_X1 U538 ( .A(n481), .B(KEYINPUT34), .Z(n482) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n518), .A2(n487), .ZN(n483) );
  XOR2_X1 U541 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  NOR2_X1 U542 ( .A1(n532), .A2(n487), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U546 ( .A1(n530), .A2(n487), .ZN(n488) );
  XOR2_X1 U547 ( .A(G22GAT), .B(n488), .Z(G1327GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n490) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT95), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n492) );
  NOR2_X1 U551 ( .A1(n514), .A2(n496), .ZN(n491) );
  XOR2_X1 U552 ( .A(n492), .B(n491), .Z(G1328GAT) );
  INV_X1 U553 ( .A(KEYINPUT40), .ZN(n494) );
  NOR2_X1 U554 ( .A1(n532), .A2(n496), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U557 ( .A1(n530), .A2(n496), .ZN(n498) );
  XNOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  NOR2_X1 U561 ( .A1(n576), .A2(n552), .ZN(n512) );
  AND2_X1 U562 ( .A1(n512), .A2(n500), .ZN(n501) );
  XOR2_X1 U563 ( .A(KEYINPUT104), .B(n501), .Z(n508) );
  NOR2_X1 U564 ( .A1(n514), .A2(n508), .ZN(n505) );
  XOR2_X1 U565 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n503) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT105), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n518), .A2(n508), .ZN(n506) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n532), .A2(n508), .ZN(n507) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n508), .A2(n530), .ZN(n510) );
  XNOR2_X1 U574 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n523) );
  NOR2_X1 U578 ( .A1(n514), .A2(n523), .ZN(n516) );
  XNOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n523), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NOR2_X1 U585 ( .A1(n532), .A2(n523), .ZN(n521) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(n521), .Z(n522) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NOR2_X1 U588 ( .A1(n530), .A2(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n534) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(n529), .B(KEYINPUT115), .Z(n548) );
  NAND2_X1 U595 ( .A1(n548), .A2(n530), .ZN(n531) );
  NOR2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n576), .A2(n544), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U600 ( .A1(n544), .A2(n562), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT117), .Z(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  INV_X1 U604 ( .A(n544), .ZN(n539) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U610 ( .A1(n544), .A2(n568), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  INV_X1 U612 ( .A(n576), .ZN(n549) );
  INV_X1 U613 ( .A(n575), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n558) );
  NOR2_X1 U615 ( .A1(n549), .A2(n558), .ZN(n550) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n550), .Z(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT120), .B(n551), .ZN(G1344GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n558), .ZN(n554) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n558), .ZN(n557) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n567), .A2(n576), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n564) );
  NAND2_X1 U629 ( .A1(n567), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .Z(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(n573), .Z(n578) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n583), .A2(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U644 ( .A(n583), .ZN(n586) );
  OR2_X1 U645 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT126), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n583), .A2(n465), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

