//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  NOR2_X1   g000(.A1(KEYINPUT2), .A2(G113), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT2), .A2(G113), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT68), .ZN(new_n189));
  OR2_X1    g003(.A1(new_n188), .A2(KEYINPUT68), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(KEYINPUT69), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n195), .B2(new_n191), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT72), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT72), .B(new_n193), .C1(new_n195), .C2(new_n191), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT65), .B(G146), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n203), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(G146), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n207), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  OAI21_X1  g029(.A(G128), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n201), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(G128), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n218), .B(new_n220), .C1(new_n206), .C2(new_n207), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n211), .A2(new_n213), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G143), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n225), .A2(KEYINPUT67), .A3(new_n218), .A4(new_n220), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n210), .A2(new_n216), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G137), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(G137), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n229), .A2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(G131), .C1(new_n239), .C2(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT71), .B1(new_n227), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n217), .B1(new_n224), .B2(G143), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT0), .A3(G128), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  OR2_X1    g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n211), .A2(new_n213), .A3(new_n207), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n209), .B1(new_n247), .B2(KEYINPUT64), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n245), .B(new_n246), .C1(new_n248), .C2(new_n204), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n234), .A2(G131), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n235), .A2(new_n250), .A3(KEYINPUT70), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT70), .B1(new_n235), .B2(new_n250), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n244), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n223), .A2(new_n226), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n216), .B1(new_n248), .B2(new_n204), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n257));
  INV_X1    g071(.A(new_n241), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n200), .A2(new_n242), .A3(new_n253), .A4(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n262), .B(KEYINPUT27), .Z(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT26), .ZN(new_n264));
  INV_X1    g078(.A(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n235), .A2(new_n250), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n249), .A2(new_n267), .A3(new_n244), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n241), .B1(new_n254), .B2(new_n255), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT30), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n242), .A2(new_n253), .A3(new_n259), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(KEYINPUT30), .ZN(new_n272));
  INV_X1    g086(.A(new_n196), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n260), .B(new_n266), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n196), .B1(new_n268), .B2(new_n269), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n260), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT28), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n251), .A2(new_n252), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n249), .A2(new_n244), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n269), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT28), .B1(new_n285), .B2(new_n200), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n266), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n274), .A2(KEYINPUT73), .A3(KEYINPUT31), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n277), .A2(new_n278), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G472), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n292), .A2(KEYINPUT32), .A3(new_n293), .A4(new_n294), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT74), .B1(new_n288), .B2(new_n289), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n260), .B1(new_n272), .B2(new_n273), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n289), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n281), .A2(new_n303), .A3(new_n266), .A4(new_n287), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n299), .A2(new_n300), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n306));
  INV_X1    g120(.A(new_n200), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n271), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n308), .B2(new_n260), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(new_n286), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n289), .A2(new_n300), .ZN(new_n311));
  AOI21_X1  g125(.A(G902), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G472), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n297), .A2(new_n298), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G128), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n318), .A2(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(KEYINPUT23), .ZN(new_n320));
  INV_X1    g134(.A(G128), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n319), .B(new_n320), .C1(G119), .C2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G119), .B(G128), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT24), .B(G110), .Z(new_n324));
  OAI22_X1  g138(.A1(new_n322), .A2(G110), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G146), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n327), .A2(new_n329), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n325), .B(new_n332), .C1(new_n206), .C2(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n322), .A2(G110), .B1(new_n323), .B2(new_n324), .ZN(new_n335));
  INV_X1    g149(.A(new_n332), .ZN(new_n336));
  AOI21_X1  g150(.A(G146), .B1(new_n330), .B2(new_n331), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT22), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(G137), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(KEYINPUT76), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n344), .B(new_n294), .C1(new_n339), .C2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G217), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(G234), .B2(new_n294), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n346), .A2(new_n348), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT77), .B1(new_n346), .B2(new_n348), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n349), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n351), .A2(G902), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n344), .B(new_n355), .C1(new_n339), .C2(new_n345), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n315), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n315), .A2(KEYINPUT78), .A3(new_n357), .ZN(new_n361));
  INV_X1    g175(.A(G469), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n251), .A2(new_n252), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G104), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(KEYINPUT82), .A3(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(KEYINPUT79), .A2(G107), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT79), .A2(G107), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n371), .A2(new_n372), .A3(G104), .ZN(new_n373));
  OAI21_X1  g187(.A(G101), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n365), .A2(G104), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(KEYINPUT3), .B2(new_n366), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(G104), .C1(new_n371), .C2(new_n372), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n265), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT67), .B1(new_n243), .B2(new_n220), .ZN(new_n382));
  NOR4_X1   g196(.A1(new_n214), .A2(new_n222), .A3(new_n217), .A4(new_n219), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n321), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT83), .B1(new_n243), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G128), .B1(new_n209), .B2(new_n215), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n387), .B(new_n388), .C1(new_n214), .C2(new_n217), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n381), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n254), .A2(new_n255), .A3(new_n380), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n364), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT84), .B1(new_n393), .B2(KEYINPUT12), .ZN(new_n394));
  INV_X1    g208(.A(new_n389), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n218), .B1(new_n206), .B2(new_n207), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n388), .B1(new_n396), .B2(new_n387), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n380), .B1(new_n398), .B2(new_n254), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n254), .A2(new_n255), .A3(new_n380), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n282), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT84), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT12), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT12), .B(new_n267), .C1(new_n399), .C2(new_n400), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n394), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT10), .B1(new_n227), .B2(new_n380), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(new_n381), .C1(new_n384), .C2(new_n390), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n265), .B1(new_n376), .B2(new_n378), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT4), .A3(new_n379), .ZN(new_n413));
  INV_X1    g227(.A(new_n375), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n366), .A2(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n378), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n417), .A3(G101), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(KEYINPUT80), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(new_n411), .B2(new_n417), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n413), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n422), .A2(new_n423), .A3(new_n283), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(KEYINPUT80), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n411), .A2(new_n420), .A3(new_n417), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n379), .A2(KEYINPUT4), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n425), .A2(new_n426), .B1(new_n427), .B2(new_n412), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT81), .B1(new_n428), .B2(new_n284), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n364), .B(new_n410), .C1(new_n424), .C2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n340), .A2(G227), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n363), .B1(new_n406), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n433), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n423), .B1(new_n422), .B2(new_n283), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n428), .A2(KEYINPUT81), .A3(new_n284), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n437), .A2(new_n438), .B1(new_n407), .B2(new_n409), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n439), .B2(new_n364), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n394), .A2(new_n404), .A3(new_n405), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(KEYINPUT87), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n410), .B1(new_n424), .B2(new_n429), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT86), .B(new_n410), .C1(new_n424), .C2(new_n429), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n282), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n433), .B1(new_n448), .B2(new_n430), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n362), .B(new_n294), .C1(new_n443), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(G469), .A2(G902), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n440), .A2(KEYINPUT85), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n434), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n448), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n441), .A2(new_n430), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n436), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(G469), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n451), .A3(new_n458), .ZN(new_n459));
  XOR2_X1   g273(.A(KEYINPUT9), .B(G234), .Z(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G221), .B1(new_n461), .B2(G902), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G214), .B1(G237), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n428), .A2(new_n196), .ZN(new_n466));
  INV_X1    g280(.A(G113), .ZN(new_n467));
  INV_X1    g281(.A(G116), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G119), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT5), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n194), .B2(new_n470), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n381), .A2(new_n472), .A3(new_n193), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n466), .A2(new_n473), .A3(new_n475), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n227), .A2(new_n328), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n283), .A2(G125), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(G224), .A3(new_n340), .ZN(new_n483));
  INV_X1    g297(.A(G224), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n480), .B(new_n481), .C1(new_n484), .C2(G953), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n474), .A2(new_n487), .A3(new_n476), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n479), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n472), .A2(new_n193), .A3(new_n380), .ZN(new_n490));
  INV_X1    g304(.A(new_n192), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n471), .B1(new_n491), .B2(new_n470), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n380), .B1(new_n193), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n475), .B(KEYINPUT8), .Z(new_n494));
  NOR3_X1   g308(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n482), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n485), .A2(new_n496), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n478), .A4(new_n483), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n294), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n489), .A2(new_n294), .A3(new_n501), .A4(new_n499), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n465), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(G234), .A2(G237), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(G952), .A3(new_n340), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT21), .B(G898), .Z(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n506), .A2(G902), .A3(G953), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n461), .A2(new_n350), .A3(G953), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n321), .B2(G143), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n207), .A2(KEYINPUT93), .A3(G128), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT13), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n520), .A2(new_n521), .B1(new_n321), .B2(G143), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n521), .B2(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G134), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n468), .A2(G122), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT92), .B(G122), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n526), .B2(new_n468), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n371), .A2(new_n372), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n518), .A2(new_n519), .B1(new_n321), .B2(G143), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n229), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n527), .A2(new_n528), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n525), .B(KEYINPUT14), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n526), .A2(new_n468), .ZN(new_n540));
  OAI21_X1  g354(.A(G107), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n530), .A2(new_n229), .ZN(new_n542));
  INV_X1    g356(.A(new_n531), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n538), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n516), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  INV_X1    g360(.A(new_n516), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n546), .B(new_n547), .C1(new_n535), .C2(new_n536), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n294), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G478), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n549), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n336), .A2(new_n337), .ZN(new_n554));
  INV_X1    g368(.A(G237), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n340), .A3(G214), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n207), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND4_X1   g373(.A1(KEYINPUT89), .A2(new_n559), .A3(KEYINPUT17), .A4(G131), .ZN(new_n560));
  INV_X1    g374(.A(G131), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n557), .B2(new_n558), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT89), .B1(new_n562), .B2(KEYINPUT17), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n554), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT90), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n559), .A2(G131), .ZN(new_n567));
  OR3_X1    g381(.A1(new_n567), .A2(KEYINPUT17), .A3(new_n562), .ZN(new_n568));
  OAI211_X1 g382(.A(KEYINPUT90), .B(new_n554), .C1(new_n560), .C2(new_n563), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G113), .B(G122), .ZN(new_n571));
  INV_X1    g385(.A(G104), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n562), .A2(KEYINPUT18), .ZN(new_n574));
  AND2_X1   g388(.A1(KEYINPUT18), .A2(G131), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n333), .B(KEYINPUT88), .Z(new_n576));
  AND2_X1   g390(.A1(new_n576), .A2(G146), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n333), .A2(new_n206), .ZN(new_n578));
  OAI221_X1 g392(.A(new_n574), .B1(new_n559), .B2(new_n575), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n570), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT91), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n570), .A2(new_n579), .A3(KEYINPUT91), .A4(new_n573), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n576), .A2(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(KEYINPUT19), .B2(new_n333), .ZN(new_n586));
  OAI221_X1 g400(.A(new_n332), .B1(new_n562), .B2(new_n567), .C1(new_n586), .C2(new_n206), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n579), .ZN(new_n588));
  INV_X1    g402(.A(new_n573), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G475), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n294), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT20), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n582), .A2(new_n583), .B1(new_n589), .B2(new_n588), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(G475), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT20), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n294), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n573), .B1(new_n570), .B2(new_n579), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n582), .B2(new_n583), .ZN(new_n601));
  OAI21_X1  g415(.A(G475), .B1(new_n601), .B2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n553), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n463), .A2(new_n515), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n360), .A2(new_n361), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  NAND2_X1  g420(.A1(new_n292), .A2(new_n294), .ZN(new_n607));
  NAND2_X1  g421(.A1(KEYINPUT95), .A2(G472), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n459), .A2(new_n462), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n357), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n597), .B1(new_n596), .B2(new_n294), .ZN(new_n612));
  NOR4_X1   g426(.A1(new_n595), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n602), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n537), .A2(new_n544), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n547), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n537), .A2(new_n544), .A3(new_n516), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(KEYINPUT33), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n545), .B2(new_n548), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n618), .A2(new_n620), .A3(G478), .A4(new_n294), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n549), .A2(new_n550), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n611), .A2(new_n515), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  INV_X1    g441(.A(new_n515), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n594), .B2(new_n630), .ZN(new_n631));
  AOI211_X1 g445(.A(KEYINPUT96), .B(KEYINPUT97), .C1(new_n593), .C2(KEYINPUT20), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n598), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n552), .A2(new_n602), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT97), .B1(new_n612), .B2(KEYINPUT96), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n594), .A2(new_n630), .A3(new_n629), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n613), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n628), .A2(new_n633), .A3(new_n634), .A4(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n611), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT98), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT35), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G107), .ZN(G9));
  NOR2_X1   g457(.A1(new_n603), .A2(new_n515), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT36), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n345), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n339), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n355), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n354), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n609), .A2(new_n610), .A3(new_n644), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n508), .B1(new_n512), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n633), .A2(new_n637), .A3(new_n634), .A4(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n505), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n315), .A2(new_n610), .A3(new_n651), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(new_n656), .B(KEYINPUT39), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n610), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n503), .A2(new_n504), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  OR3_X1    g483(.A1(new_n463), .A2(KEYINPUT40), .A3(new_n664), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n301), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n289), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n308), .A2(new_n260), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n294), .B1(new_n674), .B2(new_n266), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n297), .A2(new_n298), .A3(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n650), .A2(new_n354), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n614), .A2(new_n552), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n677), .A2(new_n464), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n671), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n207), .ZN(G45));
  AOI22_X1  g497(.A1(new_n599), .A2(new_n602), .B1(new_n622), .B2(new_n621), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(KEYINPUT100), .A3(new_n505), .A4(new_n657), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n614), .A2(new_n505), .A3(new_n623), .A4(new_n657), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n315), .A3(new_n610), .A4(new_n651), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  AND2_X1   g505(.A1(new_n315), .A2(new_n357), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n624), .A2(new_n515), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n294), .B1(new_n443), .B2(new_n449), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n462), .A3(new_n450), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT101), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n695), .A2(new_n698), .A3(new_n462), .A4(new_n450), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n692), .A2(new_n693), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND3_X1  g517(.A1(new_n692), .A2(new_n638), .A3(new_n700), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  INV_X1    g519(.A(new_n696), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n315), .A2(new_n706), .A3(new_n644), .A4(new_n651), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  NAND2_X1  g522(.A1(new_n674), .A2(KEYINPUT28), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(KEYINPUT102), .A3(new_n287), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n309), .B2(new_n286), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n289), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n278), .A3(new_n275), .ZN(new_n714));
  NOR2_X1   g528(.A1(G472), .A2(G902), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n607), .A2(G472), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n714), .A2(KEYINPUT103), .A3(new_n715), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n357), .A2(new_n718), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n700), .A2(new_n721), .A3(new_n628), .A4(new_n680), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NAND4_X1  g537(.A1(new_n718), .A2(new_n719), .A3(new_n651), .A4(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n684), .A2(new_n657), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n505), .A3(new_n706), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n668), .A2(new_n465), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n729), .B1(new_n463), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n459), .A2(KEYINPUT104), .A3(new_n730), .A4(new_n462), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n725), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n692), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n358), .B1(new_n732), .B2(new_n733), .ZN(new_n740));
  INV_X1    g554(.A(new_n738), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n735), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  INV_X1    g558(.A(new_n658), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n734), .A2(new_n692), .A3(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT106), .B(G134), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G36));
  NAND2_X1  g562(.A1(new_n455), .A2(new_n457), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n455), .A2(KEYINPUT45), .A3(new_n457), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(G469), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n451), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n451), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n450), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n462), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n730), .B(KEYINPUT108), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n664), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n599), .A2(new_n623), .A3(new_n602), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT43), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n609), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n651), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT44), .A4(new_n651), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n772), .A2(KEYINPUT107), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(KEYINPUT107), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n761), .B(new_n771), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  OAI21_X1  g590(.A(new_n759), .B1(KEYINPUT109), .B2(KEYINPUT47), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n315), .A2(new_n357), .ZN(new_n778));
  NOR2_X1   g592(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n779));
  AND2_X1   g593(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n758), .B(new_n462), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n725), .A2(new_n731), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n777), .A2(new_n778), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  AOI21_X1  g598(.A(new_n507), .B1(new_n764), .B2(new_n766), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n721), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n696), .ZN(new_n787));
  INV_X1    g601(.A(new_n669), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n465), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n787), .A2(KEYINPUT50), .A3(new_n465), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n696), .A2(new_n731), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n785), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n724), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n677), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n357), .A3(new_n508), .A4(new_n794), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n614), .A3(new_n623), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n793), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n786), .A2(new_n760), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n695), .A2(new_n450), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(new_n462), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n777), .A2(new_n781), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT114), .B1(new_n777), .B2(new_n781), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT51), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n795), .A2(new_n692), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT48), .ZN(new_n813));
  INV_X1    g627(.A(G952), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n814), .B(G953), .C1(new_n787), .C2(new_n505), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n793), .A2(KEYINPUT51), .A3(new_n797), .A4(new_n801), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n760), .B(new_n786), .C1(new_n806), .C2(new_n805), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n813), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n799), .A2(new_n624), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n811), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n678), .A2(new_n657), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n463), .B1(KEYINPUT111), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n679), .A2(new_n659), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n823), .A2(KEYINPUT111), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n824), .A2(new_n677), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n662), .A2(new_n690), .A3(new_n727), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT112), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n701), .A2(new_n704), .A3(new_n722), .A4(new_n707), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n599), .A2(new_n552), .A3(new_n602), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n515), .B1(new_n624), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n609), .A3(new_n610), .A4(new_n357), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n652), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n605), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n746), .B1(new_n739), .B2(new_n742), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n633), .A2(new_n637), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n553), .A2(new_n602), .A3(new_n657), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n731), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n661), .A2(new_n845), .B1(new_n734), .B2(new_n726), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n822), .B1(new_n833), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n315), .A2(KEYINPUT78), .A3(new_n357), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT78), .B1(new_n315), .B2(new_n357), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n838), .B1(new_n851), .B2(new_n604), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n701), .A2(new_n722), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n704), .A2(new_n707), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n846), .ZN(new_n855));
  INV_X1    g669(.A(new_n746), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n741), .B1(new_n740), .B2(new_n735), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n692), .A2(new_n734), .A3(new_n735), .A4(new_n741), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n828), .A2(KEYINPUT52), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n724), .A2(new_n725), .A3(new_n659), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n660), .A2(new_n661), .B1(new_n862), .B2(new_n706), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n830), .A3(new_n690), .A4(new_n827), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n860), .A2(new_n866), .A3(KEYINPUT53), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n821), .B1(new_n848), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT53), .B1(new_n833), .B2(new_n847), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n860), .A2(new_n866), .A3(new_n822), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT54), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT113), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n828), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT52), .B1(new_n828), .B2(KEYINPUT112), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n875), .B2(new_n860), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n847), .A2(new_n822), .A3(new_n865), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT54), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n822), .B1(new_n875), .B2(new_n860), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n847), .A2(KEYINPUT53), .A3(new_n865), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n821), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT113), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n820), .A2(new_n872), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT115), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n814), .A2(new_n340), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n820), .A2(new_n872), .A3(new_n887), .A4(new_n883), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n804), .A2(KEYINPUT49), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT110), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n788), .A2(new_n357), .A3(new_n462), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n804), .A2(KEYINPUT49), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n892), .A2(new_n893), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n464), .A3(new_n798), .A4(new_n763), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n889), .A2(new_n897), .ZN(G75));
  NAND2_X1  g712(.A1(new_n869), .A2(new_n870), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n294), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n479), .A2(new_n488), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n486), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n901), .A2(new_n904), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n340), .A2(G952), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(G51));
  NAND3_X1  g722(.A1(new_n869), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n881), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n451), .B(KEYINPUT57), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n910), .A2(new_n911), .B1(new_n449), .B2(new_n443), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n753), .B(KEYINPUT116), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n900), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n907), .B1(new_n912), .B2(new_n914), .ZN(G54));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n592), .ZN(new_n918));
  NAND3_X1  g732(.A1(KEYINPUT117), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n900), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n595), .ZN(new_n921));
  INV_X1    g735(.A(new_n907), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n900), .A2(new_n591), .A3(new_n918), .A4(new_n919), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n921), .A2(KEYINPUT118), .A3(new_n922), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n881), .B2(new_n909), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n618), .A2(new_n620), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n907), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n930), .B1(new_n872), .B2(new_n883), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(new_n932), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT119), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n933), .C1(new_n934), .C2(new_n932), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(G63));
  INV_X1    g753(.A(new_n899), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n344), .B1(new_n339), .B2(new_n345), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n907), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n647), .B(KEYINPUT120), .Z(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G66));
  OAI21_X1  g763(.A(G953), .B1(new_n510), .B2(new_n484), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n841), .B2(G953), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n902), .B1(G898), .B2(new_n340), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  AOI21_X1  g767(.A(new_n340), .B1(G227), .B2(G900), .ZN(new_n954));
  NAND2_X1  g768(.A1(G900), .A2(G953), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n272), .B(KEYINPUT121), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n586), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n775), .A2(new_n783), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n759), .A2(new_n664), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n692), .A3(new_n825), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT125), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n960), .A2(new_n963), .A3(new_n692), .A4(new_n825), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n859), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n863), .A2(new_n690), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n959), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n955), .B(new_n957), .C1(new_n967), .C2(G953), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n954), .B1(new_n968), .B2(KEYINPUT124), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT123), .ZN(new_n971));
  INV_X1    g785(.A(new_n957), .ZN(new_n972));
  INV_X1    g786(.A(new_n682), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n966), .A2(KEYINPUT62), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n863), .A2(new_n690), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n682), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n624), .A2(new_n835), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n666), .A2(new_n731), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n851), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(new_n959), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT122), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n978), .A2(new_n959), .A3(KEYINPUT122), .A4(new_n981), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n971), .B(new_n972), .C1(new_n986), .C2(G953), .ZN(new_n987));
  AOI21_X1  g801(.A(G953), .B1(new_n984), .B2(new_n985), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT123), .B1(new_n988), .B2(new_n957), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n970), .B1(new_n990), .B2(new_n968), .ZN(new_n991));
  INV_X1    g805(.A(new_n968), .ZN(new_n992));
  AOI211_X1 g806(.A(new_n992), .B(new_n969), .C1(new_n987), .C2(new_n989), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n991), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  INV_X1    g810(.A(new_n841), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n967), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT126), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n672), .A3(new_n289), .ZN(new_n1000));
  INV_X1    g814(.A(new_n274), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n302), .B(KEYINPUT127), .Z(new_n1002));
  OAI221_X1 g816(.A(new_n996), .B1(new_n1001), .B2(new_n1002), .C1(new_n876), .C2(new_n877), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1000), .A2(new_n922), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n986), .A2(new_n841), .ZN(new_n1005));
  AOI211_X1 g819(.A(new_n672), .B(new_n289), .C1(new_n1005), .C2(new_n996), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1004), .A2(new_n1006), .ZN(G57));
endmodule


