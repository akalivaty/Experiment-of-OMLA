//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT66), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n209), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  AND2_X1   g0028(.A1(new_n228), .A2(new_n211), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n222), .C1(new_n223), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n223), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G107), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G97), .ZN(new_n247));
  INV_X1    g0047(.A(G97), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G107), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n245), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n220), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n208), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G50), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n203), .A2(G20), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(new_n265), .B1(G150), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n256), .A2(new_n220), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n260), .B1(G50), .B2(new_n254), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT72), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G222), .A2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G223), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n278), .B(new_n279), .C1(G77), .C2(new_n274), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT69), .B(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n288), .B2(new_n282), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n279), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n280), .B(new_n286), .C1(new_n287), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G200), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n270), .B2(new_n271), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n294), .A2(KEYINPUT73), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n270), .B(new_n301), .C1(G179), .C2(new_n292), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n258), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n263), .A2(new_n259), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n304), .A2(new_n305), .B1(new_n254), .B2(new_n263), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G58), .A2(G68), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n209), .B1(new_n217), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n209), .A2(new_n264), .ZN(new_n310));
  INV_X1    g0110(.A(G159), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT77), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n308), .ZN(new_n314));
  OAI21_X1  g0114(.A(G20), .B1(new_n314), .B2(new_n202), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n266), .A2(G159), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n274), .B2(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT76), .B1(new_n274), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  INV_X1    g0128(.A(new_n322), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n321), .A2(new_n323), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n319), .B1(G68), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n269), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n324), .A2(KEYINPUT78), .A3(G33), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n329), .C1(new_n327), .C2(KEYINPUT78), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n216), .B1(new_n336), .B2(new_n321), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n334), .B1(new_n337), .B2(new_n319), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT79), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n331), .A2(G68), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n313), .A2(new_n318), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(KEYINPUT16), .A3(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n342), .A2(KEYINPUT79), .A3(new_n338), .A4(new_n257), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n307), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n290), .A2(G232), .ZN(new_n347));
  INV_X1    g0147(.A(new_n279), .ZN(new_n348));
  INV_X1    g0148(.A(G87), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n264), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(G223), .A2(G1698), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n287), .B2(G1698), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n352), .B2(new_n274), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n286), .B(new_n347), .C1(new_n348), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(G169), .B2(new_n354), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n345), .A2(new_n346), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n353), .A2(new_n348), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n362), .A2(new_n295), .A3(new_n286), .A4(new_n347), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n307), .B(new_n365), .C1(new_n339), .C2(new_n344), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT17), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n342), .A2(new_n257), .A3(new_n338), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT79), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n306), .B1(new_n371), .B2(new_n343), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT18), .B1(new_n372), .B2(new_n357), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(KEYINPUT17), .A3(new_n365), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n359), .A2(new_n368), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT74), .B1(new_n254), .B2(G68), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT12), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT11), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n265), .A2(G77), .B1(G20), .B2(new_n216), .ZN(new_n379));
  INV_X1    g0179(.A(G50), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n310), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n257), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n377), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n258), .A2(G68), .A3(new_n259), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n387));
  INV_X1    g0187(.A(G238), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n286), .B1(new_n388), .B2(new_n291), .ZN(new_n389));
  INV_X1    g0189(.A(G232), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n274), .B(new_n391), .C1(G226), .C2(G1698), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G97), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n348), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n389), .A2(new_n394), .A3(KEYINPUT13), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n393), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n279), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n283), .A2(new_n285), .B1(new_n290), .B2(G238), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(G169), .B(new_n387), .C1(new_n395), .C2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT13), .B1(new_n389), .B2(new_n394), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n396), .A3(new_n399), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(G179), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n403), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n387), .B1(new_n406), .B2(G169), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n386), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n395), .A2(new_n400), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n386), .B1(new_n409), .B2(G190), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n360), .B2(new_n409), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G77), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n262), .A2(new_n310), .B1(new_n209), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT70), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT71), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n209), .A2(G33), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n414), .A2(new_n415), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n257), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n413), .B1(new_n208), .B2(G20), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n258), .A2(new_n423), .B1(new_n413), .B2(new_n255), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n274), .A2(new_n276), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n426), .A2(new_n390), .B1(new_n246), .B2(new_n274), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n327), .A2(new_n388), .A3(new_n276), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n279), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n283), .A2(new_n285), .B1(new_n290), .B2(G244), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n300), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n355), .A3(new_n430), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n425), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(G200), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n429), .A2(G190), .A3(new_n430), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n422), .A4(new_n424), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n303), .A2(new_n375), .A3(new_n412), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n208), .A2(G33), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n269), .A2(new_n254), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n254), .A2(G116), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT81), .ZN(new_n447));
  AOI21_X1  g0247(.A(G20), .B1(new_n264), .B2(G97), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n442), .A2(G20), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n257), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT20), .B1(new_n449), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n445), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n274), .A2(G264), .A3(G1698), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n274), .A2(G257), .A3(new_n276), .ZN(new_n458));
  INV_X1    g0258(.A(G303), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(new_n274), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n279), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n208), .B(G45), .C1(new_n462), .C2(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n463), .B1(new_n467), .B2(new_n462), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n285), .ZN(new_n469));
  INV_X1    g0269(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G270), .A3(new_n348), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n461), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n456), .A2(new_n472), .A3(KEYINPUT21), .A4(G169), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n456), .A2(new_n472), .A3(G169), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT21), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(G200), .ZN(new_n477));
  INV_X1    g0277(.A(new_n456), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n461), .A2(G190), .A3(new_n471), .A4(new_n469), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AND4_X1   g0280(.A1(G179), .A2(new_n461), .A3(new_n469), .A4(new_n471), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n456), .ZN(new_n482));
  AND4_X1   g0282(.A1(new_n473), .A2(new_n476), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n266), .A2(G77), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT6), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n247), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g0288(.A(G97), .B(G107), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n486), .B1(new_n490), .B2(new_n209), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n246), .B1(new_n336), .B2(new_n321), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n257), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n254), .A2(G97), .ZN(new_n494));
  AND4_X1   g0294(.A1(new_n220), .A2(new_n254), .A3(new_n256), .A4(new_n440), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n325), .A2(new_n326), .A3(G244), .A4(new_n276), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n276), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n447), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n279), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT5), .B1(new_n464), .B2(new_n466), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n348), .B(G257), .C1(new_n505), .C2(new_n463), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n469), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n295), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n497), .B1(new_n509), .B2(KEYINPUT82), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n360), .B1(new_n504), .B2(new_n507), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT82), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n511), .A2(new_n512), .B1(new_n508), .B2(new_n295), .ZN(new_n513));
  INV_X1    g0313(.A(new_n508), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n355), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n300), .A2(new_n508), .B1(new_n493), .B2(new_n496), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n510), .A2(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n274), .A2(G244), .A3(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n426), .C2(new_n388), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n208), .A2(new_n284), .A3(G45), .ZN(new_n521));
  AOI21_X1  g0321(.A(G250), .B1(new_n208), .B2(G45), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n279), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n520), .A2(new_n279), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n355), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT83), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n527), .A3(new_n355), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n520), .A2(new_n279), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(new_n521), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n300), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n274), .A2(new_n209), .A3(G68), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n419), .A2(new_n248), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(KEYINPUT19), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT84), .B(G87), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n536), .A2(new_n537), .B1(new_n209), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n257), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n418), .A2(new_n255), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n418), .C2(new_n441), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n526), .A2(new_n528), .A3(new_n532), .A4(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT85), .B1(new_n441), .B2(new_n349), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT85), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n495), .A2(new_n545), .A3(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n540), .A2(new_n547), .A3(new_n541), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n524), .A2(G190), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n360), .C2(new_n524), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n483), .A2(new_n517), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n470), .A2(KEYINPUT87), .A3(G264), .A4(new_n348), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n348), .B(G264), .C1(new_n505), .C2(new_n463), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n274), .A2(G257), .A3(G1698), .ZN(new_n558));
  INV_X1    g0358(.A(G294), .ZN(new_n559));
  INV_X1    g0359(.A(G250), .ZN(new_n560));
  OAI221_X1 g0360(.A(new_n558), .B1(new_n264), .B2(new_n559), .C1(new_n426), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n279), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(new_n469), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT88), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n360), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n325), .A2(new_n326), .A3(new_n209), .A4(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n274), .A2(new_n568), .A3(new_n209), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(G20), .B2(new_n246), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n519), .A2(G20), .ZN(new_n574));
  AND2_X1   g0374(.A1(KEYINPUT86), .A2(KEYINPUT24), .ZN(new_n575));
  NOR4_X1   g0375(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(KEYINPUT86), .A2(KEYINPUT24), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n570), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(new_n570), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n257), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n254), .B2(G107), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n254), .A2(new_n581), .A3(G107), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n582), .A2(new_n584), .B1(new_n495), .B2(G107), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n563), .A2(new_n360), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT88), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n563), .A2(G190), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n565), .B(new_n587), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n563), .A2(new_n300), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n553), .A2(new_n556), .B1(new_n561), .B2(new_n279), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n355), .A3(new_n469), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n586), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n552), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n439), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT89), .ZN(G372));
  AND2_X1   g0399(.A1(new_n359), .A2(new_n373), .ZN(new_n600));
  INV_X1    g0400(.A(new_n408), .ZN(new_n601));
  INV_X1    g0401(.A(new_n434), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n411), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n368), .A2(new_n374), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT91), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n299), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n605), .A2(new_n606), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n302), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT92), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n531), .A2(KEYINPUT90), .A3(G200), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT90), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n524), .B2(new_n360), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(new_n614), .A3(new_n548), .A4(new_n549), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n532), .A2(new_n542), .A3(new_n525), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n516), .A2(new_n515), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n616), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n619), .B1(new_n551), .B2(new_n620), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n474), .A2(new_n475), .B1(new_n481), .B2(new_n456), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n595), .A2(new_n625), .A3(new_n473), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n591), .A2(new_n626), .A3(new_n618), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n517), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n439), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n611), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g0431(.A(new_n631), .B(KEYINPUT93), .Z(G369));
  NAND3_X1  g0432(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n587), .A2(new_n639), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n596), .A2(new_n640), .B1(new_n595), .B2(new_n639), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n625), .A2(new_n473), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n456), .A2(new_n638), .ZN(new_n643));
  MUX2_X1   g0443(.A(new_n642), .B(new_n483), .S(new_n643), .Z(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n644), .A3(G330), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n639), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n596), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n645), .B(new_n648), .C1(new_n595), .C2(new_n638), .ZN(G399));
  INV_X1    g0449(.A(new_n212), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n467), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G1), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n536), .A2(new_n442), .A3(new_n537), .ZN(new_n654));
  OAI22_X1  g0454(.A1(new_n653), .A2(new_n654), .B1(new_n218), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n516), .A2(new_n515), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT26), .B1(new_n617), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n620), .A2(new_n619), .A3(new_n550), .A4(new_n543), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n616), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n514), .A2(KEYINPUT82), .A3(G190), .ZN(new_n661));
  INV_X1    g0461(.A(new_n497), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n513), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n663), .A2(KEYINPUT95), .A3(new_n657), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT95), .B1(new_n663), .B2(new_n657), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n660), .B1(new_n666), .B2(new_n627), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT96), .B1(new_n667), .B2(new_n638), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n658), .A2(new_n659), .A3(new_n616), .ZN(new_n669));
  INV_X1    g0469(.A(new_n665), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n517), .A2(KEYINPUT95), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n591), .A2(new_n626), .A3(new_n618), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT96), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n639), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n638), .B1(new_n624), .B2(new_n628), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g0479(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n680));
  AOI22_X1  g0480(.A1(new_n677), .A2(KEYINPUT29), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n597), .A2(new_n639), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT31), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n508), .A2(new_n531), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(new_n593), .A3(new_n481), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n685), .A2(KEYINPUT30), .A3(new_n481), .A4(new_n593), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n472), .A2(new_n355), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n563), .A3(new_n508), .A4(new_n531), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n684), .B1(new_n692), .B2(new_n638), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n684), .A3(new_n638), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n682), .B1(new_n683), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n681), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n656), .B1(new_n698), .B2(G1), .ZN(G364));
  AND2_X1   g0499(.A1(new_n209), .A2(G13), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n208), .B1(new_n700), .B2(G45), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n651), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n220), .B1(G20), .B2(new_n300), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR4_X1   g0506(.A1(new_n209), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT98), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT98), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR4_X1   g0511(.A1(new_n209), .A2(new_n360), .A3(G179), .A4(G190), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n711), .A2(G329), .B1(G283), .B2(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT100), .Z(new_n714));
  NOR2_X1   g0514(.A1(new_n209), .A2(new_n355), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n716), .A2(new_n295), .A3(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n295), .A2(new_n360), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(G20), .A3(new_n355), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n717), .A2(G322), .B1(new_n720), .B2(G303), .ZN(new_n721));
  INV_X1    g0521(.A(G311), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n716), .A2(G190), .A3(G200), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n716), .A2(new_n360), .A3(G190), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  XOR2_X1   g0526(.A(KEYINPUT33), .B(G317), .Z(new_n727));
  OAI221_X1 g0527(.A(new_n721), .B1(new_n722), .B2(new_n724), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n718), .A2(new_n715), .ZN(new_n729));
  INV_X1    g0529(.A(G326), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n209), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n327), .B1(new_n729), .B2(new_n730), .C1(new_n732), .C2(new_n559), .ZN(new_n733));
  OR3_X1    g0533(.A1(new_n714), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n717), .ZN(new_n735));
  INV_X1    g0535(.A(new_n712), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n735), .A2(new_n215), .B1(new_n246), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n729), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n327), .B(new_n737), .C1(G50), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n710), .A2(new_n311), .ZN(new_n740));
  XOR2_X1   g0540(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n741));
  XNOR2_X1  g0541(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n726), .A2(new_n216), .B1(new_n724), .B2(new_n413), .ZN(new_n743));
  INV_X1    g0543(.A(new_n536), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(new_n720), .ZN(new_n745));
  INV_X1    g0545(.A(new_n732), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G97), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n739), .A2(new_n742), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n706), .B1(new_n734), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n705), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n650), .A2(new_n327), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n754), .A2(G355), .B1(new_n442), .B2(new_n650), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT97), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n650), .A2(new_n274), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n219), .A2(new_n282), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n759), .B(new_n760), .C1(new_n245), .C2(new_n282), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n704), .B(new_n749), .C1(new_n753), .C2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n752), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n644), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n644), .A2(G330), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n644), .A2(G330), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n704), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n765), .B1(new_n766), .B2(new_n768), .ZN(G396));
  NAND2_X1  g0569(.A1(new_n434), .A2(KEYINPUT101), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT101), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n425), .A2(new_n432), .A3(new_n771), .A4(new_n433), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(new_n437), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n678), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n425), .A2(new_n638), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n770), .A2(new_n437), .A3(new_n776), .A4(new_n772), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n434), .B2(new_n639), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n775), .B1(new_n678), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n697), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n703), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n780), .B2(new_n779), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n706), .A2(new_n751), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n703), .B1(G77), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G283), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n785), .A2(new_n726), .B1(new_n735), .B2(new_n559), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G116), .B2(new_n723), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n736), .A2(new_n349), .B1(new_n719), .B2(new_n246), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n274), .B(new_n788), .C1(G303), .C2(new_n738), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n711), .A2(G311), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n787), .A2(new_n747), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n725), .A2(G150), .B1(new_n738), .B2(G137), .ZN(new_n792));
  INV_X1    g0592(.A(G143), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n792), .B1(new_n793), .B2(new_n735), .C1(new_n311), .C2(new_n724), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT34), .Z(new_n795));
  NOR2_X1   g0595(.A1(new_n736), .A2(new_n216), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n327), .B(new_n796), .C1(G50), .C2(new_n720), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n797), .B1(new_n215), .B2(new_n732), .C1(new_n798), .C2(new_n710), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n791), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n784), .B1(new_n800), .B2(new_n705), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n778), .B2(new_n751), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n782), .A2(new_n802), .ZN(G384));
  INV_X1    g0603(.A(new_n490), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT35), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT35), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n805), .A2(G116), .A3(new_n221), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT36), .Z(new_n808));
  NAND3_X1  g0608(.A1(new_n219), .A2(G77), .A3(new_n308), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n201), .A2(G68), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n208), .B(G13), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT38), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n366), .B1(new_n372), .B2(new_n357), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n371), .A2(new_n343), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n636), .B1(new_n815), .B2(new_n307), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT37), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n345), .A2(new_n358), .ZN(new_n818));
  INV_X1    g0618(.A(new_n636), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n345), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT37), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n818), .A2(new_n820), .A3(new_n821), .A4(new_n366), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n817), .A2(KEYINPUT103), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n375), .A2(new_n816), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT103), .B1(new_n817), .B2(new_n822), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n813), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n333), .B1(KEYINPUT16), .B2(new_n332), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n307), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n819), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n375), .A2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n306), .B(new_n364), .C1(new_n371), .C2(new_n343), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n828), .A2(new_n307), .B1(new_n357), .B2(new_n636), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT37), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n822), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n832), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT39), .B1(new_n827), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n366), .A2(new_n367), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT17), .B1(new_n372), .B2(new_n365), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n830), .B1(new_n600), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n834), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n821), .B1(new_n843), .B2(new_n366), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n372), .A2(new_n357), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n845), .A2(new_n816), .A3(new_n833), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n846), .B2(new_n821), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n813), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n848), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n838), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n601), .A2(new_n639), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n600), .A2(new_n819), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n773), .A2(new_n638), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n678), .B2(new_n774), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n386), .A2(new_n638), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT102), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n408), .A2(new_n411), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n405), .A2(new_n407), .A3(new_n857), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n857), .A2(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n848), .A2(new_n837), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n854), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n853), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n681), .A2(new_n439), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n611), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n867), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n827), .A2(new_n837), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n683), .A2(new_n696), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n872), .A2(KEYINPUT40), .A3(new_n778), .A4(new_n862), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n692), .A2(new_n684), .A3(new_n638), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(new_n693), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n552), .A2(new_n596), .A3(new_n638), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n778), .B(new_n862), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n848), .B2(new_n837), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n875), .B1(KEYINPUT40), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n439), .A2(new_n872), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(G330), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n870), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n208), .B2(new_n700), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n870), .A2(new_n885), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n812), .B1(new_n887), .B2(new_n888), .ZN(G367));
  NAND2_X1  g0689(.A1(new_n759), .A2(new_n241), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(new_n753), .C1(new_n212), .C2(new_n418), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT106), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n893), .A2(new_n894), .A3(new_n704), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n548), .A2(new_n639), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n618), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n616), .B2(new_n896), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n717), .A2(G150), .B1(G77), .B2(new_n712), .ZN(new_n899));
  INV_X1    g0699(.A(G137), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n899), .B1(new_n215), .B2(new_n719), .C1(new_n710), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n732), .A2(new_n216), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n274), .B1(new_n729), .B2(new_n793), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n311), .A2(new_n726), .B1(new_n724), .B2(new_n201), .ZN(new_n904));
  NOR4_X1   g0704(.A1(new_n901), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT108), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT107), .B1(new_n720), .B2(G116), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT46), .Z(new_n908));
  OAI22_X1  g0708(.A1(new_n726), .A2(new_n559), .B1(new_n724), .B2(new_n785), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n735), .A2(new_n459), .B1(new_n729), .B2(new_n722), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n327), .B1(new_n732), .B2(new_n246), .C1(new_n736), .C2(new_n248), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(G317), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n913), .B2(new_n710), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n906), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT47), .Z(new_n916));
  OAI221_X1 g0716(.A(new_n895), .B1(new_n764), .B2(new_n898), .C1(new_n916), .C2(new_n706), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n672), .B1(new_n497), .B2(new_n638), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n620), .B2(new_n638), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n648), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT42), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n595), .B(new_n672), .C1(new_n497), .C2(new_n638), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n639), .B1(new_n922), .B2(new_n620), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT104), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT105), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n919), .A2(new_n645), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n648), .B1(new_n595), .B2(new_n638), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n919), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT44), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n919), .A2(new_n934), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(new_n645), .ZN(new_n940));
  INV_X1    g0740(.A(new_n646), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n648), .B1(new_n641), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(new_n767), .Z(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n698), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n698), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n651), .B(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n702), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n917), .B1(new_n933), .B2(new_n947), .ZN(G387));
  NAND2_X1  g0748(.A1(new_n943), .A2(new_n702), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n641), .A2(new_n764), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n724), .A2(new_n216), .B1(new_n413), .B2(new_n719), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n327), .B(new_n951), .C1(G97), .C2(new_n712), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n725), .A2(new_n263), .B1(new_n738), .B2(G159), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n380), .B2(new_n735), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n711), .A2(G150), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n418), .A2(new_n732), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n952), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n274), .B1(new_n712), .B2(G116), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n732), .A2(new_n785), .B1(new_n719), .B2(new_n559), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n725), .A2(G311), .B1(new_n738), .B2(G322), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n961), .B1(new_n459), .B2(new_n724), .C1(new_n913), .C2(new_n735), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT48), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n963), .B2(new_n962), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT49), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n959), .B1(new_n730), .B2(new_n710), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n958), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n705), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n263), .A2(new_n380), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT50), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n282), .B1(new_n216), .B2(new_n413), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n972), .A2(new_n654), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n759), .B1(new_n238), .B2(new_n282), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n754), .A2(new_n654), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n212), .A2(G107), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n753), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n970), .A2(new_n703), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n698), .A2(new_n943), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n651), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n698), .A2(new_n943), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n949), .B1(new_n950), .B2(new_n980), .C1(new_n982), .C2(new_n983), .ZN(G393));
  NAND2_X1  g0784(.A1(new_n919), .A2(new_n752), .ZN(new_n985));
  INV_X1    g0785(.A(new_n759), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n753), .B1(new_n248), .B2(new_n212), .C1(new_n986), .C2(new_n252), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n703), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT109), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n327), .B1(new_n732), .B2(new_n442), .C1(new_n736), .C2(new_n246), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n726), .A2(new_n459), .B1(new_n724), .B2(new_n559), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G283), .C2(new_n720), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n711), .A2(G322), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n717), .A2(G311), .B1(new_n738), .B2(G317), .ZN(new_n994));
  XNOR2_X1  g0794(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n717), .A2(G159), .B1(new_n738), .B2(G150), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT51), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n726), .A2(new_n201), .B1(new_n724), .B2(new_n262), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G68), .B2(new_n720), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n711), .A2(G143), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n732), .A2(new_n413), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n327), .B(new_n1003), .C1(G87), .C2(new_n712), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n997), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n989), .B1(new_n1006), .B2(new_n705), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n940), .A2(new_n702), .B1(new_n985), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n944), .A2(new_n651), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n940), .B1(new_n698), .B2(new_n943), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(G390));
  INV_X1    g0811(.A(new_n778), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n668), .B2(new_n676), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n862), .B1(new_n1013), .B2(new_n855), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n852), .B1(new_n827), .B2(new_n837), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT111), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(new_n1015), .A3(KEYINPUT111), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n838), .A2(new_n849), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n851), .B1(new_n856), .B2(new_n863), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1018), .A2(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n697), .A2(new_n778), .A3(new_n862), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT112), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1021), .B1(new_n838), .B2(new_n849), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1019), .ZN(new_n1026));
  AOI21_X1  g0826(.A(KEYINPUT111), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT112), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1023), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1023), .B(new_n1025), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT113), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT113), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1034), .A2(new_n1035), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1024), .A2(new_n1031), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n439), .A2(new_n697), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n611), .A2(new_n868), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n862), .B1(new_n697), .B2(new_n778), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1030), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1013), .A2(new_n855), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n856), .B2(new_n1042), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1037), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n651), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1037), .A2(new_n702), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT114), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT114), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1037), .A2(new_n1055), .A3(new_n702), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n703), .B1(new_n263), .B2(new_n783), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n724), .A2(new_n248), .B1(new_n349), .B2(new_n719), .ZN(new_n1059));
  OR4_X1    g0859(.A1(new_n274), .A2(new_n1059), .A3(new_n796), .A4(new_n1003), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G107), .A2(new_n725), .B1(new_n717), .B2(G116), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n785), .B2(new_n729), .C1(new_n710), .C2(new_n559), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT54), .B(G143), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1064), .A2(new_n723), .B1(new_n725), .B2(G137), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n201), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G128), .A2(new_n738), .B1(new_n1066), .B2(new_n712), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n746), .A2(G159), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n327), .B1(new_n717), .B2(G132), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G150), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n719), .A2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1073));
  XNOR2_X1  g0873(.A(new_n1072), .B(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(G125), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n710), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1060), .A2(new_n1062), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1058), .B1(new_n1077), .B2(new_n705), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n850), .B2(new_n751), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1052), .A2(new_n1057), .A3(new_n1079), .ZN(G378));
  INV_X1    g0880(.A(KEYINPUT57), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT118), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n270), .A2(new_n819), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n299), .B2(new_n302), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n299), .A2(new_n302), .A3(new_n1083), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(G330), .B1(new_n880), .B2(KEYINPUT40), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n873), .B1(new_n827), .B2(new_n837), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1091), .A2(KEYINPUT117), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT117), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n858), .A2(new_n857), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n860), .A2(new_n861), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n778), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n683), .B2(new_n696), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n832), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT38), .B1(new_n832), .B2(new_n836), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT40), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n682), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1094), .B1(new_n875), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1090), .B1(new_n1093), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT117), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1082), .B1(new_n1109), .B2(new_n867), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT119), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1109), .B2(new_n867), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n875), .A2(new_n1103), .A3(new_n1094), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1107), .B1(new_n1106), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n875), .A2(new_n1103), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1090), .B1(new_n1115), .B2(KEYINPUT117), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1111), .B(new_n867), .C1(new_n1114), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n867), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n867), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT119), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1122), .A2(new_n1124), .A3(new_n1117), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1039), .B1(new_n1037), .B2(new_n1047), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1081), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT120), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT120), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1130), .B(new_n1081), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1051), .A2(new_n1040), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1081), .B1(new_n1133), .B2(new_n1123), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n652), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n703), .B1(new_n1066), .B2(new_n783), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n467), .A2(new_n274), .ZN(new_n1138));
  AOI211_X1 g0938(.A(G50), .B(new_n1138), .C1(new_n264), .C2(new_n288), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n248), .A2(new_n726), .B1(new_n735), .B2(new_n246), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n413), .B2(new_n719), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n736), .A2(new_n215), .B1(new_n442), .B2(new_n729), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n902), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n785), .B2(new_n710), .C1(new_n418), .C2(new_n724), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT58), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n711), .A2(G124), .ZN(new_n1147));
  AOI211_X1 g0947(.A(G33), .B(G41), .C1(new_n712), .C2(G159), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n720), .A2(new_n1064), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT116), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n735), .A2(new_n1151), .B1(new_n724), .B2(new_n900), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n726), .A2(new_n798), .B1(new_n729), .B2(new_n1075), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n732), .A2(new_n1071), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT59), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1147), .B(new_n1148), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1155), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1146), .B1(new_n1145), .B2(new_n1144), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1137), .B1(new_n1160), .B2(new_n705), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1107), .B2(new_n751), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n702), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1136), .A2(new_n1165), .ZN(G375));
  AOI22_X1  g0966(.A1(G107), .A2(new_n723), .B1(new_n725), .B2(G116), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(KEYINPUT121), .A2(new_n1167), .B1(new_n711), .B2(G303), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1168), .B(new_n957), .C1(KEYINPUT121), .C2(new_n1167), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n720), .A2(G97), .B1(new_n738), .B2(G294), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n274), .B1(new_n712), .B2(G77), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n785), .C2(new_n735), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n717), .A2(G137), .B1(new_n720), .B2(G159), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n327), .B1(new_n712), .B2(G58), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n380), .C2(new_n732), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n723), .A2(G150), .B1(new_n738), .B2(G132), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n726), .B2(new_n1063), .C1(new_n1151), .C2(new_n710), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1169), .A2(new_n1172), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n705), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1179), .B(new_n703), .C1(G68), .C2(new_n783), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n863), .B2(new_n750), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1045), .B2(new_n702), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1046), .A2(new_n946), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(G381));
  INV_X1    g0985(.A(G378), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1136), .A2(new_n1186), .A3(new_n1165), .ZN(new_n1187));
  OR4_X1    g0987(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1188));
  OR4_X1    g0988(.A1(G387), .A2(new_n1187), .A3(G381), .A4(new_n1188), .ZN(G407));
  OAI211_X1 g0989(.A(G407), .B(G213), .C1(G343), .C2(new_n1187), .ZN(G409));
  XNOR2_X1  g0990(.A(G393), .B(G396), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(G390), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(G387), .B(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n637), .A2(G213), .ZN(new_n1195));
  INV_X1    g0995(.A(G384), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT125), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1046), .A2(KEYINPUT60), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1184), .A2(KEYINPUT60), .A3(new_n1046), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n651), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1197), .B1(new_n1201), .B2(new_n1182), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1196), .A2(KEYINPUT125), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1136), .A2(G378), .A3(new_n1165), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1132), .A2(new_n946), .A3(new_n1125), .A4(new_n1119), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT122), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1133), .A2(new_n1123), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT123), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n701), .B1(new_n1210), .B2(KEYINPUT123), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1163), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT122), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1164), .A2(new_n1214), .A3(new_n946), .A4(new_n1132), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1209), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT124), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1186), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1207), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1217), .B1(new_n1216), .B2(new_n1186), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1195), .B(new_n1206), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1220), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n1218), .A3(new_n1207), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1225), .A2(KEYINPUT126), .A3(new_n1195), .A4(new_n1206), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT62), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1195), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n637), .A2(G213), .A3(G2897), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1206), .B(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT61), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1221), .A2(KEYINPUT62), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1194), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT63), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1223), .A2(new_n1226), .A3(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1221), .A2(new_n1235), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n1231), .A3(new_n1193), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(G405));
  INV_X1    g1039(.A(KEYINPUT127), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1207), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G378), .B1(new_n1136), .B2(new_n1165), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1242), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(KEYINPUT127), .A3(new_n1207), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(new_n1245), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(KEYINPUT127), .A3(new_n1207), .A4(new_n1206), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(new_n1193), .ZN(G402));
endmodule


