//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT93), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT93), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT15), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT96), .ZN(new_n207));
  INV_X1    g006(.A(G43gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(G50gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n206), .B(new_n209), .C1(new_n202), .C2(new_n207), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT94), .B(G36gat), .Z(new_n212));
  AND2_X1   g011(.A1(new_n212), .A2(G29gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT95), .ZN(new_n214));
  NOR2_X1   g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n215), .B(KEYINPUT14), .Z(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(KEYINPUT95), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n205), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G1gat), .B2(new_n223), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(G8gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n219), .A2(new_n229), .A3(new_n220), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n222), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n219), .A2(new_n220), .A3(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n228), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n237), .A2(new_n232), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n233), .B(KEYINPUT13), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n232), .A4(new_n233), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT11), .B(G169gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(G197gat), .ZN(new_n244));
  XOR2_X1   g043(.A(G113gat), .B(G141gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT12), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n236), .A2(new_n240), .A3(new_n247), .A4(new_n241), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G190gat), .ZN(new_n253));
  AND2_X1   g052(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT28), .ZN(new_n257));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT26), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n265), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n257), .A2(new_n258), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT68), .ZN(new_n268));
  INV_X1    g067(.A(new_n258), .ZN(new_n269));
  INV_X1    g068(.A(new_n262), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n270), .B1(new_n260), .B2(new_n259), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n269), .B1(new_n271), .B2(new_n263), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n257), .A4(new_n266), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT23), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n259), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n275), .A2(G169gat), .A3(G176gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n258), .A2(KEYINPUT24), .ZN(new_n282));
  NOR2_X1   g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n269), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n284), .B2(KEYINPUT24), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT25), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n270), .B2(KEYINPUT67), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n281), .A2(new_n285), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n259), .A2(KEYINPUT23), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n262), .B(new_n291), .C1(new_n292), .C2(new_n259), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n253), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT24), .A3(new_n258), .ZN(new_n296));
  INV_X1    g095(.A(new_n282), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n290), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n268), .A2(new_n274), .B1(new_n289), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G113gat), .ZN(new_n302));
  INV_X1    g101(.A(G113gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G120gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G127gat), .B(G134gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G127gat), .B(G134gat), .Z(new_n312));
  OAI211_X1 g111(.A(new_n306), .B(new_n305), .C1(new_n312), .C2(new_n308), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT70), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n315));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n310), .B1(new_n316), .B2(KEYINPUT69), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(KEYINPUT1), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI221_X4 g118(.A(KEYINPUT1), .B1(new_n302), .B2(new_n304), .C1(new_n310), .C2(KEYINPUT69), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n300), .A2(new_n314), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n289), .A2(new_n299), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT27), .B(G183gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n265), .B1(new_n324), .B2(new_n253), .ZN(new_n325));
  INV_X1    g124(.A(new_n266), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n273), .B1(new_n327), .B2(new_n272), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n257), .A2(new_n266), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n264), .A2(new_n258), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT68), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n323), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n321), .A2(new_n314), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n322), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT34), .ZN(new_n336));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT64), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n335), .B2(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n338), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n334), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT32), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n346), .B2(KEYINPUT32), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G15gat), .B(G43gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(G71gat), .ZN(new_n355));
  INV_X1    g154(.A(G99gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n350), .A2(new_n351), .A3(new_n353), .A4(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n353), .B(new_n357), .C1(new_n348), .C2(new_n349), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT72), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(KEYINPUT33), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n346), .A2(KEYINPUT32), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n344), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n358), .B2(new_n360), .ZN(new_n365));
  INV_X1    g164(.A(new_n344), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(KEYINPUT36), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT36), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n365), .A2(new_n366), .ZN(new_n370));
  AOI211_X1 g169(.A(new_n363), .B(new_n344), .C1(new_n358), .C2(new_n360), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT0), .B(G57gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(G85gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G155gat), .B(G162gat), .ZN(new_n379));
  XOR2_X1   g178(.A(G141gat), .B(G148gat), .Z(new_n380));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G141gat), .B(G148gat), .ZN(new_n383));
  INV_X1    g182(.A(G162gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT81), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G162gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n387), .A3(G155gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n383), .B1(new_n388), .B2(KEYINPUT2), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n382), .B1(new_n379), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n311), .A2(new_n313), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT84), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n394), .A3(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n391), .B2(new_n390), .ZN(new_n397));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n389), .A2(new_n379), .ZN(new_n402));
  INV_X1    g201(.A(new_n382), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(new_n321), .B2(new_n314), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT83), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n393), .A2(new_n406), .A3(new_n395), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT70), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT70), .B1(new_n311), .B2(new_n313), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n390), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT4), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n404), .A2(KEYINPUT3), .ZN(new_n415));
  XOR2_X1   g214(.A(KEYINPUT82), .B(KEYINPUT3), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n390), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n415), .A2(new_n418), .A3(new_n313), .A4(new_n311), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n419), .A2(new_n398), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n414), .A2(KEYINPUT85), .A3(new_n420), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n401), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n411), .A2(new_n406), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(new_n419), .C1(new_n396), .C2(new_n406), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n427), .A2(KEYINPUT5), .A3(new_n399), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n378), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n414), .A2(KEYINPUT85), .A3(new_n420), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT85), .B1(new_n414), .B2(new_n420), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n428), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n377), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT6), .B(new_n378), .C1(new_n425), .C2(new_n428), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n440));
  NAND2_X1  g239(.A1(G226gat), .A2(G233gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n290), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n279), .A2(new_n270), .A3(new_n280), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n285), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n288), .B(new_n291), .C1(new_n292), .C2(new_n259), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n286), .A2(new_n296), .A3(new_n297), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n267), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n442), .A2(KEYINPUT29), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n300), .A2(new_n442), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT77), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT75), .B(G218gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G211gat), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT22), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT74), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT22), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G197gat), .B(G204gat), .Z(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(G211gat), .A2(G218gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(G211gat), .A2(G218gat), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT76), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G211gat), .ZN(new_n467));
  INV_X1    g266(.A(G218gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT76), .ZN(new_n470));
  NAND2_X1  g269(.A1(G211gat), .A2(G218gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n461), .A2(new_n463), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n459), .B1(G211gat), .B2(new_n453), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n466), .A2(new_n472), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n474), .A2(new_n475), .A3(new_n462), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n452), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n461), .A2(new_n466), .A3(new_n472), .A4(new_n463), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n474), .B2(new_n462), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT77), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n440), .B1(new_n451), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n289), .A2(new_n299), .B1(new_n272), .B2(new_n327), .ZN(new_n483));
  INV_X1    g282(.A(new_n450), .ZN(new_n484));
  OAI22_X1  g283(.A1(new_n332), .A2(new_n441), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n477), .A2(new_n480), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(KEYINPUT80), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT78), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n441), .C1(new_n300), .C2(KEYINPUT29), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT29), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n442), .B1(new_n332), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT78), .B1(new_n483), .B2(new_n441), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n481), .B(new_n490), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT79), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n441), .B1(new_n300), .B2(KEYINPUT29), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n489), .B1(new_n449), .B2(new_n442), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT79), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n481), .A4(new_n490), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n488), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G8gat), .B(G36gat), .ZN(new_n502));
  INV_X1    g301(.A(G64gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G92gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n501), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n506), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n507), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n439), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT29), .B1(new_n390), .B2(new_n417), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n480), .B2(new_n477), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n404), .A2(new_n491), .A3(new_n478), .A4(new_n479), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(G228gat), .A3(G233gat), .A4(new_n415), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n404), .A2(new_n416), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n486), .B2(new_n517), .ZN(new_n525));
  NAND2_X1  g324(.A1(G228gat), .A2(G233gat), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT87), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n519), .A2(new_n523), .ZN(new_n528));
  OAI211_X1 g327(.A(KEYINPUT87), .B(new_n526), .C1(new_n518), .C2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n522), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G22gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n526), .B1(new_n518), .B2(new_n528), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n521), .B1(new_n535), .B2(new_n529), .ZN(new_n536));
  INV_X1    g335(.A(G22gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n532), .A2(KEYINPUT88), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  XOR2_X1   g340(.A(G78gat), .B(G106gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT31), .ZN(new_n543));
  INV_X1    g342(.A(G50gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT86), .Z(new_n546));
  NAND3_X1  g345(.A1(new_n539), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n538), .A3(new_n545), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n516), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n373), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT89), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT91), .B(KEYINPUT37), .Z(new_n554));
  AOI211_X1 g353(.A(new_n554), .B(new_n488), .C1(new_n495), .C2(new_n500), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT37), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n495), .A2(new_n500), .ZN(new_n557));
  INV_X1    g356(.A(new_n488), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT38), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n554), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT38), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n498), .A2(new_n486), .A3(new_n490), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(KEYINPUT37), .C1(new_n486), .C2(new_n451), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(new_n506), .A3(new_n566), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n501), .A2(KEYINPUT38), .A3(new_n506), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n439), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(KEYINPUT90), .A2(KEYINPUT40), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n427), .A2(new_n399), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n396), .B(new_n398), .C1(new_n391), .C2(new_n390), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n572), .A2(KEYINPUT39), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT39), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n427), .A2(new_n575), .A3(new_n399), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n377), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n571), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n572), .A2(KEYINPUT39), .A3(new_n573), .ZN(new_n579));
  INV_X1    g378(.A(new_n571), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n579), .A2(new_n377), .A3(new_n580), .A4(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n377), .B1(new_n434), .B2(new_n435), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n514), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n549), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT92), .B1(new_n570), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n514), .A2(new_n584), .B1(new_n547), .B2(new_n548), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n562), .B1(new_n556), .B2(new_n501), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n507), .B1(new_n590), .B2(KEYINPUT38), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n568), .B1(new_n591), .B2(new_n566), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n588), .B(new_n589), .C1(new_n592), .C2(new_n439), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n368), .A2(new_n372), .B1(new_n550), .B2(new_n516), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n553), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n370), .A2(new_n371), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n549), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n599), .B1(new_n601), .B2(new_n516), .ZN(new_n602));
  INV_X1    g401(.A(new_n516), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n603), .A2(KEYINPUT35), .A3(new_n600), .A4(new_n549), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n252), .B1(new_n598), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT97), .B(G57gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G64gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n503), .A2(G57gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(G71gat), .ZN(new_n612));
  INV_X1    g411(.A(G78gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(G71gat), .A2(G78gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT9), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G57gat), .B(G64gat), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT9), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n614), .A2(new_n616), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n611), .A2(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n620), .A2(new_n621), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n609), .A2(new_n610), .B1(new_n615), .B2(new_n617), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT98), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n227), .B1(new_n628), .B2(KEYINPUT21), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n294), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n624), .A2(new_n627), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT99), .B(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G211gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n634), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT102), .B(KEYINPUT7), .ZN(new_n644));
  NAND2_X1  g443(.A1(G85gat), .A2(G92gat), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G99gat), .A2(G106gat), .ZN(new_n647));
  INV_X1    g446(.A(G85gat), .ZN(new_n648));
  AOI22_X1  g447(.A1(KEYINPUT8), .A2(new_n647), .B1(new_n648), .B2(new_n505), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G99gat), .B(G106gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  NAND3_X1  g452(.A1(new_n222), .A2(new_n230), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n651), .B(new_n652), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n219), .A2(new_n220), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G134gat), .B(G162gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G190gat), .B(G218gat), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n660), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n643), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G230gat), .A2(G233gat), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n628), .B2(new_n656), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n635), .A2(new_n653), .A3(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n656), .A2(new_n622), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT104), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n656), .A2(new_n673), .A3(new_n622), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n669), .A2(new_n670), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n628), .A2(new_n656), .A3(KEYINPUT10), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n667), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n675), .A2(new_n666), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(G120gat), .B(G148gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G176gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(G204gat), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n679), .B2(new_n680), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n665), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n607), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n437), .A2(new_n438), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g493(.A1(new_n690), .A2(new_n515), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(KEYINPUT105), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(KEYINPUT105), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(G8gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT16), .B(G8gat), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n695), .A2(KEYINPUT42), .A3(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n699), .B(new_n702), .C1(KEYINPUT42), .C2(new_n701), .ZN(G1325gat));
  INV_X1    g502(.A(new_n373), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n691), .A2(G15gat), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(G15gat), .B1(new_n691), .B2(new_n600), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n690), .A2(new_n549), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT106), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n708), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(new_n643), .ZN(new_n712));
  INV_X1    g511(.A(new_n688), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n664), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n607), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(G29gat), .A3(new_n439), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT45), .Z(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n719), .B(new_n664), .C1(new_n598), .C2(new_n606), .ZN(new_n720));
  INV_X1    g519(.A(new_n593), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n567), .A2(new_n569), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n692), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n589), .B1(new_n723), .B2(new_n588), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT108), .B(new_n595), .C1(new_n721), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT108), .B1(new_n594), .B2(new_n595), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n606), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n663), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n660), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n720), .B1(new_n719), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n251), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n249), .A2(KEYINPUT107), .A3(new_n250), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n714), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n732), .A2(new_n692), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G29gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n718), .A2(new_n740), .ZN(G1328gat));
  NOR2_X1   g540(.A1(new_n515), .A2(new_n212), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n607), .A2(new_n715), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT46), .Z(new_n744));
  NAND2_X1  g543(.A1(new_n594), .A2(new_n595), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n605), .B1(new_n747), .B2(new_n725), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n719), .B1(new_n748), .B2(new_n664), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n598), .A2(new_n606), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(KEYINPUT44), .A3(new_n730), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n749), .A2(new_n514), .A3(new_n738), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n212), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n744), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT109), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n744), .A2(new_n756), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1329gat));
  INV_X1    g557(.A(new_n600), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n208), .B1(new_n716), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n749), .A2(G43gat), .A3(new_n738), .A4(new_n751), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n760), .B(new_n762), .C1(new_n763), .C2(new_n373), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1330gat));
  NAND4_X1  g565(.A1(new_n732), .A2(G50gat), .A3(new_n550), .A4(new_n738), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n544), .B1(new_n716), .B2(new_n549), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n767), .A2(KEYINPUT48), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT48), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(G1331gat));
  INV_X1    g570(.A(new_n665), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n736), .A2(new_n713), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n728), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n439), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(new_n608), .ZN(G1332gat));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n774), .A2(new_n777), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n515), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT49), .B(G64gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n782), .B2(new_n785), .ZN(G1333gat));
  OAI211_X1 g585(.A(G71gat), .B(new_n704), .C1(new_n778), .C2(new_n780), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n612), .B1(new_n774), .B2(new_n759), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT50), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n791), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1334gat));
  OAI21_X1  g592(.A(new_n550), .B1(new_n778), .B2(new_n780), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g594(.A1(new_n737), .A2(new_n712), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT112), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n688), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n749), .A2(new_n751), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(G85gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n728), .A2(new_n730), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT51), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n728), .A2(new_n803), .A3(new_n730), .A4(new_n797), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n692), .A3(new_n688), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n692), .A2(new_n800), .B1(new_n806), .B2(new_n648), .ZN(G1336gat));
  NAND4_X1  g606(.A1(new_n749), .A2(new_n514), .A3(new_n751), .A4(new_n798), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G92gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT113), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n515), .A2(G92gat), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n802), .A2(new_n688), .A3(new_n804), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n813), .A3(KEYINPUT52), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n809), .B(new_n812), .C1(KEYINPUT113), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1337gat));
  NAND3_X1  g616(.A1(new_n732), .A2(new_n704), .A3(new_n798), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT114), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n799), .A2(new_n820), .A3(new_n704), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n821), .A3(G99gat), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n805), .A2(new_n356), .A3(new_n600), .A4(new_n688), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1338gat));
  NAND4_X1  g623(.A1(new_n802), .A2(new_n550), .A3(new_n688), .A4(new_n804), .ZN(new_n825));
  INV_X1    g624(.A(G106gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n732), .A2(G106gat), .A3(new_n550), .A4(new_n798), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1339gat));
  NOR3_X1   g632(.A1(new_n665), .A2(new_n688), .A3(new_n736), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n677), .A2(new_n678), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n666), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n677), .A2(new_n667), .A3(new_n678), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n685), .B1(new_n679), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n237), .A2(new_n232), .A3(new_n239), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n237), .A2(KEYINPUT115), .A3(new_n232), .A4(new_n239), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n233), .B1(new_n231), .B2(new_n232), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n246), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n250), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n843), .A2(new_n851), .A3(new_n686), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT116), .B1(new_n853), .B2(new_n664), .ZN(new_n854));
  INV_X1    g653(.A(new_n852), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT55), .B1(new_n838), .B2(new_n840), .ZN(new_n856));
  INV_X1    g655(.A(new_n686), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n730), .A4(new_n851), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n736), .A2(new_n858), .B1(new_n688), .B2(new_n851), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n854), .B(new_n860), .C1(new_n861), .C2(new_n730), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n834), .B1(new_n862), .B2(new_n712), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n601), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n439), .A2(new_n514), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n303), .A3(new_n736), .ZN(new_n868));
  OAI21_X1  g667(.A(G113gat), .B1(new_n866), .B2(new_n252), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1340gat));
  OAI21_X1  g669(.A(G120gat), .B1(new_n866), .B2(new_n713), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(KEYINPUT117), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(KEYINPUT117), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n688), .A2(new_n301), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n874), .B(KEYINPUT118), .Z(new_n875));
  OAI22_X1  g674(.A1(new_n872), .A2(new_n873), .B1(new_n866), .B2(new_n875), .ZN(G1341gat));
  NOR2_X1   g675(.A1(new_n866), .A2(new_n712), .ZN(new_n877));
  XNOR2_X1  g676(.A(KEYINPUT119), .B(G127gat), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n877), .B(new_n878), .ZN(G1342gat));
  NOR3_X1   g678(.A1(new_n866), .A2(G134gat), .A3(new_n664), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT56), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n866), .B2(new_n664), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G1343gat));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n736), .A2(new_n858), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n851), .A2(new_n688), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n730), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n860), .A2(new_n854), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n712), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n834), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n549), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n886), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT120), .B(new_n895), .C1(new_n863), .C2(new_n549), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n843), .A2(new_n251), .A3(new_n686), .A4(new_n852), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n888), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT121), .B1(new_n898), .B2(new_n664), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  AOI211_X1 g699(.A(new_n900), .B(new_n730), .C1(new_n897), .C2(new_n888), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n890), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n643), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT57), .B(new_n550), .C1(new_n904), .C2(new_n834), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n894), .A2(new_n896), .A3(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n373), .A2(new_n865), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n251), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G141gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n907), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(G141gat), .A3(new_n252), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  XOR2_X1   g711(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n906), .A2(new_n736), .A3(new_n907), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n911), .B1(new_n916), .B2(G141gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(G1344gat));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n906), .A2(new_n907), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n919), .B(G148gat), .C1(new_n920), .C2(new_n713), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT57), .B1(new_n863), .B2(new_n549), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n898), .A2(new_n664), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n858), .A2(new_n730), .A3(new_n851), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n643), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n665), .A2(new_n251), .A3(new_n688), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n895), .B(new_n550), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n922), .A2(new_n688), .A3(new_n907), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G148gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT59), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n921), .A2(new_n930), .ZN(new_n931));
  OR3_X1    g730(.A1(new_n910), .A2(G148gat), .A3(new_n713), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1345gat));
  INV_X1    g732(.A(new_n910), .ZN(new_n934));
  AOI21_X1  g733(.A(G155gat), .B1(new_n934), .B2(new_n643), .ZN(new_n935));
  INV_X1    g734(.A(new_n920), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n643), .A2(G155gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G1346gat));
  NAND2_X1  g737(.A1(new_n385), .A2(new_n387), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n920), .A2(new_n939), .A3(new_n664), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n934), .A2(new_n730), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(G1347gat));
  NOR2_X1   g741(.A1(new_n692), .A2(new_n515), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n864), .A2(new_n943), .ZN(new_n944));
  OR3_X1    g743(.A1(new_n944), .A2(G169gat), .A3(new_n737), .ZN(new_n945));
  OAI21_X1  g744(.A(G169gat), .B1(new_n944), .B2(new_n252), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1348gat));
  INV_X1    g746(.A(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n688), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g749(.A1(new_n948), .A2(new_n324), .A3(new_n643), .ZN(new_n951));
  OAI21_X1  g750(.A(G183gat), .B1(new_n944), .B2(new_n712), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(KEYINPUT123), .A3(new_n952), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g753(.A1(new_n948), .A2(new_n730), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G190gat), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(KEYINPUT124), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(KEYINPUT124), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n957), .A2(KEYINPUT124), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n955), .A2(G190gat), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n958), .B(new_n961), .C1(G190gat), .C2(new_n955), .ZN(G1351gat));
  AND2_X1   g761(.A1(new_n373), .A2(new_n943), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n922), .A2(new_n251), .A3(new_n927), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G197gat), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n893), .A2(new_n963), .ZN(new_n966));
  INV_X1    g765(.A(G197gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n967), .A3(new_n736), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT125), .Z(G1352gat));
  XOR2_X1   g769(.A(KEYINPUT126), .B(G204gat), .Z(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n966), .A2(new_n688), .A3(new_n972), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  AND2_X1   g773(.A1(new_n922), .A2(new_n927), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(new_n688), .A3(new_n963), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n974), .B1(new_n972), .B2(new_n976), .ZN(G1353gat));
  NAND3_X1  g776(.A1(new_n966), .A2(new_n467), .A3(new_n643), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n643), .A3(new_n963), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  AOI21_X1  g781(.A(G218gat), .B1(new_n966), .B2(new_n730), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n975), .A2(new_n963), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n730), .A2(new_n453), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n985), .B(KEYINPUT127), .Z(new_n986));
  AOI21_X1  g785(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(G1355gat));
endmodule


