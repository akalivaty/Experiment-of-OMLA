//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT0), .B(G128), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT65), .A2(G134), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(G137), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n200), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n201), .A2(new_n202), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT11), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n207), .A2(new_n210), .A3(G131), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n204), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT65), .A2(G134), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n209), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT11), .B1(new_n216), .B2(new_n205), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n215), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n200), .B1(new_n218), .B2(G137), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n212), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n199), .B1(new_n211), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n205), .B1(new_n218), .B2(G137), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n212), .B(new_n219), .C1(new_n222), .C2(new_n200), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n192), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n195), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n192), .A2(new_n194), .A3(new_n224), .A4(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n189), .A2(new_n230), .A3(new_n224), .A4(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n218), .A2(G137), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n209), .A2(G134), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n223), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n221), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT68), .B(G119), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G116), .ZN(new_n242));
  INV_X1    g056(.A(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT2), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n238), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT68), .A2(G119), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT68), .A2(G119), .ZN(new_n250));
  OAI21_X1  g064(.A(G116), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n240), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n253), .A2(KEYINPUT69), .A3(new_n244), .A4(new_n246), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n242), .A2(new_n257), .A3(new_n247), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(new_n247), .A3(new_n252), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n255), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n256), .B1(new_n255), .B2(new_n261), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n237), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n255), .A2(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n255), .A2(new_n256), .A3(new_n261), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n221), .A4(new_n236), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n187), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT74), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n237), .A2(new_n262), .A3(new_n263), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n266), .A2(new_n267), .B1(new_n221), .B2(new_n236), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT28), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n237), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n262), .A2(new_n263), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT28), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n270), .B1(new_n278), .B2(KEYINPUT74), .ZN(new_n279));
  INV_X1    g093(.A(G237), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G210), .ZN(new_n282));
  INV_X1    g096(.A(G101), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n284), .B(new_n285), .Z(new_n286));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n223), .A2(new_n232), .A3(new_n235), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n190), .A2(new_n198), .ZN(new_n290));
  OAI21_X1  g104(.A(G131), .B1(new_n207), .B2(new_n210), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(new_n223), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n288), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n237), .A2(new_n295), .A3(new_n288), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n221), .A2(KEYINPUT30), .A3(new_n236), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n221), .A2(KEYINPUT72), .A3(KEYINPUT30), .A4(new_n236), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n275), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n297), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n268), .ZN(new_n305));
  INV_X1    g119(.A(new_n286), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT29), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n287), .B2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n273), .A2(new_n277), .A3(KEYINPUT29), .A4(new_n286), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n309), .B(KEYINPUT76), .Z(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G472), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n279), .B2(new_n286), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT74), .B1(new_n269), .B2(new_n276), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n273), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n286), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT75), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT31), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT73), .B1(new_n271), .B2(new_n306), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n268), .A2(new_n323), .A3(new_n286), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n304), .A2(new_n321), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n304), .A2(new_n322), .A3(new_n324), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT31), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n315), .A2(new_n320), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n313), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n327), .B(new_n325), .C1(new_n319), .C2(KEYINPUT75), .ZN(new_n331));
  AOI211_X1 g145(.A(new_n314), .B(new_n286), .C1(new_n316), .C2(new_n318), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n313), .B(new_n329), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n312), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G116), .B(G122), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT14), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G116), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT14), .A3(G122), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(G107), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G107), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT85), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT85), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G107), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n336), .ZN(new_n347));
  XNOR2_X1  g161(.A(G128), .B(G143), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n218), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n218), .A2(new_n348), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n341), .B(new_n347), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT95), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n204), .B1(new_n348), .B2(KEYINPUT13), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n191), .A2(G128), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(KEYINPUT13), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n346), .B(new_n336), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n349), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT9), .B(G234), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT82), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G217), .A3(new_n281), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n359), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G902), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G478), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n365), .B(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G475), .A2(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n280), .A2(new_n281), .A3(G214), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(G143), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT18), .A2(G131), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n372), .B(new_n373), .Z(new_n374));
  XNOR2_X1  g188(.A(G125), .B(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n193), .ZN(new_n376));
  INV_X1    g190(.A(G140), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT79), .B1(new_n377), .B2(G125), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT78), .B(G125), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n377), .ZN(new_n381));
  INV_X1    g195(.A(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT78), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n376), .B1(new_n390), .B2(new_n193), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n374), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n378), .B1(new_n386), .B2(G140), .ZN(new_n393));
  AOI211_X1 g207(.A(KEYINPUT79), .B(new_n377), .C1(new_n383), .C2(new_n385), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT19), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT19), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n375), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n193), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n381), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n400));
  OR3_X1    g214(.A1(new_n386), .A2(KEYINPUT16), .A3(G140), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(G146), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n372), .B(G131), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n399), .B1(new_n398), .B2(new_n402), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n392), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT91), .ZN(new_n409));
  XNOR2_X1  g223(.A(G113), .B(G122), .ZN(new_n410));
  INV_X1    g224(.A(G104), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(new_n392), .C1(new_n406), .C2(new_n407), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n402), .ZN(new_n417));
  AOI21_X1  g231(.A(G146), .B1(new_n400), .B2(new_n401), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n372), .A2(new_n420), .A3(new_n212), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n419), .B(new_n421), .C1(KEYINPUT17), .C2(new_n405), .ZN(new_n422));
  XOR2_X1   g236(.A(new_n412), .B(KEYINPUT92), .Z(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n392), .A3(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n416), .A2(KEYINPUT93), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT93), .B1(new_n416), .B2(new_n424), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT20), .B(new_n370), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n416), .A2(new_n424), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n370), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n424), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT94), .B1(new_n422), .B2(new_n392), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n412), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n422), .A2(KEYINPUT94), .A3(new_n392), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G475), .B1(new_n436), .B2(G902), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n369), .A2(new_n427), .A3(new_n431), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n281), .A2(G952), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(G234), .B2(G237), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G898), .Z(new_n442));
  INV_X1    g256(.A(G234), .ZN(new_n443));
  OAI211_X1 g257(.A(G902), .B(G953), .C1(new_n443), .C2(new_n280), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n241), .A2(new_n448), .A3(G116), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(G113), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n261), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT3), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n344), .A2(G107), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n342), .A2(KEYINPUT85), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n452), .B(G104), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT86), .B(G101), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n342), .A2(G104), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n342), .A2(G104), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(KEYINPUT3), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n343), .A2(new_n345), .A3(new_n411), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G101), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n451), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  XOR2_X1   g280(.A(G110), .B(G122), .Z(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n283), .B1(new_n455), .B2(new_n459), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n460), .A2(KEYINPUT4), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n472), .B2(new_n469), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n466), .B(new_n468), .C1(new_n275), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n449), .A2(G113), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n449), .A2(new_n477), .A3(G113), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n447), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n464), .B1(new_n479), .B2(new_n261), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n467), .B(KEYINPUT8), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n460), .A2(new_n463), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(new_n451), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n232), .A2(new_n386), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n199), .A2(new_n380), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G224), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(G953), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n490), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n486), .B2(new_n487), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n488), .A2(KEYINPUT7), .A3(new_n490), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n485), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n473), .B1(new_n266), .B2(new_n267), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n467), .B1(new_n499), .B2(new_n465), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n474), .A3(KEYINPUT6), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n502), .B(new_n467), .C1(new_n499), .C2(new_n465), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n491), .A2(new_n493), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G210), .B1(G237), .B2(G902), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n498), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n498), .B2(new_n505), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n445), .B(new_n446), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n438), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  INV_X1    g326(.A(G221), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n513), .A2(new_n443), .A3(G953), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n512), .B(new_n514), .Z(new_n515));
  NAND2_X1  g329(.A1(new_n241), .A2(G128), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT23), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n241), .B2(G128), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n249), .A2(new_n250), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT77), .A3(new_n226), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n226), .A2(KEYINPUT23), .A3(G119), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G110), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n516), .B1(new_n239), .B2(G128), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT24), .B(G110), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n525), .B(new_n528), .C1(new_n417), .C2(new_n418), .ZN(new_n529));
  INV_X1    g343(.A(G110), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n522), .A2(new_n530), .A3(new_n523), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n527), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n376), .A3(new_n402), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n529), .A2(new_n534), .A3(KEYINPUT80), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT80), .B1(new_n529), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n515), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n515), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n529), .A2(new_n534), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT80), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(new_n364), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT81), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G217), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(G234), .B2(new_n364), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n542), .A2(new_n544), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n537), .A2(KEYINPUT25), .A3(new_n364), .A4(new_n541), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT81), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n545), .B(new_n547), .C1(new_n548), .C2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n547), .A2(G902), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n537), .A2(new_n541), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G469), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n471), .B(new_n199), .C1(new_n472), .C2(new_n469), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n483), .A2(KEYINPUT10), .A3(new_n232), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n211), .A2(new_n220), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT87), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(new_n464), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT10), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n232), .A2(KEYINPUT87), .A3(new_n460), .A4(new_n463), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n559), .A2(new_n560), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT88), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n559), .A2(KEYINPUT88), .A3(new_n560), .A4(new_n566), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n562), .A2(new_n464), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n563), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n560), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n281), .A2(G227), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G140), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT83), .B(G110), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n571), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n560), .B1(new_n559), .B2(new_n566), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n571), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n556), .B(new_n364), .C1(new_n582), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n571), .A2(new_n577), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n581), .B(KEYINPUT84), .Z(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n581), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n569), .B2(new_n570), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n584), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(G469), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n556), .A2(new_n364), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n586), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n513), .B1(new_n361), .B2(new_n364), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n335), .A2(new_n511), .A3(new_n555), .A4(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(new_n456), .Z(G3));
  NAND3_X1  g417(.A1(new_n427), .A2(new_n431), .A3(new_n437), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n363), .A2(KEYINPUT33), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n363), .A2(KEYINPUT33), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(G478), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(G478), .A2(G902), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n363), .A2(new_n366), .A3(new_n364), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n446), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n509), .B2(KEYINPUT96), .ZN(new_n613));
  INV_X1    g427(.A(new_n506), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n497), .A2(new_n474), .A3(new_n484), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n364), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n614), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n619), .A3(new_n507), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n613), .A2(new_n620), .A3(new_n445), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n611), .A2(new_n621), .A3(KEYINPUT97), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n604), .A2(new_n610), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n613), .A2(new_n620), .A3(new_n445), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n600), .A2(new_n554), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n364), .B1(new_n331), .B2(new_n332), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n629), .A2(G472), .B1(new_n328), .B2(new_n329), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(KEYINPUT93), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n428), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n416), .A2(KEYINPUT93), .A3(new_n424), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT20), .B1(new_n638), .B2(new_n370), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n427), .A2(new_n437), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n368), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n625), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n631), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n538), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n539), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n552), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n551), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n630), .A2(new_n511), .A3(new_n601), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  NAND3_X1  g467(.A1(new_n650), .A2(new_n599), .A3(new_n597), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT32), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n333), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n657), .B2(new_n312), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n613), .A2(new_n620), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n441), .B1(new_n444), .B2(G900), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n642), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n226), .ZN(G30));
  NAND2_X1  g479(.A1(new_n604), .A2(new_n368), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  INV_X1    g481(.A(G472), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n306), .B1(new_n271), .B2(new_n272), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n326), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n668), .B1(new_n670), .B2(new_n364), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n667), .B1(new_n657), .B2(new_n672), .ZN(new_n673));
  AOI211_X1 g487(.A(KEYINPUT99), .B(new_n671), .C1(new_n656), .C2(new_n333), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n661), .B(KEYINPUT39), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n601), .A2(new_n677), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n666), .B(new_n675), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n446), .B1(new_n678), .B2(new_n676), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n650), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n508), .A2(new_n509), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n679), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  NOR2_X1   g502(.A1(new_n624), .A2(new_n662), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n660), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n193), .ZN(G48));
  OAI221_X1 g505(.A(new_n364), .B1(KEYINPUT100), .B2(new_n556), .C1(new_n582), .C2(new_n585), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n556), .A2(KEYINPUT100), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n571), .A2(new_n584), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n694), .A2(new_n591), .B1(new_n592), .B2(new_n577), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n693), .B1(new_n695), .B2(G902), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n692), .A2(new_n696), .A3(new_n599), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n335), .A2(new_n555), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n627), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT41), .B(G113), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT101), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n699), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n643), .A2(new_n335), .A3(new_n555), .A4(new_n697), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  AND3_X1   g518(.A1(new_n659), .A2(new_n697), .A3(new_n445), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n438), .B1(new_n551), .B2(new_n649), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n335), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n668), .B1(new_n308), .B2(new_n310), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n656), .B2(new_n333), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n659), .A2(new_n697), .A3(new_n445), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(KEYINPUT102), .A3(new_n706), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  NAND2_X1  g530(.A1(new_n629), .A2(G472), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n278), .A2(new_n306), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n327), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n325), .B1(new_n719), .B2(KEYINPUT103), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n326), .A2(KEYINPUT31), .B1(new_n278), .B2(new_n306), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n329), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n555), .A2(new_n717), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n604), .A2(new_n368), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n705), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  AND2_X1   g543(.A1(new_n659), .A2(new_n697), .ZN(new_n730));
  INV_X1    g544(.A(new_n325), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n721), .B2(new_n722), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g548(.A1(G472), .A2(new_n629), .B1(new_n734), .B2(new_n329), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT104), .B1(new_n735), .B2(new_n650), .ZN(new_n736));
  AND4_X1   g550(.A1(KEYINPUT104), .A2(new_n717), .A3(new_n650), .A4(new_n724), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n689), .B(new_n730), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n335), .A2(new_n740), .A3(new_n555), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT107), .B1(new_n711), .B2(new_n554), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n594), .A2(new_n743), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n587), .A2(new_n589), .B1(new_n592), .B2(new_n584), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(KEYINPUT105), .A3(G469), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n586), .A3(new_n596), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n599), .A3(new_n604), .A4(new_n610), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n618), .A2(new_n507), .A3(new_n446), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n662), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n748), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n741), .A2(new_n742), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT105), .B1(new_n745), .B2(G469), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n588), .B1(new_n571), .B2(new_n577), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n591), .B(new_n583), .C1(new_n569), .C2(new_n570), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n743), .A4(new_n556), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n586), .A2(new_n596), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n598), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n611), .A3(new_n751), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n711), .A3(new_n554), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n755), .B1(new_n764), .B2(KEYINPUT42), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n711), .A2(new_n554), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n748), .A2(new_n752), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(KEYINPUT106), .A3(new_n749), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n754), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n212), .ZN(G33));
  NAND3_X1  g585(.A1(new_n427), .A2(new_n368), .A3(new_n437), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n772), .A2(new_n639), .A3(new_n750), .A4(new_n662), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n335), .A2(new_n555), .A3(new_n773), .A4(new_n762), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  NAND3_X1  g589(.A1(new_n641), .A2(new_n431), .A3(new_n610), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n630), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n650), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT110), .ZN(new_n783));
  INV_X1    g597(.A(new_n750), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(KEYINPUT110), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n590), .A2(new_n593), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n745), .A2(KEYINPUT108), .A3(KEYINPUT45), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n556), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n790), .A2(new_n791), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n595), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT46), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n586), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n599), .A3(new_n677), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT109), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n780), .A2(new_n781), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n783), .A2(KEYINPUT111), .A3(new_n784), .A4(new_n785), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n788), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n599), .ZN(new_n806));
  XNOR2_X1  g620(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n799), .A2(new_n599), .A3(new_n807), .ZN(new_n810));
  AOI211_X1 g624(.A(new_n624), .B(new_n662), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n335), .A2(new_n555), .A3(new_n750), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT102), .B1(new_n713), .B2(new_n706), .ZN(new_n816));
  AND4_X1   g630(.A1(KEYINPUT102), .A2(new_n705), .A3(new_n335), .A4(new_n706), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n627), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n335), .A2(new_n555), .A3(new_n697), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n728), .B(new_n703), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n815), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n725), .A2(new_n712), .A3(new_n666), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n698), .B2(new_n627), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n715), .A2(new_n824), .A3(KEYINPUT114), .A4(new_n703), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n624), .B1(new_n369), .B2(new_n604), .ZN(new_n827));
  INV_X1    g641(.A(new_n510), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n630), .A4(new_n628), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n602), .A2(new_n774), .A3(new_n651), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n717), .A2(new_n724), .A3(new_n650), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT104), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n717), .A2(new_n724), .A3(KEYINPUT104), .A4(new_n650), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n748), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n640), .A2(new_n641), .A3(new_n369), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n711), .A2(new_n654), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n751), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n830), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n770), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n650), .A2(new_n662), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n762), .A2(new_n659), .A3(new_n727), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n841), .B(new_n842), .C1(new_n673), .C2(new_n674), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n658), .B(new_n659), .C1(new_n663), .C2(new_n689), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n738), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n738), .A3(new_n844), .A4(KEYINPUT52), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n826), .A2(new_n840), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n822), .A2(new_n825), .B1(new_n847), .B2(new_n848), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(KEYINPUT53), .A3(new_n840), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n850), .A2(new_n856), .A3(new_n851), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n853), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n778), .A2(new_n440), .A3(new_n726), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n730), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n686), .A2(new_n446), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n697), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT50), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n860), .A2(new_n865), .A3(new_n697), .A4(new_n862), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n697), .A2(new_n784), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n675), .A2(new_n440), .A3(new_n555), .A4(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n604), .A2(new_n610), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n864), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n692), .A2(new_n696), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n598), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n809), .A2(new_n810), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n784), .A3(new_n860), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n778), .A2(new_n440), .A3(new_n867), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n736), .B2(new_n737), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n871), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n871), .A2(new_n875), .A3(KEYINPUT51), .A4(new_n877), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n741), .A2(new_n742), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT48), .Z(new_n884));
  XOR2_X1   g698(.A(new_n439), .B(KEYINPUT119), .Z(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n868), .B2(new_n624), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n861), .A2(new_n880), .A3(new_n881), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT115), .B(KEYINPUT53), .C1(new_n854), .C2(new_n840), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n856), .B1(new_n850), .B2(new_n851), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n889), .B1(new_n892), .B2(new_n855), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n894));
  INV_X1    g708(.A(new_n754), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n764), .A2(new_n755), .A3(KEYINPUT42), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT106), .B1(new_n768), .B2(new_n749), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n821), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(KEYINPUT118), .A3(new_n715), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n839), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n900), .A2(new_n849), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT53), .B1(new_n839), .B2(new_n901), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n898), .A2(new_n715), .A3(new_n899), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n903), .A2(new_n907), .B1(new_n851), .B2(new_n850), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n894), .B1(new_n908), .B2(new_n889), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n859), .B(new_n888), .C1(new_n893), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT120), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n872), .B(KEYINPUT49), .Z(new_n914));
  NOR3_X1   g728(.A1(new_n914), .A2(new_n686), .A3(new_n776), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n554), .A2(new_n612), .A3(new_n598), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT113), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n675), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n913), .A2(KEYINPUT121), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(G75));
  NOR2_X1   g737(.A1(new_n908), .A2(new_n364), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(G210), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n501), .A2(new_n503), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n504), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n925), .B2(new_n926), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n281), .A2(G952), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT122), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(G51));
  OR3_X1    g748(.A1(new_n908), .A2(KEYINPUT123), .A3(new_n889), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT123), .B1(new_n908), .B2(new_n889), .ZN(new_n936));
  INV_X1    g750(.A(new_n908), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n935), .B(new_n936), .C1(new_n937), .C2(KEYINPUT54), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n595), .B(KEYINPUT57), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n695), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n924), .A2(new_n795), .A3(new_n794), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n932), .B1(new_n942), .B2(new_n943), .ZN(G54));
  NAND3_X1  g758(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n945));
  INV_X1    g759(.A(new_n638), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n932), .ZN(G60));
  XOR2_X1   g763(.A(new_n608), .B(KEYINPUT59), .Z(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n605), .B2(new_n606), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n938), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n933), .ZN(new_n953));
  INV_X1    g767(.A(new_n909), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n858), .A2(KEYINPUT54), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n950), .B1(new_n956), .B2(new_n859), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n605), .A2(new_n606), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n952), .B(new_n953), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(G63));
  NAND2_X1  g774(.A1(G217), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT124), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n937), .A2(new_n648), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n937), .A2(new_n963), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n537), .A2(new_n541), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n953), .B(new_n964), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g782(.A(new_n281), .B1(new_n442), .B2(G224), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n826), .A2(new_n602), .A3(new_n651), .A4(new_n829), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT125), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n971), .B2(new_n281), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n927), .B1(G898), .B2(new_n281), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT126), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G69));
  NAND3_X1  g789(.A1(new_n788), .A2(new_n802), .A3(new_n803), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n882), .A2(new_n659), .A3(new_n727), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n801), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n738), .A2(new_n844), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n813), .A2(new_n774), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n898), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n281), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n297), .A2(new_n302), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n395), .A2(new_n397), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(G227), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(G900), .A3(G953), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n983), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n990));
  INV_X1    g804(.A(new_n986), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n766), .A2(new_n678), .A3(new_n784), .A4(new_n827), .ZN(new_n992));
  NAND2_X1  g806(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n687), .A2(new_n980), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n687), .A2(new_n980), .ZN(new_n995));
  XNOR2_X1  g809(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n995), .A2(new_n996), .B1(new_n811), .B2(new_n812), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n804), .A2(new_n992), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n990), .B(new_n991), .C1(new_n998), .C2(G953), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n989), .A2(new_n999), .ZN(G72));
  INV_X1    g814(.A(new_n932), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n982), .B2(new_n971), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1004), .A2(new_n268), .A3(new_n306), .A4(new_n304), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1003), .B1(new_n998), .B2(new_n971), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n286), .A3(new_n305), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n305), .A2(new_n306), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n326), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n858), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1010));
  AND4_X1   g824(.A1(new_n1001), .A2(new_n1005), .A3(new_n1007), .A4(new_n1010), .ZN(G57));
endmodule


