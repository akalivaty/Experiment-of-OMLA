//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021;
  INV_X1    g000(.A(G43gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G43gat), .A2(G50gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OR3_X1    g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n204), .A2(new_n214), .A3(new_n205), .ZN(new_n215));
  AND4_X1   g014(.A1(new_n207), .A2(new_n210), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(KEYINPUT85), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n218), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n211), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n207), .B1(new_n220), .B2(new_n208), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT17), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n208), .ZN(new_n223));
  INV_X1    g022(.A(new_n207), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n213), .A4(new_n215), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G22gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G15gat), .ZN(new_n231));
  INV_X1    g030(.A(G15gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT87), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n231), .B2(new_n233), .ZN(new_n236));
  INV_X1    g035(.A(G1gat), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(KEYINPUT16), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n233), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT87), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(G8gat), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G8gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n241), .A3(G1gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n235), .A2(new_n236), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n245), .B(new_n246), .C1(new_n247), .C2(new_n239), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n229), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n225), .A2(new_n227), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n244), .A2(new_n251), .A3(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(G229gat), .A2(G233gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT88), .Z(new_n254));
  NAND4_X1  g053(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(KEYINPUT13), .Z(new_n256));
  INV_X1    g055(.A(new_n252), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n251), .B1(new_n244), .B2(new_n248), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT18), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT89), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G141gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT11), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G169gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G197gat), .ZN(new_n269));
  INV_X1    g068(.A(G169gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n267), .B(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G197gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT12), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT12), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n269), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n260), .B(new_n263), .C1(new_n264), .C2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n277), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n276), .B1(new_n269), .B2(new_n273), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n255), .A2(new_n259), .A3(new_n264), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n222), .A2(new_n228), .B1(new_n244), .B2(new_n248), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n257), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT18), .B1(new_n285), .B2(new_n254), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n255), .A2(new_n259), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n282), .B(new_n283), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n291));
  AND2_X1   g090(.A1(G57gat), .A2(G64gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G57gat), .A2(G64gat), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT91), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n297));
  INV_X1    g096(.A(G71gat), .ZN(new_n298));
  INV_X1    g097(.A(G78gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT90), .B1(G71gat), .B2(G78gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(G71gat), .A2(G78gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n296), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI211_X1 g104(.A(KEYINPUT91), .B(new_n303), .C1(new_n300), .C2(new_n301), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n295), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(G71gat), .A2(G78gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n294), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n249), .B1(new_n290), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n290), .ZN(new_n313));
  NAND2_X1  g112(.A1(G231gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n310), .A2(new_n290), .A3(new_n314), .ZN(new_n317));
  XNOR2_X1  g116(.A(G127gat), .B(G155gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n316), .B2(new_n317), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n312), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  INV_X1    g122(.A(new_n312), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n311), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(new_n325), .A3(new_n311), .ZN(new_n328));
  XOR2_X1   g127(.A(G183gat), .B(G211gat), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n328), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n329), .B1(new_n332), .B2(new_n326), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT96), .ZN(new_n336));
  NAND3_X1  g135(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n337));
  OR2_X1    g136(.A1(G99gat), .A2(G106gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT95), .ZN(new_n339));
  NAND2_X1  g138(.A1(G99gat), .A2(G106gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(G99gat), .A2(G106gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(G99gat), .A2(G106gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT95), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(KEYINPUT8), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT94), .ZN(new_n347));
  INV_X1    g146(.A(G85gat), .ZN(new_n348));
  INV_X1    g147(.A(G92gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n347), .B1(new_n346), .B2(new_n350), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n348), .B2(new_n349), .ZN(new_n355));
  OAI211_X1 g154(.A(G85gat), .B(G92gat), .C1(KEYINPUT93), .C2(KEYINPUT7), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n355), .A2(new_n356), .B1(KEYINPUT93), .B2(KEYINPUT7), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n345), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT8), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(G99gat), .B2(G106gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(G85gat), .A2(G92gat), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT94), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n341), .A2(new_n344), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(new_n356), .ZN(new_n366));
  NAND2_X1  g165(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n358), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n216), .A2(new_n221), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n337), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n222), .A2(new_n228), .B1(new_n369), .B2(new_n358), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G190gat), .B(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n336), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G134gat), .B(G162gat), .Z(new_n378));
  AOI21_X1  g177(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n374), .B2(new_n376), .ZN(new_n381));
  OAI211_X1 g180(.A(KEYINPUT96), .B(new_n375), .C1(new_n372), .C2(new_n373), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n380), .B(KEYINPUT92), .Z(new_n384));
  NOR2_X1   g183(.A1(new_n374), .A2(new_n376), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT97), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n383), .B2(new_n387), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n364), .A2(new_n368), .A3(new_n365), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n365), .B1(new_n364), .B2(new_n368), .ZN(new_n394));
  INV_X1    g193(.A(new_n301), .ZN(new_n395));
  NOR3_X1   g194(.A1(KEYINPUT90), .A2(G71gat), .A3(G78gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n304), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT91), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n302), .A2(new_n296), .A3(new_n304), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n294), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n309), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n393), .A2(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n358), .A2(new_n369), .A3(new_n307), .A4(new_n309), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n400), .A2(new_n401), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n406), .A2(KEYINPUT10), .A3(new_n369), .A4(new_n358), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G230gat), .A2(G233gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n402), .B2(new_n404), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G120gat), .B(G148gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT98), .ZN(new_n414));
  XOR2_X1   g213(.A(G176gat), .B(G204gat), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  INV_X1    g217(.A(new_n409), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n419), .B1(new_n405), .B2(new_n407), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n418), .B1(new_n420), .B2(new_n411), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n417), .A2(KEYINPUT99), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT99), .B1(new_n417), .B2(new_n421), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n335), .A2(new_n392), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428));
  OR2_X1    g227(.A1(G113gat), .A2(G120gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT1), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT67), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT67), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT1), .ZN(new_n433));
  NAND2_X1  g232(.A1(G113gat), .A2(G120gat), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n429), .A2(new_n431), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G127gat), .B(G134gat), .Z(new_n436));
  OAI21_X1  g235(.A(new_n428), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n429), .A2(new_n434), .ZN(new_n438));
  XNOR2_X1  g237(.A(G127gat), .B(G134gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n438), .A2(KEYINPUT68), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n430), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n437), .A2(new_n441), .B1(new_n442), .B2(new_n436), .ZN(new_n443));
  NOR2_X1   g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT23), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT23), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(G169gat), .B2(G176gat), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT24), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n448), .A2(new_n449), .B1(G183gat), .B2(G190gat), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT65), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n451));
  OAI221_X1 g250(.A(new_n445), .B1(new_n444), .B2(new_n447), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n445), .B1(new_n447), .B2(new_n444), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT25), .ZN(new_n454));
  NAND2_X1  g253(.A1(G183gat), .A2(G190gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT64), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT64), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n452), .A2(KEYINPUT25), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT26), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(new_n444), .ZN(new_n466));
  INV_X1    g265(.A(G183gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT27), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT27), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G183gat), .ZN(new_n470));
  INV_X1    g269(.A(G190gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT28), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT66), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n472), .B2(KEYINPUT66), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n455), .B(new_n466), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  AOI211_X1 g276(.A(new_n427), .B(new_n443), .C1(new_n462), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n477), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n437), .A2(new_n441), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n442), .A2(new_n436), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n450), .A2(new_n451), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT25), .B1(new_n484), .B2(new_n453), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n454), .A2(new_n461), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(new_n443), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n478), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT34), .ZN(new_n490));
  NAND2_X1  g289(.A1(G227gat), .A2(G233gat), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n489), .A2(KEYINPUT72), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n483), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n479), .A2(KEYINPUT69), .A3(new_n482), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n493), .A2(new_n490), .A3(new_n491), .A4(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n491), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT34), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n492), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G15gat), .B(G43gat), .Z(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT70), .ZN(new_n502));
  XNOR2_X1  g301(.A(G71gat), .B(G99gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(KEYINPUT33), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT32), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n510));
  INV_X1    g309(.A(new_n491), .ZN(new_n511));
  AOI221_X4 g310(.A(new_n507), .B1(KEYINPUT33), .B2(new_n504), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n500), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT32), .B1(new_n489), .B2(new_n491), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(new_n504), .C1(KEYINPUT33), .C2(new_n505), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n492), .A2(new_n497), .A3(new_n499), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT79), .B(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G228gat), .A2(G233gat), .ZN(new_n522));
  XOR2_X1   g321(.A(G155gat), .B(G162gat), .Z(new_n523));
  INV_X1    g322(.A(G141gat), .ZN(new_n524));
  INV_X1    g323(.A(G148gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G141gat), .A2(G148gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n523), .B1(KEYINPUT2), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n528), .ZN(new_n530));
  XNOR2_X1  g329(.A(G155gat), .B(G162gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT2), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT75), .B(G155gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(G162gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n529), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(G211gat), .A2(G218gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(G211gat), .A2(G218gat), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G197gat), .B(G204gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(KEYINPUT22), .B2(new_n537), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n539), .B(new_n541), .C1(KEYINPUT22), .C2(new_n537), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT29), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n536), .B1(new_n545), .B2(KEYINPUT3), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n522), .B1(new_n546), .B2(KEYINPUT78), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT3), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n529), .B(new_n548), .C1(new_n532), .C2(new_n535), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(new_n544), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n553), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n521), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G78gat), .B(G106gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G50gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(G22gat), .A3(new_n555), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n560), .B(KEYINPUT77), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n554), .A2(new_n555), .A3(new_n521), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n556), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G226gat), .A2(G233gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n486), .A2(new_n485), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n466), .A2(new_n455), .ZN(new_n569));
  INV_X1    g368(.A(new_n476), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(new_n474), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n567), .B1(new_n572), .B2(KEYINPUT29), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n567), .B(KEYINPUT73), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n568), .B2(new_n571), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n479), .A2(KEYINPUT74), .A3(new_n574), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n573), .A2(new_n577), .A3(new_n552), .A4(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n552), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n574), .B1(new_n479), .B2(new_n550), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n572), .A2(new_n567), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n584));
  XNOR2_X1  g383(.A(G8gat), .B(G36gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G64gat), .B(G92gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n579), .A2(new_n583), .A3(new_n584), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n579), .A2(new_n583), .A3(new_n588), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT30), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n579), .B2(new_n583), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n519), .A2(new_n566), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT4), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n482), .A2(new_n595), .A3(new_n536), .ZN(new_n596));
  INV_X1    g395(.A(new_n535), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n523), .A2(new_n528), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n530), .A2(new_n533), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n597), .A2(new_n598), .B1(new_n599), .B2(new_n523), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT4), .B1(new_n443), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT76), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n443), .A2(new_n600), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n595), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT76), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n443), .A2(new_n600), .A3(KEYINPUT4), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n536), .A2(KEYINPUT3), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n482), .A3(new_n549), .ZN(new_n609));
  NAND2_X1  g408(.A1(G225gat), .A2(G233gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT5), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n602), .A2(new_n607), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n482), .A2(new_n536), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n443), .A2(new_n600), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n604), .A2(new_n606), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n609), .A2(new_n610), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n616), .B(KEYINPUT5), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G1gat), .B(G29gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT0), .ZN(new_n622));
  XNOR2_X1  g421(.A(G57gat), .B(G85gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT6), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n613), .A2(new_n619), .A3(new_n624), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n620), .A2(KEYINPUT6), .A3(new_n625), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT83), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n624), .B1(new_n613), .B2(new_n619), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n629), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT35), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n594), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n514), .A3(new_n516), .ZN(new_n640));
  OAI211_X1 g439(.A(KEYINPUT71), .B(new_n517), .C1(new_n509), .C2(new_n512), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n566), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT84), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT84), .A4(new_n566), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n593), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n638), .B1(new_n650), .B2(KEYINPUT35), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT36), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n640), .B2(new_n641), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT36), .B1(new_n513), .B2(new_n518), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n566), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n602), .A2(new_n607), .A3(new_n609), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n611), .ZN(new_n659));
  INV_X1    g458(.A(new_n609), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n617), .B2(KEYINPUT76), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n610), .B1(new_n661), .B2(new_n607), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n482), .A2(new_n536), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n603), .A3(new_n610), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n658), .B1(new_n664), .B2(KEYINPUT80), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(KEYINPUT80), .B2(new_n664), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n659), .B(new_n624), .C1(new_n662), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT81), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n626), .B(new_n589), .C1(new_n591), .C2(new_n592), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n667), .A2(KEYINPUT81), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n633), .A2(KEYINPUT6), .ZN(new_n675));
  AOI211_X1 g474(.A(new_n627), .B(new_n624), .C1(new_n613), .C2(new_n619), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n675), .A2(new_n628), .B1(new_n676), .B2(KEYINPUT83), .ZN(new_n677));
  INV_X1    g476(.A(new_n590), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT37), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n579), .A2(new_n583), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n680), .A2(new_n587), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n574), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n572), .B2(KEYINPUT29), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n479), .A2(G226gat), .A3(G233gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n679), .B1(new_n687), .B2(new_n552), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n573), .A2(new_n577), .A3(new_n580), .A4(new_n578), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n678), .B1(new_n681), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n680), .A2(new_n587), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n679), .B1(new_n579), .B2(new_n583), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n683), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n677), .A2(new_n691), .A3(new_n632), .A4(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n656), .B1(new_n674), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n656), .A2(new_n646), .A3(new_n593), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n655), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n289), .B(new_n426), .C1(new_n651), .C2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n646), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(new_n237), .ZN(G1324gat));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n593), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT102), .ZN(new_n707));
  OAI21_X1  g506(.A(G8gat), .B1(new_n701), .B2(new_n593), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT101), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n705), .B(KEYINPUT100), .Z(new_n710));
  AND2_X1   g509(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n707), .B(new_n709), .C1(KEYINPUT42), .C2(new_n711), .ZN(G1325gat));
  OAI21_X1  g511(.A(G15gat), .B1(new_n701), .B2(new_n655), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n519), .A2(new_n232), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n701), .B2(new_n714), .ZN(G1326gat));
  OR3_X1    g514(.A1(new_n701), .A2(KEYINPUT103), .A3(new_n566), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT103), .B1(new_n701), .B2(new_n566), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  INV_X1    g519(.A(new_n392), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n334), .A2(new_n721), .A3(new_n425), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n289), .B(new_n722), .C1(new_n651), .C2(new_n700), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(G29gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n725), .A3(new_n647), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  INV_X1    g526(.A(new_n289), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n334), .A2(new_n728), .A3(new_n425), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n650), .A2(KEYINPUT35), .ZN(new_n731));
  INV_X1    g530(.A(new_n638), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n667), .A2(KEYINPUT81), .A3(new_n672), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n672), .B1(new_n667), .B2(KEYINPUT81), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n735), .A2(new_n736), .A3(new_n670), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n688), .A2(new_n689), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n738), .A2(new_n587), .A3(new_n680), .A4(new_n682), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n694), .A2(new_n590), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n635), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n566), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n697), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n734), .B1(new_n743), .B2(new_n655), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n655), .B(new_n734), .C1(new_n696), .C2(new_n698), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n733), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n392), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n392), .B1(new_n651), .B2(new_n700), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT44), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n730), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n647), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n727), .B1(new_n754), .B2(new_n725), .ZN(G1328gat));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757));
  INV_X1    g556(.A(G36gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n648), .A2(new_n758), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n723), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n757), .B1(new_n723), .B2(new_n759), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n753), .A2(new_n648), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(G36gat), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n756), .A3(new_n761), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(KEYINPUT107), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(KEYINPUT107), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(G1329gat));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n519), .A2(new_n202), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n723), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(KEYINPUT108), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n655), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n202), .B1(new_n753), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n775), .B2(new_n771), .ZN(new_n776));
  INV_X1    g575(.A(new_n771), .ZN(new_n777));
  AOI211_X1 g576(.A(new_n655), .B(new_n730), .C1(new_n750), .C2(new_n752), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n777), .B(new_n772), .C1(new_n778), .C2(new_n202), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1330gat));
  NAND2_X1  g579(.A1(new_n750), .A2(new_n752), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(new_n656), .A3(new_n729), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n566), .A2(G50gat), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n782), .A2(G50gat), .B1(new_n724), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n785));
  AOI21_X1  g584(.A(new_n203), .B1(new_n753), .B2(new_n656), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n724), .B2(new_n783), .ZN(new_n788));
  NOR4_X1   g587(.A1(new_n723), .A2(KEYINPUT110), .A3(G50gat), .A4(new_n566), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT48), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n784), .A2(new_n785), .B1(new_n786), .B2(new_n790), .ZN(G1331gat));
  NAND2_X1  g590(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n651), .B1(new_n792), .B2(new_n745), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n334), .A2(new_n721), .A3(new_n728), .A4(new_n425), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n647), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n648), .ZN(new_n798));
  NOR2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  AND2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n799), .B2(new_n798), .ZN(G1333gat));
  NAND3_X1  g601(.A1(new_n795), .A2(new_n298), .A3(new_n519), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n793), .A2(new_n655), .A3(new_n794), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n298), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g605(.A1(new_n795), .A2(new_n656), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT111), .B(G78gat), .Z(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1335gat));
  NOR2_X1   g608(.A1(new_n646), .A2(G85gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n745), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n721), .B1(new_n811), .B2(new_n733), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n334), .A2(new_n289), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT51), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815));
  INV_X1    g614(.A(new_n813), .ZN(new_n816));
  NOR4_X1   g615(.A1(new_n793), .A2(new_n815), .A3(new_n721), .A4(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n814), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n747), .A2(new_n392), .A3(new_n813), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n815), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n812), .A2(KEYINPUT51), .A3(new_n813), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT112), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n425), .B(new_n810), .C1(new_n819), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n813), .A2(new_n425), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n750), .B2(new_n752), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n647), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G85gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(G1336gat));
  AOI21_X1  g628(.A(new_n349), .B1(new_n826), .B2(new_n648), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n424), .A2(G92gat), .A3(new_n593), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n821), .B2(new_n822), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT52), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n831), .B1(new_n814), .B2(new_n817), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n593), .B(new_n825), .C1(new_n750), .C2(new_n752), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n349), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n834), .A2(new_n838), .ZN(G1337gat));
  AOI21_X1  g638(.A(G99gat), .B1(new_n513), .B2(new_n518), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n425), .B(new_n840), .C1(new_n819), .C2(new_n823), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n774), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G99gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1338gat));
  XNOR2_X1  g643(.A(KEYINPUT113), .B(G106gat), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n845), .B1(new_n826), .B2(new_n656), .ZN(new_n846));
  OR3_X1    g645(.A1(new_n566), .A2(new_n424), .A3(G106gat), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT114), .Z(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n821), .B2(new_n822), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT53), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n814), .B2(new_n817), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n566), .B(new_n825), .C1(new_n750), .C2(new_n752), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n845), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n855), .ZN(G1339gat));
  NAND4_X1  g655(.A1(new_n278), .A2(new_n263), .A3(new_n259), .A4(new_n255), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n285), .A2(new_n254), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n257), .A2(new_n258), .A3(new_n256), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n274), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n422), .B2(new_n423), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n405), .A2(new_n407), .A3(new_n419), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n410), .A2(KEYINPUT54), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n416), .B1(new_n420), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(KEYINPUT55), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n405), .A2(new_n407), .A3(new_n419), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(new_n420), .A3(new_n865), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n408), .A2(new_n865), .A3(new_n409), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n418), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n289), .A2(new_n417), .A3(new_n867), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n392), .B1(new_n862), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n383), .A2(new_n387), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT97), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n389), .A3(new_n861), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n417), .A3(new_n867), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n335), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n334), .A2(new_n721), .A3(new_n728), .A4(new_n424), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n646), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n644), .A2(new_n645), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n593), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n289), .ZN(new_n887));
  INV_X1    g686(.A(G113gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n594), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n883), .A2(G113gat), .A3(new_n890), .A4(new_n289), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n889), .A2(KEYINPUT115), .A3(new_n891), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1340gat));
  NOR2_X1   g695(.A1(new_n424), .A2(G120gat), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT116), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n890), .ZN(new_n900));
  OAI21_X1  g699(.A(G120gat), .B1(new_n900), .B2(new_n424), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1341gat));
  INV_X1    g701(.A(G127gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n903), .A3(new_n334), .ZN(new_n904));
  OAI21_X1  g703(.A(G127gat), .B1(new_n900), .B2(new_n335), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1342gat));
  INV_X1    g705(.A(G134gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n721), .A2(new_n648), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n885), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT56), .Z(new_n910));
  OAI21_X1  g709(.A(G134gat), .B1(new_n900), .B2(new_n721), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1343gat));
  NAND2_X1  g711(.A1(new_n655), .A2(new_n656), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT118), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n593), .A3(new_n883), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n524), .B1(new_n915), .B2(new_n728), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n867), .A2(new_n417), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n873), .A2(KEYINPUT117), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n919), .B(new_n868), .C1(new_n870), .C2(new_n872), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n917), .A2(new_n918), .A3(new_n289), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n392), .B1(new_n921), .B2(new_n862), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n335), .B1(new_n922), .B2(new_n880), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n566), .B1(new_n923), .B2(new_n882), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n655), .A2(new_n647), .A3(new_n593), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n566), .B1(new_n881), .B2(new_n882), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n289), .A2(G141gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n916), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g731(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n933));
  XOR2_X1   g732(.A(new_n932), .B(new_n933), .Z(G1344gat));
  INV_X1    g733(.A(KEYINPUT59), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n874), .A2(new_n862), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n721), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n878), .A2(new_n879), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n334), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n882), .ZN(new_n940));
  OAI211_X1 g739(.A(KEYINPUT57), .B(new_n656), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n941), .B1(new_n924), .B2(KEYINPUT57), .ZN(new_n942));
  INV_X1    g741(.A(new_n927), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n425), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT120), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n525), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(KEYINPUT120), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n935), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n930), .A2(new_n424), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(KEYINPUT59), .A3(new_n525), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n425), .A2(new_n525), .ZN(new_n951));
  OAI22_X1  g750(.A1(new_n948), .A2(new_n950), .B1(new_n915), .B2(new_n951), .ZN(G1345gat));
  OR3_X1    g751(.A1(new_n915), .A2(new_n534), .A3(new_n335), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n534), .B1(new_n930), .B2(new_n335), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT121), .ZN(G1346gat));
  OAI21_X1  g755(.A(G162gat), .B1(new_n930), .B2(new_n721), .ZN(new_n957));
  INV_X1    g756(.A(G162gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n914), .A2(new_n958), .A3(new_n883), .A4(new_n908), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1347gat));
  NAND2_X1  g759(.A1(new_n881), .A2(new_n882), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n884), .A2(new_n648), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(KEYINPUT122), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(KEYINPUT122), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n646), .B(new_n961), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n965), .A2(G169gat), .A3(new_n728), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n647), .A2(new_n593), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(new_n566), .A3(new_n519), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n961), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G169gat), .B1(new_n971), .B2(new_n728), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT124), .Z(new_n973));
  NAND2_X1  g772(.A1(new_n968), .A2(new_n973), .ZN(G1348gat));
  OAI21_X1  g773(.A(G176gat), .B1(new_n971), .B2(new_n424), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n424), .A2(G176gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n965), .B2(new_n976), .ZN(G1349gat));
  OAI21_X1  g776(.A(G183gat), .B1(new_n971), .B2(new_n335), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n334), .A2(new_n468), .A3(new_n470), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n965), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g780(.A(G190gat), .B1(new_n971), .B2(new_n721), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n392), .A2(new_n471), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n965), .B2(new_n984), .ZN(G1351gat));
  AND2_X1   g784(.A1(new_n655), .A2(new_n969), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n928), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(new_n272), .A3(new_n289), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n942), .A2(new_n986), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n728), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(G197gat), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n990), .A2(new_n989), .A3(new_n728), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(G1352gat));
  INV_X1    g793(.A(new_n987), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n995), .A2(G204gat), .A3(new_n424), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n996), .B(KEYINPUT62), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n942), .A2(new_n425), .A3(new_n986), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(G204gat), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n997), .A2(new_n999), .ZN(G1353gat));
  NAND2_X1  g799(.A1(new_n923), .A2(new_n882), .ZN(new_n1001));
  AOI21_X1  g800(.A(KEYINPUT57), .B1(new_n1001), .B2(new_n656), .ZN(new_n1002));
  AOI211_X1 g801(.A(new_n925), .B(new_n566), .C1(new_n881), .C2(new_n882), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n334), .B(new_n986), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(KEYINPUT126), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n1006));
  NAND4_X1  g805(.A1(new_n942), .A2(new_n1006), .A3(new_n334), .A4(new_n986), .ZN(new_n1007));
  NAND4_X1  g806(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(KEYINPUT127), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n1007), .A2(G211gat), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1011));
  NAND4_X1  g810(.A1(new_n1010), .A2(new_n1011), .A3(KEYINPUT63), .A4(new_n1005), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT63), .ZN(new_n1013));
  INV_X1    g812(.A(new_n1005), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1007), .A2(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1009), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  OR3_X1    g816(.A1(new_n995), .A2(G211gat), .A3(new_n335), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(new_n1018), .ZN(G1354gat));
  OAI21_X1  g818(.A(G218gat), .B1(new_n990), .B2(new_n721), .ZN(new_n1020));
  OR2_X1    g819(.A1(new_n721), .A2(G218gat), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1020), .B1(new_n995), .B2(new_n1021), .ZN(G1355gat));
endmodule


