//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  XOR2_X1   g000(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT27), .Z(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT67), .B1(new_n195), .B2(G116), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(G119), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n201), .B1(new_n196), .B2(new_n199), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT68), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT2), .B(G113), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(new_n208), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT1), .B1(new_n216), .B2(G146), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT66), .A3(KEYINPUT1), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT64), .A2(G143), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT64), .A2(G143), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n220), .A2(G143), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n219), .A2(new_n222), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g042(.A1(KEYINPUT64), .A2(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT64), .A2(G143), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G146), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n221), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n214), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n217), .A2(new_n218), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(G128), .A3(new_n222), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n225), .A2(new_n227), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT69), .A3(new_n233), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT65), .B(G131), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G137), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G134), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n242), .B2(G137), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n243), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n243), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n242), .A2(G137), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n235), .A2(new_n240), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n231), .A2(new_n221), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n238), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(new_n243), .A3(new_n245), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(new_n248), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n255), .B(new_n258), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n253), .A2(KEYINPUT71), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT71), .B1(new_n253), .B2(new_n262), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n213), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n213), .A2(new_n253), .A3(new_n262), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n252), .B1(new_n234), .B2(new_n228), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n262), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n212), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT28), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n194), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n253), .B2(new_n262), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n270), .A2(KEYINPUT30), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n212), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(new_n268), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT31), .A4(new_n194), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n278), .A2(new_n280), .A3(new_n194), .A4(new_n268), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n274), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n187), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n267), .A2(new_n273), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n193), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n282), .A2(new_n283), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n282), .A2(new_n283), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT32), .A3(new_n286), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n278), .A2(new_n268), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT29), .B1(new_n295), .B2(new_n193), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n253), .A2(new_n262), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n253), .A2(KEYINPUT71), .A3(new_n262), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n212), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n194), .B(new_n273), .C1(new_n302), .C2(KEYINPUT28), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n296), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n297), .B1(new_n296), .B2(new_n303), .ZN(new_n305));
  INV_X1    g119(.A(new_n268), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n213), .B1(new_n253), .B2(new_n262), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT28), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n194), .A2(KEYINPUT29), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n267), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT74), .B(G902), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n304), .A2(new_n305), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G472), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n288), .B(new_n294), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n311), .B2(G234), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n311), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n195), .B2(G128), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n215), .A2(KEYINPUT23), .A3(G119), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n321), .B(new_n322), .C1(G119), .C2(new_n215), .ZN(new_n323));
  XNOR2_X1  g137(.A(G119), .B(G128), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT24), .B(G110), .Z(new_n325));
  AOI22_X1  g139(.A1(new_n323), .A2(G110), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G125), .B(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n329), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(G146), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(G146), .B1(new_n328), .B2(new_n330), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n326), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT75), .B(G110), .ZN(new_n335));
  OAI22_X1  g149(.A1(new_n323), .A2(new_n335), .B1(new_n324), .B2(new_n325), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(KEYINPUT77), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n328), .A2(new_n339), .A3(G146), .A4(new_n330), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n342));
  OAI221_X1 g156(.A(new_n342), .B1(new_n325), .B2(new_n324), .C1(new_n323), .C2(new_n335), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n327), .A2(new_n220), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n334), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G137), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n347), .A2(KEYINPUT78), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(KEYINPUT78), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n348), .B2(new_n349), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n334), .B(new_n353), .C1(new_n341), .C2(new_n345), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n319), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n318), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n343), .A2(new_n344), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n338), .A2(new_n340), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(new_n337), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n353), .B1(new_n362), .B2(new_n334), .ZN(new_n363));
  INV_X1    g177(.A(new_n356), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n311), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n355), .A2(new_n356), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n317), .A2(G902), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n315), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT88), .ZN(new_n374));
  XNOR2_X1  g188(.A(G113), .B(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT86), .B(G104), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(new_n216), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT64), .B(G143), .ZN(new_n382));
  INV_X1    g196(.A(G214), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n383), .A2(G237), .A3(G953), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n223), .A2(new_n224), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT83), .B1(new_n387), .B2(new_n379), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n381), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n241), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT84), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n385), .B1(new_n382), .B2(new_n384), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n380), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n392), .B1(new_n395), .B2(new_n241), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n241), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n327), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(KEYINPUT19), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n398), .B(new_n361), .C1(G146), .C2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n389), .A2(KEYINPUT18), .A3(G131), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT18), .A2(G131), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n327), .B(new_n220), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n378), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n407), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n391), .A2(new_n396), .A3(new_n410), .A4(new_n397), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n332), .A2(new_n333), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n391), .A2(new_n396), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(new_n415), .B2(KEYINPUT17), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n412), .B1(new_n416), .B2(KEYINPUT87), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n410), .B1(new_n391), .B2(new_n396), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(new_n414), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n409), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n408), .B1(new_n421), .B2(new_n378), .ZN(new_n422));
  NOR2_X1   g236(.A1(G475), .A2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n374), .B(KEYINPUT20), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT84), .B1(new_n389), .B2(new_n390), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n395), .A2(new_n392), .A3(new_n241), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT17), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT87), .A3(new_n413), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n420), .A3(new_n411), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n407), .A3(new_n378), .ZN(new_n431));
  INV_X1    g245(.A(new_n408), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n424), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT88), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n434), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n425), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n431), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n378), .B1(new_n430), .B2(new_n407), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G475), .ZN(new_n442));
  XNOR2_X1  g256(.A(G116), .B(G122), .ZN(new_n443));
  INV_X1    g257(.A(G107), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n445), .B(KEYINPUT90), .Z(new_n446));
  NAND2_X1  g260(.A1(new_n387), .A2(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n215), .A2(G143), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n242), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n242), .B1(new_n447), .B2(new_n448), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT14), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n198), .A3(G122), .ZN(new_n453));
  INV_X1    g267(.A(G122), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT14), .B1(new_n454), .B2(G116), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(G116), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n457), .A2(G107), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT91), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  OAI221_X1 g275(.A(new_n446), .B1(new_n450), .B2(new_n451), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n443), .B(new_n444), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n449), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT13), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT89), .B1(new_n447), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n387), .A2(new_n467), .A3(KEYINPUT13), .A4(G128), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n447), .A2(new_n465), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n466), .A2(new_n468), .A3(new_n448), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n464), .B1(new_n470), .B2(G134), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT9), .B(G234), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n316), .A3(G953), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n462), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n462), .B2(new_n472), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n311), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G478), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT15), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI221_X1 g294(.A(new_n311), .B1(KEYINPUT15), .B2(new_n478), .C1(new_n475), .C2(new_n476), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(G234), .A2(G237), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(G952), .A3(new_n189), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT92), .Z(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n319), .A2(G953), .A3(new_n484), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT21), .B(G898), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n490), .B(KEYINPUT93), .Z(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n437), .A2(new_n442), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G101), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT79), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT3), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n444), .A4(G104), .ZN(new_n498));
  INV_X1    g312(.A(G104), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n499), .A2(KEYINPUT79), .A3(G107), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT3), .B1(new_n499), .B2(G107), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n495), .B(new_n498), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n499), .A2(G107), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n444), .A2(G104), .ZN(new_n504));
  OAI21_X1  g318(.A(G101), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT10), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n235), .A2(new_n240), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n215), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n510));
  INV_X1    g324(.A(new_n221), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n387), .B2(G146), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n233), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n502), .A2(new_n505), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n260), .A2(new_n261), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G101), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(KEYINPUT4), .A3(new_n502), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n512), .A2(new_n254), .B1(new_n238), .B2(new_n257), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT4), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n522), .A3(G101), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n509), .A2(new_n516), .A3(new_n517), .A4(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G110), .B(G140), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n189), .A2(G227), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n526), .B(new_n527), .Z(new_n528));
  NAND3_X1  g342(.A1(new_n239), .A2(new_n233), .A3(new_n506), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n517), .B1(new_n515), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(KEYINPUT12), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n532), .B(new_n517), .C1(new_n515), .C2(new_n529), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n525), .B(new_n528), .C1(new_n531), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n535));
  INV_X1    g349(.A(new_n517), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n514), .A2(new_n228), .A3(new_n234), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n231), .A2(new_n221), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT1), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n382), .B2(new_n220), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n540), .B2(new_n215), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n506), .B1(new_n541), .B2(new_n233), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n536), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n532), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n530), .A2(KEYINPUT12), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT80), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n525), .A4(new_n528), .ZN(new_n548));
  INV_X1    g362(.A(new_n528), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n520), .A2(new_n523), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n550), .A2(new_n521), .B1(new_n507), .B2(new_n515), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n517), .B1(new_n551), .B2(new_n509), .ZN(new_n552));
  INV_X1    g366(.A(new_n525), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n535), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G469), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n311), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n438), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n546), .A2(new_n525), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n549), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n516), .A2(new_n524), .ZN(new_n562));
  INV_X1    g376(.A(new_n509), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n536), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n525), .A3(new_n528), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(G469), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n557), .A2(new_n559), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G221), .B1(new_n473), .B2(G902), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G214), .B1(G237), .B2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n550), .A2(new_n212), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT5), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n205), .B2(new_n207), .ZN(new_n573));
  OAI21_X1  g387(.A(G113), .B1(new_n202), .B2(KEYINPUT5), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n211), .B(new_n514), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(G110), .B(G122), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT81), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n577), .B(KEYINPUT81), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n581), .A3(new_n575), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(KEYINPUT6), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n206), .A2(KEYINPUT68), .ZN(new_n584));
  AOI211_X1 g398(.A(new_n204), .B(new_n201), .C1(new_n199), .C2(new_n196), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT5), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n574), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n210), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n588), .A2(new_n514), .B1(new_n550), .B2(new_n212), .ZN(new_n589));
  OR3_X1    g403(.A1(new_n589), .A2(KEYINPUT6), .A3(new_n581), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n521), .A2(G125), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n329), .B1(new_n228), .B2(new_n234), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G224), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(G953), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n593), .B(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n583), .A2(new_n590), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(KEYINPUT7), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n591), .A2(new_n592), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(G125), .B1(new_n239), .B2(new_n233), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n258), .A2(G125), .A3(new_n255), .ZN(new_n602));
  OAI211_X1 g416(.A(KEYINPUT7), .B(new_n596), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n582), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n210), .B(new_n514), .C1(new_n586), .C2(new_n587), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n581), .A2(KEYINPUT8), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT8), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n579), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n206), .A2(KEYINPUT5), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n210), .B1(new_n587), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n609), .B1(new_n611), .B2(new_n506), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT82), .B1(new_n605), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n588), .A2(new_n506), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT82), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n587), .A2(new_n610), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n211), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(new_n514), .B1(new_n606), .B2(new_n608), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n604), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(G210), .B1(G237), .B2(G902), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n598), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n598), .B2(new_n621), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n570), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n569), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n373), .A2(new_n494), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G101), .ZN(G3));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n285), .B2(new_n319), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n293), .A2(KEYINPUT94), .A3(new_n311), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n632), .A2(G472), .B1(new_n286), .B2(new_n293), .ZN(new_n633));
  INV_X1    g447(.A(new_n569), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n372), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n477), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT96), .B(G478), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n639));
  AND2_X1   g453(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n640));
  OR4_X1    g454(.A1(new_n475), .A2(new_n476), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(KEYINPUT95), .B(KEYINPUT33), .C1(new_n475), .C2(new_n476), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n319), .A2(new_n478), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n437), .B2(new_n442), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n625), .A2(new_n492), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n635), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT34), .B(G104), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  AOI21_X1  g465(.A(new_n482), .B1(new_n441), .B2(G475), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n425), .A2(new_n435), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n436), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n653), .B1(new_n425), .B2(new_n435), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n647), .B(new_n652), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n425), .A2(new_n435), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT97), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n436), .A3(new_n654), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n662), .A2(KEYINPUT98), .A3(new_n647), .A4(new_n652), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n635), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT35), .B(G107), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  OAI21_X1  g480(.A(new_n346), .B1(KEYINPUT36), .B2(new_n353), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n362), .A2(new_n334), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n667), .A2(new_n369), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n358), .B(new_n311), .C1(new_n363), .C2(new_n364), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n317), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n357), .A2(new_n358), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT99), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n670), .B1(new_n359), .B2(new_n366), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n633), .A2(new_n494), .A3(new_n626), .A4(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  NAND3_X1  g497(.A1(new_n319), .A2(G953), .A3(new_n484), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n486), .B1(G900), .B2(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n652), .B(new_n685), .C1(new_n655), .C2(new_n656), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n678), .B1(new_n367), .B2(new_n671), .ZN(new_n688));
  AOI211_X1 g502(.A(KEYINPUT99), .B(new_n670), .C1(new_n359), .C2(new_n366), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n625), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n288), .A2(new_n294), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n305), .A2(new_n312), .ZN(new_n693));
  INV_X1    g507(.A(new_n304), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n314), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n634), .B(new_n691), .C1(new_n692), .C2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n687), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XNOR2_X1  g513(.A(new_n685), .B(KEYINPUT39), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n634), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n279), .A2(new_n194), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n193), .B1(new_n306), .B2(new_n307), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n438), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G472), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n288), .A2(new_n294), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n482), .B1(new_n437), .B2(new_n442), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n623), .A2(new_n624), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n570), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n712), .A2(new_n713), .A3(new_n680), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n702), .A2(new_n708), .A3(new_n709), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n382), .ZN(G45));
  AND2_X1   g530(.A1(new_n646), .A2(new_n685), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n697), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  NAND2_X1  g533(.A1(new_n555), .A2(new_n311), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n568), .A3(new_n557), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n315), .A2(new_n372), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n648), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT41), .B(G113), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  AOI21_X1  g541(.A(new_n724), .B1(new_n659), .B2(new_n663), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n198), .ZN(G18));
  NAND4_X1  g543(.A1(new_n494), .A2(new_n315), .A3(new_n691), .A4(new_n723), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  AOI211_X1 g545(.A(new_n482), .B(new_n625), .C1(new_n437), .C2(new_n442), .ZN(new_n732));
  OAI21_X1  g546(.A(G472), .B1(new_n285), .B2(new_n319), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n371), .A2(KEYINPUT102), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n367), .A2(new_n735), .A3(new_n370), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n194), .B1(new_n267), .B2(new_n308), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n281), .B2(new_n284), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT101), .B1(new_n739), .B2(new_n287), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT101), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n291), .A2(new_n292), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n741), .B(new_n286), .C1(new_n742), .C2(new_n738), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n733), .A2(new_n737), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n722), .A2(new_n492), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n732), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NAND2_X1  g561(.A1(new_n437), .A2(new_n442), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n722), .A2(new_n625), .ZN(new_n749));
  INV_X1    g563(.A(new_n645), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n685), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n740), .A2(new_n743), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(KEYINPUT103), .A3(new_n680), .A4(new_n733), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n733), .A2(new_n740), .A3(new_n743), .A4(new_n680), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT103), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n751), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n329), .ZN(G27));
  NAND2_X1  g572(.A1(new_n598), .A2(new_n621), .ZN(new_n759));
  INV_X1    g573(.A(new_n622), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n598), .A2(new_n621), .A3(new_n622), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n568), .A3(new_n570), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n565), .A2(KEYINPUT104), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT104), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n564), .A2(new_n765), .A3(new_n525), .A4(new_n528), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n561), .A2(new_n764), .A3(G469), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n557), .A2(new_n559), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT105), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n557), .A2(KEYINPUT105), .A3(new_n559), .A4(new_n767), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n763), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n315), .A2(new_n772), .A3(new_n372), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n717), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n315), .A2(new_n772), .A3(new_n372), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n646), .A2(new_n685), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT106), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n772), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT32), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n285), .B2(new_n287), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n294), .C1(new_n314), .C2(new_n313), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n737), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(KEYINPUT42), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NOR2_X1   g604(.A1(new_n776), .A2(new_n686), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n242), .ZN(G36));
  OR3_X1    g606(.A1(new_n748), .A2(KEYINPUT43), .A3(new_n645), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT43), .B1(new_n748), .B2(new_n645), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n633), .A2(new_n690), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n561), .A2(new_n565), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n561), .A2(new_n764), .A3(KEYINPUT45), .A4(new_n766), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT107), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  OAI221_X1 g617(.A(G469), .B1(KEYINPUT45), .B2(new_n799), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n559), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT46), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n804), .A2(KEYINPUT46), .A3(new_n559), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n557), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n568), .A3(new_n700), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n797), .B1(new_n795), .B2(new_n796), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n623), .A2(new_n624), .A3(new_n713), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n798), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(KEYINPUT108), .B(G137), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n813), .B(new_n814), .ZN(G39));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n809), .A2(KEYINPUT47), .A3(new_n568), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT47), .B1(new_n809), .B2(new_n568), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n812), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n777), .A2(new_n372), .A3(new_n315), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n816), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n819), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n817), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n822), .B(KEYINPUT109), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(KEYINPUT110), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G140), .ZN(G42));
  NAND2_X1  g645(.A1(new_n721), .A2(new_n557), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT111), .Z(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT49), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n748), .A3(new_n645), .ZN(new_n835));
  INV_X1    g649(.A(new_n708), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n737), .A2(new_n568), .A3(new_n570), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n712), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n480), .A2(new_n481), .A3(new_n685), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n441), .B2(G475), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n812), .A2(new_n680), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n315), .A2(new_n843), .A3(new_n634), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n655), .A2(new_n656), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n812), .A2(new_n680), .A3(new_n842), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n569), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n662), .A3(KEYINPUT112), .A4(new_n315), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n791), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n753), .A2(new_n756), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n782), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n746), .B(new_n730), .C1(new_n648), .C2(new_n724), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n728), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n748), .A2(new_n482), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n647), .B1(new_n857), .B2(new_n646), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n627), .B(new_n681), .C1(new_n635), .C2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n854), .A2(new_n789), .A3(new_n856), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n696), .B1(new_n686), .B2(new_n777), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n757), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n770), .A2(new_n771), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n677), .A2(new_n568), .A3(new_n685), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n708), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n625), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n748), .A2(new_n483), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n757), .A2(new_n862), .A3(new_n872), .A4(new_n869), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n839), .B1(new_n861), .B2(new_n874), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n786), .A2(new_n777), .A3(new_n781), .A4(new_n779), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n776), .A2(new_n777), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT42), .B1(new_n877), .B2(new_n774), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n878), .B2(new_n778), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n659), .A2(new_n663), .ZN(new_n880));
  INV_X1    g694(.A(new_n724), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n315), .A2(new_n691), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n723), .A2(new_n437), .A3(new_n442), .A4(new_n493), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n724), .A2(new_n648), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n732), .A2(new_n744), .A3(new_n745), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT114), .B1(new_n879), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n751), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n852), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(new_n698), .A3(new_n718), .A4(new_n870), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n872), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n863), .A2(KEYINPUT52), .A3(new_n870), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n850), .A2(new_n853), .A3(new_n851), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n896), .A2(new_n839), .A3(new_n859), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT114), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n789), .A2(new_n856), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n889), .A2(new_n895), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n875), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT113), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n875), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n895), .A2(new_n897), .A3(new_n789), .A4(new_n856), .ZN(new_n905));
  OAI211_X1 g719(.A(KEYINPUT113), .B(new_n839), .C1(new_n861), .C2(new_n874), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n902), .B1(new_n907), .B2(KEYINPUT54), .ZN(new_n908));
  NOR4_X1   g722(.A1(new_n763), .A2(new_n832), .A3(new_n371), .A4(new_n486), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n646), .A3(new_n836), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(G952), .A3(new_n189), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n487), .A2(new_n793), .A3(new_n744), .A4(new_n794), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n749), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n795), .A2(new_n486), .A3(new_n832), .A4(new_n763), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n787), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(KEYINPUT48), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(KEYINPUT48), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n833), .A2(new_n568), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n812), .B(new_n912), .C1(new_n827), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n909), .A2(new_n836), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n921), .A2(new_n748), .A3(new_n750), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n914), .B2(new_n852), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n712), .A2(new_n713), .A3(new_n723), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT115), .Z(new_n925));
  AOI21_X1  g739(.A(KEYINPUT50), .B1(new_n925), .B2(new_n912), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n925), .A2(new_n912), .A3(KEYINPUT50), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n920), .B(new_n923), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT51), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n918), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n927), .B2(new_n926), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n923), .B(KEYINPUT116), .C1(new_n927), .C2(new_n926), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n933), .A2(KEYINPUT51), .A3(new_n934), .A4(new_n920), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n908), .A2(new_n936), .A3(KEYINPUT117), .ZN(new_n937));
  NOR2_X1   g751(.A1(G952), .A2(G953), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT118), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT117), .B1(new_n908), .B2(new_n936), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n838), .B1(new_n940), .B2(new_n941), .ZN(G75));
  INV_X1    g756(.A(KEYINPUT119), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n583), .A2(new_n590), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(new_n597), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT55), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n901), .A2(new_n319), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n622), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n943), .B(new_n946), .C1(new_n948), .C2(KEYINPUT56), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n189), .A2(G952), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n948), .A2(KEYINPUT56), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n946), .B1(new_n953), .B2(new_n943), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n943), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G51));
  NOR2_X1   g770(.A1(new_n947), .A2(new_n804), .ZN(new_n957));
  INV_X1    g771(.A(new_n555), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n901), .B(KEYINPUT54), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n558), .B(KEYINPUT57), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n957), .B1(new_n962), .B2(KEYINPUT120), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT54), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n901), .B(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n555), .B1(new_n965), .B2(new_n960), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n950), .B1(new_n963), .B2(new_n968), .ZN(G54));
  AND4_X1   g783(.A1(KEYINPUT58), .A2(new_n901), .A3(G475), .A4(new_n319), .ZN(new_n970));
  INV_X1    g784(.A(new_n422), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n951), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n971), .B2(new_n970), .ZN(G60));
  INV_X1    g787(.A(new_n643), .ZN(new_n974));
  NAND2_X1  g788(.A1(G478), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT59), .Z(new_n976));
  OR2_X1    g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n951), .B1(new_n965), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n908), .A2(new_n976), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n974), .ZN(G63));
  INV_X1    g794(.A(KEYINPUT121), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n981), .A2(KEYINPUT61), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT122), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT60), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n875), .B2(new_n900), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n951), .B1(new_n989), .B2(new_n368), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n667), .A2(new_n669), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n901), .A2(new_n991), .A3(new_n987), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n984), .B(new_n985), .C1(new_n990), .C2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n901), .A2(new_n991), .A3(new_n987), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n995), .B(new_n951), .C1(new_n368), .C2(new_n989), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n984), .B1(new_n996), .B2(new_n985), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n983), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n985), .B1(new_n990), .B2(new_n992), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(KEYINPUT122), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n982), .A3(new_n993), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n998), .A2(new_n1001), .ZN(G66));
  OAI21_X1  g816(.A(G953), .B1(new_n489), .B2(new_n594), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT123), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n888), .A2(new_n859), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n944), .B1(G898), .B2(new_n189), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G69));
  NOR2_X1   g822(.A1(new_n786), .A2(new_n868), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n791), .B1(new_n810), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n813), .A2(new_n1010), .A3(new_n789), .A4(new_n863), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(G953), .B1(new_n1012), .B2(new_n830), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n189), .A2(G900), .ZN(new_n1014));
  OAI21_X1  g828(.A(KEYINPUT125), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n825), .A2(new_n829), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n189), .B1(new_n1016), .B2(new_n1011), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT125), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1014), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n276), .A2(new_n277), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(new_n401), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n701), .A2(new_n821), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n373), .B(new_n1025), .C1(new_n646), .C2(new_n857), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n813), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT124), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n813), .A2(KEYINPUT124), .A3(new_n1026), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n715), .A2(new_n863), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT62), .Z(new_n1033));
  AND3_X1   g847(.A1(new_n1031), .A2(new_n830), .A3(new_n1033), .ZN(new_n1034));
  OR3_X1    g848(.A1(new_n1034), .A2(G953), .A3(new_n1023), .ZN(new_n1035));
  NAND2_X1  g849(.A1(G227), .A2(G900), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(G953), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1024), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n1021), .A2(G953), .A3(new_n1036), .A4(new_n1023), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT63), .Z(new_n1042));
  NAND2_X1  g856(.A1(new_n295), .A2(new_n193), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n703), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n907), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1012), .A2(new_n830), .A3(new_n1005), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n1046), .A2(new_n1042), .ZN(new_n1047));
  XNOR2_X1  g861(.A(new_n295), .B(KEYINPUT126), .ZN(new_n1048));
  OR2_X1    g862(.A1(new_n1048), .A2(new_n194), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1045), .B(new_n951), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1048), .A2(new_n194), .ZN(new_n1051));
  NAND4_X1  g865(.A1(new_n1031), .A2(new_n830), .A3(new_n1005), .A4(new_n1033), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1051), .B1(new_n1052), .B2(new_n1042), .ZN(new_n1053));
  OR2_X1    g867(.A1(new_n1053), .A2(KEYINPUT127), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1053), .A2(KEYINPUT127), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1050), .B1(new_n1054), .B2(new_n1055), .ZN(G57));
endmodule


