

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U547 ( .A1(G651), .A2(G543), .ZN(n641) );
  NOR2_X1 U548 ( .A1(n720), .A2(n999), .ZN(n680) );
  NOR2_X1 U549 ( .A1(n737), .A2(n736), .ZN(n739) );
  AND2_X1 U550 ( .A1(n728), .A2(n727), .ZN(n729) );
  INV_X1 U551 ( .A(G2104), .ZN(n513) );
  INV_X1 U552 ( .A(G2105), .ZN(n514) );
  INV_X1 U553 ( .A(n969), .ZN(n681) );
  AND2_X1 U554 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U555 ( .A1(n684), .A2(n683), .ZN(n686) );
  XOR2_X1 U556 ( .A(n720), .B(KEYINPUT96), .Z(n707) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n704) );
  AND2_X1 U558 ( .A1(n735), .A2(n734), .ZN(n736) );
  INV_X1 U559 ( .A(KEYINPUT101), .ZN(n738) );
  INV_X1 U560 ( .A(KEYINPUT32), .ZN(n731) );
  XNOR2_X1 U561 ( .A(n731), .B(KEYINPUT103), .ZN(n732) );
  XNOR2_X1 U562 ( .A(n733), .B(n732), .ZN(n792) );
  XNOR2_X1 U563 ( .A(n517), .B(KEYINPUT65), .ZN(n546) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n759) );
  INV_X1 U565 ( .A(KEYINPUT105), .ZN(n808) );
  NAND2_X1 U566 ( .A1(n514), .A2(n513), .ZN(n515) );
  NOR2_X1 U567 ( .A1(G651), .A2(n632), .ZN(n639) );
  XNOR2_X2 U568 ( .A(n515), .B(KEYINPUT17), .ZN(n882) );
  NAND2_X1 U569 ( .A1(G138), .A2(n882), .ZN(n520) );
  INV_X1 U570 ( .A(G2105), .ZN(n516) );
  NAND2_X1 U571 ( .A1(n516), .A2(G2104), .ZN(n517) );
  INV_X1 U572 ( .A(n546), .ZN(n518) );
  INV_X1 U573 ( .A(n518), .ZN(n880) );
  NAND2_X1 U574 ( .A1(G102), .A2(n880), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n520), .A2(n519), .ZN(n525) );
  NOR2_X2 U576 ( .A1(G2104), .A2(n514), .ZN(n875) );
  NAND2_X1 U577 ( .A1(G126), .A2(n875), .ZN(n523) );
  NAND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XNOR2_X2 U579 ( .A(n521), .B(KEYINPUT67), .ZN(n876) );
  NAND2_X1 U580 ( .A1(G114), .A2(n876), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U583 ( .A(KEYINPUT89), .B(n526), .Z(G164) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  INV_X1 U585 ( .A(G651), .ZN(n528) );
  NOR2_X1 U586 ( .A1(n632), .A2(n528), .ZN(n644) );
  NAND2_X1 U587 ( .A1(G78), .A2(n644), .ZN(n527) );
  XOR2_X1 U588 ( .A(KEYINPUT70), .B(n527), .Z(n534) );
  NOR2_X1 U589 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n529), .Z(n640) );
  NAND2_X1 U591 ( .A1(G65), .A2(n640), .ZN(n531) );
  NAND2_X1 U592 ( .A1(G53), .A2(n639), .ZN(n530) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U594 ( .A(KEYINPUT71), .B(n532), .Z(n533) );
  NOR2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n641), .A2(G91), .ZN(n535) );
  NAND2_X1 U597 ( .A1(n536), .A2(n535), .ZN(G299) );
  NAND2_X1 U598 ( .A1(G85), .A2(n641), .ZN(n538) );
  NAND2_X1 U599 ( .A1(G72), .A2(n644), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G60), .A2(n640), .ZN(n540) );
  NAND2_X1 U602 ( .A1(G47), .A2(n639), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  OR2_X1 U604 ( .A1(n542), .A2(n541), .ZN(G290) );
  NAND2_X1 U605 ( .A1(G113), .A2(n876), .ZN(n544) );
  NAND2_X1 U606 ( .A1(G137), .A2(n882), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n545), .B(KEYINPUT68), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G101), .A2(n546), .ZN(n547) );
  XNOR2_X1 U610 ( .A(KEYINPUT66), .B(n547), .ZN(n549) );
  INV_X1 U611 ( .A(KEYINPUT23), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G125), .A2(n875), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT64), .ZN(n677) );
  BUF_X1 U617 ( .A(n677), .Z(G160) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  NAND2_X1 U621 ( .A1(G64), .A2(n640), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G52), .A2(n639), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n641), .A2(G90), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT69), .B(n557), .Z(n559) );
  NAND2_X1 U626 ( .A1(n644), .A2(G77), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n560), .Z(n561) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U630 ( .A1(G89), .A2(n641), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT4), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G76), .A2(n644), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G63), .A2(n640), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G51), .A2(n639), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U643 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n575) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U645 ( .A(n575), .B(n574), .ZN(G223) );
  INV_X1 U646 ( .A(G223), .ZN(n827) );
  NAND2_X1 U647 ( .A1(n827), .A2(G567), .ZN(n576) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U649 ( .A1(G56), .A2(n640), .ZN(n577) );
  XOR2_X1 U650 ( .A(KEYINPUT14), .B(n577), .Z(n584) );
  NAND2_X1 U651 ( .A1(G81), .A2(n641), .ZN(n578) );
  XNOR2_X1 U652 ( .A(n578), .B(KEYINPUT12), .ZN(n579) );
  XNOR2_X1 U653 ( .A(n579), .B(KEYINPUT74), .ZN(n581) );
  NAND2_X1 U654 ( .A1(G68), .A2(n644), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U656 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  NOR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n639), .A2(G43), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n586), .A2(n585), .ZN(n969) );
  INV_X1 U660 ( .A(G860), .ZN(n599) );
  OR2_X1 U661 ( .A1(n969), .A2(n599), .ZN(G153) );
  INV_X1 U662 ( .A(G171), .ZN(G301) );
  NAND2_X1 U663 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G54), .A2(n639), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G66), .A2(n640), .ZN(n588) );
  NAND2_X1 U666 ( .A1(G79), .A2(n644), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U668 ( .A1(G92), .A2(n641), .ZN(n589) );
  XNOR2_X1 U669 ( .A(KEYINPUT75), .B(n589), .ZN(n590) );
  NOR2_X1 U670 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U672 ( .A(n594), .B(KEYINPUT15), .ZN(n984) );
  OR2_X1 U673 ( .A1(n984), .A2(G868), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(G284) );
  INV_X1 U675 ( .A(G868), .ZN(n657) );
  NOR2_X1 U676 ( .A1(G286), .A2(n657), .ZN(n598) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U678 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n600), .A2(n984), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n969), .ZN(n604) );
  NAND2_X1 U683 ( .A1(G868), .A2(n984), .ZN(n602) );
  NOR2_X1 U684 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U686 ( .A(KEYINPUT77), .B(n605), .Z(G282) );
  NAND2_X1 U687 ( .A1(G111), .A2(n876), .ZN(n606) );
  XNOR2_X1 U688 ( .A(n606), .B(KEYINPUT78), .ZN(n609) );
  NAND2_X1 U689 ( .A1(G123), .A2(n875), .ZN(n607) );
  XNOR2_X1 U690 ( .A(n607), .B(KEYINPUT18), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U692 ( .A1(G135), .A2(n882), .ZN(n611) );
  NAND2_X1 U693 ( .A1(G99), .A2(n880), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n932) );
  XNOR2_X1 U696 ( .A(n932), .B(G2096), .ZN(n615) );
  INV_X1 U697 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G61), .A2(n640), .ZN(n617) );
  NAND2_X1 U700 ( .A1(G86), .A2(n641), .ZN(n616) );
  NAND2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n644), .A2(G73), .ZN(n618) );
  XOR2_X1 U703 ( .A(KEYINPUT2), .B(n618), .Z(n619) );
  NOR2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n639), .A2(G48), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n622), .A2(n621), .ZN(G305) );
  NAND2_X1 U707 ( .A1(G88), .A2(n641), .ZN(n624) );
  NAND2_X1 U708 ( .A1(G75), .A2(n644), .ZN(n623) );
  NAND2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G62), .A2(n640), .ZN(n626) );
  NAND2_X1 U711 ( .A1(G50), .A2(n639), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U713 ( .A1(n628), .A2(n627), .ZN(G166) );
  NAND2_X1 U714 ( .A1(G49), .A2(n639), .ZN(n630) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U717 ( .A1(n640), .A2(n631), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n632), .A2(G87), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(G288) );
  XNOR2_X1 U720 ( .A(n969), .B(KEYINPUT79), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n984), .A2(G559), .ZN(n635) );
  XOR2_X1 U722 ( .A(n636), .B(n635), .Z(n915) );
  XNOR2_X1 U723 ( .A(KEYINPUT19), .B(KEYINPUT83), .ZN(n638) );
  XNOR2_X1 U724 ( .A(G305), .B(KEYINPUT82), .ZN(n637) );
  XNOR2_X1 U725 ( .A(n638), .B(n637), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G55), .A2(n639), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G67), .A2(n640), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G93), .A2(n641), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n644), .A2(G80), .ZN(n645) );
  XOR2_X1 U731 ( .A(KEYINPUT80), .B(n645), .Z(n646) );
  NOR2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U734 ( .A(n650), .B(KEYINPUT81), .ZN(n916) );
  XOR2_X1 U735 ( .A(n651), .B(n916), .Z(n653) );
  INV_X1 U736 ( .A(G299), .ZN(n973) );
  XNOR2_X1 U737 ( .A(n973), .B(G166), .ZN(n652) );
  XNOR2_X1 U738 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U739 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U740 ( .A(n655), .B(G288), .ZN(n894) );
  XOR2_X1 U741 ( .A(n915), .B(n894), .Z(n656) );
  NAND2_X1 U742 ( .A1(n656), .A2(G868), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n916), .A2(n657), .ZN(n658) );
  NAND2_X1 U744 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U745 ( .A(KEYINPUT84), .B(n660), .Z(G295) );
  NAND2_X1 U746 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XNOR2_X1 U747 ( .A(n661), .B(KEYINPUT20), .ZN(n662) );
  XNOR2_X1 U748 ( .A(n662), .B(KEYINPUT85), .ZN(n663) );
  NAND2_X1 U749 ( .A1(n663), .A2(G2090), .ZN(n664) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n665), .A2(G2072), .ZN(n666) );
  XNOR2_X1 U752 ( .A(KEYINPUT86), .B(n666), .ZN(G158) );
  XOR2_X1 U753 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G108), .A2(G120), .ZN(n667) );
  NOR2_X1 U756 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U757 ( .A1(G69), .A2(n668), .ZN(n913) );
  NAND2_X1 U758 ( .A1(G567), .A2(n913), .ZN(n673) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U761 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U762 ( .A1(G96), .A2(n671), .ZN(n914) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n914), .ZN(n672) );
  NAND2_X1 U764 ( .A1(n673), .A2(n672), .ZN(n831) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n674) );
  XOR2_X1 U766 ( .A(KEYINPUT87), .B(n674), .Z(n675) );
  NOR2_X1 U767 ( .A1(n831), .A2(n675), .ZN(n676) );
  XNOR2_X1 U768 ( .A(KEYINPUT88), .B(n676), .ZN(n830) );
  NAND2_X1 U769 ( .A1(G36), .A2(n830), .ZN(G176) );
  XOR2_X1 U770 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NAND2_X1 U771 ( .A1(G40), .A2(n677), .ZN(n758) );
  INV_X1 U772 ( .A(n758), .ZN(n678) );
  NAND2_X2 U773 ( .A1(n759), .A2(n678), .ZN(n720) );
  INV_X1 U774 ( .A(G1996), .ZN(n999) );
  INV_X1 U775 ( .A(KEYINPUT26), .ZN(n679) );
  XNOR2_X1 U776 ( .A(n680), .B(n679), .ZN(n684) );
  NAND2_X1 U777 ( .A1(n720), .A2(G1341), .ZN(n682) );
  NOR2_X1 U778 ( .A1(n686), .A2(n984), .ZN(n685) );
  XNOR2_X1 U779 ( .A(n685), .B(KEYINPUT99), .ZN(n692) );
  NAND2_X1 U780 ( .A1(n686), .A2(n984), .ZN(n690) );
  NAND2_X1 U781 ( .A1(G2067), .A2(n707), .ZN(n688) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n720), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U786 ( .A(n693), .B(KEYINPUT100), .ZN(n698) );
  NAND2_X1 U787 ( .A1(G2072), .A2(n707), .ZN(n694) );
  XNOR2_X1 U788 ( .A(n694), .B(KEYINPUT27), .ZN(n696) );
  XOR2_X1 U789 ( .A(KEYINPUT98), .B(G1956), .Z(n949) );
  NOR2_X1 U790 ( .A1(n707), .A2(n949), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n699), .A2(n973), .ZN(n697) );
  NAND2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n699), .A2(n973), .ZN(n700) );
  XNOR2_X1 U795 ( .A(n700), .B(KEYINPUT28), .ZN(n701) );
  INV_X1 U796 ( .A(n701), .ZN(n702) );
  NAND2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n705) );
  XNOR2_X1 U798 ( .A(n705), .B(n704), .ZN(n712) );
  XOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .Z(n706) );
  XNOR2_X1 U800 ( .A(KEYINPUT97), .B(n706), .ZN(n1001) );
  NAND2_X1 U801 ( .A1(n707), .A2(n1001), .ZN(n710) );
  INV_X1 U802 ( .A(G1961), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n708), .A2(n720), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n710), .A2(n709), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n716), .A2(G171), .ZN(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n735) );
  NOR2_X1 U807 ( .A1(G2084), .A2(n720), .ZN(n740) );
  NAND2_X1 U808 ( .A1(G8), .A2(n720), .ZN(n800) );
  NOR2_X1 U809 ( .A1(G1966), .A2(n800), .ZN(n737) );
  NOR2_X1 U810 ( .A1(n740), .A2(n737), .ZN(n713) );
  NAND2_X1 U811 ( .A1(G8), .A2(n713), .ZN(n714) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n714), .ZN(n715) );
  NOR2_X1 U813 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U814 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U815 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U816 ( .A(KEYINPUT31), .B(n719), .Z(n734) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n800), .ZN(n722) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U819 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U820 ( .A1(n723), .A2(G303), .ZN(n725) );
  AND2_X1 U821 ( .A1(n734), .A2(n725), .ZN(n724) );
  NAND2_X1 U822 ( .A1(n735), .A2(n724), .ZN(n728) );
  INV_X1 U823 ( .A(n725), .ZN(n726) );
  OR2_X1 U824 ( .A1(n726), .A2(G286), .ZN(n727) );
  XNOR2_X1 U825 ( .A(n729), .B(KEYINPUT102), .ZN(n730) );
  NAND2_X1 U826 ( .A1(n730), .A2(G8), .ZN(n733) );
  XNOR2_X1 U827 ( .A(n739), .B(n738), .ZN(n743) );
  NAND2_X1 U828 ( .A1(G8), .A2(n740), .ZN(n741) );
  XOR2_X1 U829 ( .A(KEYINPUT95), .B(n741), .Z(n742) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n791) );
  INV_X1 U831 ( .A(KEYINPUT33), .ZN(n744) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NAND2_X1 U833 ( .A1(n744), .A2(n976), .ZN(n745) );
  INV_X1 U834 ( .A(n800), .ZN(n751) );
  NOR2_X1 U835 ( .A1(n745), .A2(n800), .ZN(n747) );
  AND2_X1 U836 ( .A1(n791), .A2(n747), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n792), .A2(n746), .ZN(n756) );
  INV_X1 U838 ( .A(n747), .ZN(n750) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n975) );
  NOR2_X1 U840 ( .A1(G303), .A2(G1971), .ZN(n748) );
  NOR2_X1 U841 ( .A1(n975), .A2(n748), .ZN(n749) );
  OR2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n975), .A2(n751), .ZN(n752) );
  NAND2_X1 U844 ( .A1(n752), .A2(KEYINPUT33), .ZN(n753) );
  AND2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U847 ( .A(n757), .B(KEYINPUT104), .ZN(n790) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n987) );
  NOR2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n822) );
  XNOR2_X1 U850 ( .A(KEYINPUT37), .B(G2067), .ZN(n819) );
  NAND2_X1 U851 ( .A1(G140), .A2(n882), .ZN(n761) );
  NAND2_X1 U852 ( .A1(G104), .A2(n880), .ZN(n760) );
  NAND2_X1 U853 ( .A1(n761), .A2(n760), .ZN(n763) );
  XOR2_X1 U854 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n762) );
  XNOR2_X1 U855 ( .A(n763), .B(n762), .ZN(n768) );
  NAND2_X1 U856 ( .A1(G128), .A2(n875), .ZN(n765) );
  NAND2_X1 U857 ( .A1(G116), .A2(n876), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U859 ( .A(KEYINPUT35), .B(n766), .Z(n767) );
  NOR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U861 ( .A(KEYINPUT36), .B(n769), .ZN(n858) );
  NOR2_X1 U862 ( .A1(n819), .A2(n858), .ZN(n931) );
  NAND2_X1 U863 ( .A1(n822), .A2(n931), .ZN(n817) );
  NAND2_X1 U864 ( .A1(G119), .A2(n875), .ZN(n771) );
  NAND2_X1 U865 ( .A1(G107), .A2(n876), .ZN(n770) );
  NAND2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U867 ( .A1(n880), .A2(G95), .ZN(n772) );
  XOR2_X1 U868 ( .A(KEYINPUT92), .B(n772), .Z(n773) );
  NOR2_X1 U869 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n882), .A2(G131), .ZN(n775) );
  NAND2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n870) );
  NAND2_X1 U872 ( .A1(n870), .A2(G1991), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G129), .A2(n875), .ZN(n778) );
  NAND2_X1 U874 ( .A1(G117), .A2(n876), .ZN(n777) );
  NAND2_X1 U875 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n880), .A2(G105), .ZN(n779) );
  XOR2_X1 U877 ( .A(KEYINPUT38), .B(n779), .Z(n780) );
  NOR2_X1 U878 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U879 ( .A(KEYINPUT93), .B(n782), .Z(n784) );
  NAND2_X1 U880 ( .A1(n882), .A2(G141), .ZN(n783) );
  NAND2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n891) );
  NAND2_X1 U882 ( .A1(n891), .A2(G1996), .ZN(n785) );
  AND2_X1 U883 ( .A1(n786), .A2(n785), .ZN(n928) );
  XOR2_X1 U884 ( .A(n822), .B(KEYINPUT94), .Z(n787) );
  NOR2_X1 U885 ( .A1(n928), .A2(n787), .ZN(n814) );
  INV_X1 U886 ( .A(n814), .ZN(n788) );
  AND2_X1 U887 ( .A1(n817), .A2(n788), .ZN(n805) );
  AND2_X1 U888 ( .A1(n987), .A2(n805), .ZN(n789) );
  NAND2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n807) );
  NAND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n799) );
  NOR2_X1 U891 ( .A1(G2090), .A2(G303), .ZN(n793) );
  NAND2_X1 U892 ( .A1(G8), .A2(n793), .ZN(n797) );
  NOR2_X1 U893 ( .A1(G1981), .A2(G305), .ZN(n794) );
  XOR2_X1 U894 ( .A(n794), .B(KEYINPUT24), .Z(n795) );
  NOR2_X1 U895 ( .A1(n800), .A2(n795), .ZN(n801) );
  INV_X1 U896 ( .A(n801), .ZN(n796) );
  AND2_X1 U897 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n803) );
  OR2_X1 U899 ( .A1(n801), .A2(n800), .ZN(n802) );
  AND2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n809), .B(n808), .ZN(n811) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n986) );
  NAND2_X1 U905 ( .A1(n986), .A2(n822), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n825) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n891), .ZN(n924) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n870), .ZN(n933) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n933), .A2(n812), .ZN(n813) );
  NOR2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n924), .A2(n815), .ZN(n816) );
  XNOR2_X1 U913 ( .A(KEYINPUT39), .B(n816), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n858), .A2(n819), .ZN(n820) );
  XNOR2_X1 U916 ( .A(n820), .B(KEYINPUT106), .ZN(n938) );
  NAND2_X1 U917 ( .A1(n821), .A2(n938), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U923 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G188) );
  XNOR2_X1 U926 ( .A(KEYINPUT107), .B(n831), .ZN(G319) );
  XOR2_X1 U927 ( .A(G2100), .B(G2678), .Z(n833) );
  XNOR2_X1 U928 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U930 ( .A(KEYINPUT42), .B(G2090), .Z(n835) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U933 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U934 ( .A(KEYINPUT43), .B(G2096), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n841) );
  XOR2_X1 U936 ( .A(G2084), .B(G2078), .Z(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U938 ( .A(G1976), .B(G1971), .Z(n843) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1966), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(n844), .B(G2474), .Z(n846) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U944 ( .A(KEYINPUT41), .B(G1981), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1961), .B(G1956), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(G229) );
  NAND2_X1 U948 ( .A1(n875), .A2(G124), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U950 ( .A1(G112), .A2(n876), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G136), .A2(n882), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G100), .A2(n880), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U955 ( .A1(n857), .A2(n856), .ZN(G162) );
  XNOR2_X1 U956 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n858), .B(KEYINPUT48), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n872) );
  NAND2_X1 U959 ( .A1(G127), .A2(n875), .ZN(n862) );
  NAND2_X1 U960 ( .A1(G115), .A2(n876), .ZN(n861) );
  NAND2_X1 U961 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n863), .B(KEYINPUT47), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G139), .A2(n882), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n880), .A2(G103), .ZN(n866) );
  XOR2_X1 U966 ( .A(KEYINPUT112), .B(n866), .Z(n867) );
  NOR2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n919) );
  XOR2_X1 U968 ( .A(n932), .B(n919), .Z(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U970 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U971 ( .A(G164), .B(G162), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n889) );
  NAND2_X1 U973 ( .A1(G130), .A2(n875), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U976 ( .A(KEYINPUT110), .B(n879), .ZN(n887) );
  NAND2_X1 U977 ( .A1(n880), .A2(G106), .ZN(n881) );
  XOR2_X1 U978 ( .A(KEYINPUT111), .B(n881), .Z(n884) );
  NAND2_X1 U979 ( .A1(n882), .A2(G142), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U981 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U982 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U983 ( .A(n889), .B(n888), .Z(n890) );
  XNOR2_X1 U984 ( .A(n890), .B(G160), .ZN(n892) );
  XNOR2_X1 U985 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U986 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U987 ( .A(n969), .B(n894), .ZN(n896) );
  XNOR2_X1 U988 ( .A(G171), .B(n984), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U990 ( .A(G286), .B(n897), .Z(n898) );
  NOR2_X1 U991 ( .A1(G37), .A2(n898), .ZN(G397) );
  XOR2_X1 U992 ( .A(G2451), .B(G2430), .Z(n900) );
  XNOR2_X1 U993 ( .A(G2438), .B(G2443), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n906) );
  XOR2_X1 U995 ( .A(G2435), .B(G2454), .Z(n902) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n904) );
  XOR2_X1 U998 ( .A(G2446), .B(G2427), .Z(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n907), .ZN(n918) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n918), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(G225) );
  XOR2_X1 U1008 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1010 ( .A(G120), .ZN(G236) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G325) );
  INV_X1 U1015 ( .A(G325), .ZN(G261) );
  NOR2_X1 U1016 ( .A1(n915), .A2(G860), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n917), .B(n916), .ZN(G145) );
  INV_X1 U1018 ( .A(n918), .ZN(G401) );
  XOR2_X1 U1019 ( .A(G2072), .B(n919), .Z(n921) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(KEYINPUT50), .B(n922), .ZN(n927) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1025 ( .A(KEYINPUT51), .B(n925), .Z(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n940) );
  XNOR2_X1 U1027 ( .A(G2084), .B(G160), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT115), .B(n936), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1035 ( .A(KEYINPUT52), .B(n941), .Z(n942) );
  NOR2_X1 U1036 ( .A1(KEYINPUT55), .A2(n942), .ZN(n944) );
  INV_X1 U1037 ( .A(G29), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n1028) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G21), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G1961), .B(G5), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n958) );
  XOR2_X1 U1042 ( .A(KEYINPUT126), .B(G4), .Z(n948) );
  XNOR2_X1 U1043 ( .A(G1348), .B(KEYINPUT59), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(n948), .B(n947), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(n949), .B(G20), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G1981), .B(G6), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT60), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n965) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n962) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1060 ( .A(KEYINPUT61), .B(n966), .Z(n967) );
  NOR2_X1 U1061 ( .A1(G16), .A2(n967), .ZN(n1025) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT121), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1064 ( .A(G1341), .B(KEYINPUT124), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(n969), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1961), .B(G301), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n983) );
  XOR2_X1 U1068 ( .A(G1956), .B(n973), .Z(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(G303), .B(G1971), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n978), .B(KEYINPUT122), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT123), .B(n981), .Z(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n993) );
  XOR2_X1 U1076 ( .A(n984), .B(G1348), .Z(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT57), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1084 ( .A(KEYINPUT125), .B(n996), .Z(n1022) );
  XNOR2_X1 U1085 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n1017) );
  XNOR2_X1 U1086 ( .A(G2067), .B(G26), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G33), .B(G2072), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(G32), .B(n999), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(G28), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(G27), .B(n1001), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(KEYINPUT116), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G25), .B(G1991), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT117), .B(n1009), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT53), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(G2084), .B(G34), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1011), .B(KEYINPUT54), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G35), .B(G2090), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(n1017), .B(n1016), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(G29), .B(KEYINPUT119), .Z(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT120), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(G11), .A2(n1023), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(n1026), .B(KEYINPUT127), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1029), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

