//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0005(.A1(G58), .A2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  AND4_X1   g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT66), .B(G244), .Z(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G77), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n215), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n213), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n215), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT65), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n225), .B(new_n231), .C1(new_n224), .C2(new_n223), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT68), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT70), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT70), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n252), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n210), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n203), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(new_n211), .B2(G68), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n254), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT11), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n251), .A2(new_n253), .A3(new_n210), .A4(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n214), .A2(G20), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT71), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(G68), .A3(new_n268), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n271), .B(new_n272), .C1(new_n264), .C2(G68), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(KEYINPUT79), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(KEYINPUT79), .B2(new_n273), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n263), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT14), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT76), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n284), .A3(G274), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(G238), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n279), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n285), .A2(new_n287), .A3(new_n279), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G33), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n292), .A2(new_n294), .A3(G232), .A4(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n292), .A2(new_n294), .A3(G226), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G97), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n278), .B1(new_n291), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n285), .A2(new_n287), .A3(new_n279), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n301), .B(new_n278), .C1(new_n303), .C2(new_n288), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n277), .B(G169), .C1(new_n302), .C2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n301), .B1(new_n303), .B2(new_n288), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT13), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(G179), .A3(new_n304), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n304), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n277), .B1(new_n311), .B2(G169), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n276), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(G190), .A3(new_n304), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT77), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n308), .A2(KEYINPUT77), .A3(G190), .A4(new_n304), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n308), .B2(new_n304), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n276), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT3), .B(G33), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(G232), .A3(new_n296), .ZN(new_n324));
  INV_X1    g0124(.A(G107), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(G1698), .ZN(new_n326));
  INV_X1    g0126(.A(G238), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n324), .B1(new_n325), .B2(new_n323), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n300), .ZN(new_n329));
  INV_X1    g0129(.A(new_n285), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n300), .A2(new_n282), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n221), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n329), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G190), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n266), .A2(G77), .A3(new_n268), .ZN(new_n339));
  XOR2_X1   g0139(.A(new_n339), .B(KEYINPUT73), .Z(new_n340));
  XOR2_X1   g0140(.A(KEYINPUT8), .B(G58), .Z(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT15), .B(G87), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n257), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n264), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n344), .A2(new_n254), .B1(new_n203), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n334), .A2(G200), .A3(new_n336), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n338), .A2(new_n340), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n337), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G169), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n334), .A2(new_n351), .A3(new_n336), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n340), .A2(new_n346), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT74), .B1(new_n348), .B2(new_n354), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n313), .B(new_n322), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT10), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n341), .A2(new_n256), .B1(G150), .B2(new_n259), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n202), .B2(new_n211), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n254), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n266), .A2(G50), .A3(new_n268), .ZN(new_n362));
  INV_X1    g0162(.A(G50), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n345), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT75), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n365), .A2(new_n366), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT9), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n365), .A2(new_n366), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n323), .A2(G222), .A3(new_n296), .ZN(new_n375));
  INV_X1    g0175(.A(G223), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n375), .B1(new_n203), .B2(new_n323), .C1(new_n326), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n300), .ZN(new_n378));
  XOR2_X1   g0178(.A(KEYINPUT69), .B(G226), .Z(new_n379));
  AOI21_X1  g0179(.A(new_n330), .B1(new_n331), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G200), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n381), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n358), .B1(new_n374), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT10), .B(new_n384), .C1(new_n370), .C2(new_n373), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n268), .A2(new_n341), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n389), .A2(new_n265), .B1(new_n264), .B2(new_n341), .ZN(new_n390));
  INV_X1    g0190(.A(new_n254), .ZN(new_n391));
  INV_X1    g0191(.A(G58), .ZN(new_n392));
  INV_X1    g0192(.A(G68), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n394), .B2(new_n206), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n259), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n323), .B2(G20), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n293), .A2(G33), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n401));
  OAI211_X1 g0201(.A(KEYINPUT7), .B(new_n211), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n397), .B1(new_n403), .B2(G68), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n391), .B1(new_n404), .B2(KEYINPUT16), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n393), .B1(new_n399), .B2(new_n402), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n397), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n390), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n292), .A2(new_n294), .A3(G223), .A4(new_n296), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n292), .A2(new_n294), .A3(G226), .A4(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n300), .ZN(new_n414));
  INV_X1    g0214(.A(G274), .ZN(new_n415));
  INV_X1    g0215(.A(new_n210), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(new_n283), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n331), .A2(G232), .B1(new_n417), .B2(new_n282), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G169), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n414), .A2(new_n418), .A3(G179), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT18), .B1(new_n409), .B2(new_n423), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n414), .A2(new_n418), .A3(G190), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n319), .B1(new_n414), .B2(new_n418), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n292), .A2(new_n294), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n428), .B2(new_n211), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n398), .B(G20), .C1(new_n292), .C2(new_n294), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n397), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(KEYINPUT16), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(new_n408), .A3(new_n254), .ZN(new_n434));
  INV_X1    g0234(.A(new_n390), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n427), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n427), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n435), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(new_n422), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n424), .A2(new_n438), .A3(new_n439), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n381), .A2(new_n351), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n378), .A2(new_n349), .A3(new_n380), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n365), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n357), .A2(new_n388), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n292), .A2(new_n294), .A3(G257), .A4(new_n296), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n292), .A2(new_n294), .A3(G264), .A4(G1698), .ZN(new_n452));
  INV_X1    g0252(.A(G303), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n451), .B(new_n452), .C1(new_n453), .C2(new_n323), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n300), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT5), .B(G41), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n214), .A2(G45), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n456), .A2(new_n458), .B1(new_n416), .B2(new_n283), .ZN(new_n459));
  OR2_X1    g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  NAND2_X1  g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n459), .A2(G270), .B1(new_n417), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(KEYINPUT21), .A3(G169), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n349), .B2(new_n464), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT85), .ZN(new_n467));
  AOI21_X1  g0267(.A(G20), .B1(new_n255), .B2(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT84), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT20), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n468), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT83), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G20), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n254), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n254), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n470), .A2(new_n471), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI221_X1 g0280(.A(new_n472), .B1(new_n470), .B2(new_n471), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n264), .A2(new_n474), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n265), .B1(new_n214), .B2(G33), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(new_n474), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n466), .A2(new_n467), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n467), .B1(new_n466), .B2(new_n485), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n351), .B1(new_n455), .B2(new_n463), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT86), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT21), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n485), .A2(KEYINPUT86), .A3(new_n489), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n464), .A2(G200), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n383), .B2(new_n464), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n485), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n488), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT80), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n259), .A2(G77), .ZN(new_n502));
  XNOR2_X1  g0302(.A(G97), .B(G107), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  INV_X1    g0304(.A(G97), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n503), .A2(new_n504), .B1(new_n325), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n502), .B1(new_n507), .B2(new_n211), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n325), .B1(new_n399), .B2(new_n402), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n254), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n483), .A2(G97), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n264), .A2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n292), .A2(new_n294), .A3(G244), .A4(new_n296), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n323), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n323), .A2(G250), .A3(G1698), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n469), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n300), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n462), .A2(new_n417), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n459), .A2(G257), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n520), .A2(new_n300), .B1(G257), .B2(new_n459), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G190), .A3(new_n522), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n514), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n524), .A2(new_n351), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n349), .A3(new_n522), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n501), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n345), .A2(new_n325), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT25), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(G107), .B2(new_n483), .ZN(new_n536));
  NOR2_X1   g0336(.A1(KEYINPUT87), .A2(G20), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n292), .A2(new_n294), .A3(G87), .A4(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT22), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT88), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n211), .B2(G107), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT23), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n541), .B(new_n544), .C1(new_n211), .C2(G107), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G87), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n548), .A2(KEYINPUT87), .A3(G20), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n549), .A2(KEYINPUT22), .A3(new_n292), .A4(new_n294), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT24), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n539), .A2(new_n538), .B1(new_n543), .B2(new_n545), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT89), .B1(new_n558), .B2(new_n254), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT89), .ZN(new_n560));
  AOI211_X1 g0360(.A(new_n560), .B(new_n391), .C1(new_n553), .C2(new_n557), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n536), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT90), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n459), .A2(G264), .B1(new_n417), .B2(new_n462), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n292), .A2(new_n294), .A3(G257), .A4(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n292), .A2(new_n294), .A3(G250), .A4(new_n296), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G294), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n300), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n563), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n564), .A2(new_n569), .A3(new_n563), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(G169), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n564), .A2(new_n569), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(new_n349), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n562), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n547), .A2(new_n552), .A3(KEYINPUT24), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n556), .B1(new_n554), .B2(new_n555), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n254), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n560), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n558), .A2(KEYINPUT89), .A3(new_n254), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n564), .A2(new_n563), .A3(new_n569), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n383), .B1(new_n585), .B2(new_n570), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n574), .A2(new_n319), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n536), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n528), .A2(new_n532), .A3(new_n501), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n257), .B2(new_n505), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n323), .A2(new_n211), .A3(G68), .ZN(new_n593));
  NOR3_X1   g0393(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n594), .B(KEYINPUT81), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n211), .B1(new_n298), .B2(new_n591), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n592), .B(new_n593), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n254), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n343), .A2(new_n345), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n483), .A2(G87), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n417), .A2(new_n458), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n284), .A2(G250), .A3(new_n457), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n292), .A2(new_n294), .A3(G244), .A4(G1698), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n292), .A2(new_n294), .A3(G238), .A4(new_n296), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n255), .C2(new_n474), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n608), .B2(new_n300), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n319), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n300), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n603), .A2(new_n604), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT82), .B1(new_n614), .B2(new_n383), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n609), .A2(new_n616), .A3(G190), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n609), .A2(new_n349), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n351), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n343), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n483), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n599), .A2(new_n623), .A3(new_n600), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n611), .A2(new_n618), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n578), .A2(new_n589), .A3(new_n590), .A4(new_n625), .ZN(new_n626));
  NOR4_X1   g0426(.A1(new_n450), .A2(new_n500), .A3(new_n533), .A4(new_n626), .ZN(G372));
  AOI211_X1 g0427(.A(new_n276), .B(new_n320), .C1(new_n316), .C2(new_n317), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n313), .B1(new_n628), .B2(new_n354), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n438), .A2(new_n439), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT92), .ZN(new_n632));
  AOI221_X4 g0432(.A(KEYINPUT18), .B1(new_n420), .B2(new_n421), .C1(new_n434), .C2(new_n435), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n441), .B1(new_n440), .B2(new_n422), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n424), .A2(KEYINPUT92), .A3(new_n442), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n388), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n447), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n624), .A2(new_n620), .A3(new_n619), .ZN(new_n640));
  INV_X1    g0440(.A(new_n532), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT26), .B1(new_n625), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n614), .A2(KEYINPUT82), .A3(new_n383), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n616), .B1(new_n609), .B2(G190), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n614), .A2(G200), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(new_n600), .A3(new_n599), .A4(new_n601), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n640), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n648), .A2(new_n649), .A3(new_n532), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n640), .B1(new_n642), .B2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n532), .A2(new_n589), .A3(new_n528), .A4(new_n625), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n466), .A2(new_n485), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n495), .A2(new_n653), .A3(new_n578), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n651), .B1(new_n655), .B2(KEYINPUT91), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT91), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n652), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n639), .B1(new_n450), .B2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n214), .A2(new_n211), .A3(G13), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(G213), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n494), .A2(new_n493), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT86), .B1(new_n485), .B2(new_n489), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n485), .B(new_n667), .C1(new_n670), .C2(new_n466), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n672));
  INV_X1    g0472(.A(new_n667), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n671), .B1(new_n500), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n562), .A2(new_n667), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n578), .A2(new_n678), .A3(new_n589), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT93), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n578), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n667), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n677), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n673), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n488), .A2(new_n495), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n681), .A2(new_n689), .A3(new_n673), .A4(new_n682), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(G399));
  INV_X1    g0491(.A(KEYINPUT81), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n594), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G116), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n227), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n208), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  INV_X1    g0499(.A(new_n651), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n652), .B1(new_n689), .B2(new_n684), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n667), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n667), .B1(new_n656), .B2(new_n658), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(KEYINPUT29), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n464), .A2(new_n614), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n575), .A3(KEYINPUT30), .A4(new_n526), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT94), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n521), .A2(new_n523), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n455), .A2(new_n612), .A3(new_n463), .A4(new_n613), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT30), .A4(new_n575), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n455), .A2(new_n463), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n526), .A3(new_n609), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n576), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(G179), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n524), .A3(new_n574), .A4(new_n614), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n708), .A2(new_n713), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n667), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(KEYINPUT21), .A2(new_n489), .B1(new_n715), .B2(G179), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT85), .B1(new_n672), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n466), .A2(new_n467), .A3(new_n485), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n670), .A2(new_n731), .A3(new_n498), .ZN(new_n732));
  AND4_X1   g0532(.A1(new_n590), .A2(new_n578), .A3(new_n589), .A4(new_n625), .ZN(new_n733));
  INV_X1    g0533(.A(new_n533), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n732), .A2(new_n733), .A3(new_n734), .A4(new_n673), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n723), .A2(KEYINPUT95), .A3(new_n724), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n727), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n705), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n699), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n226), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n214), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n695), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n677), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n675), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n228), .A2(new_n323), .ZN(new_n748));
  INV_X1    g0548(.A(G355), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n749), .B1(G116), .B2(new_n228), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n245), .A2(new_n281), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n227), .A2(new_n323), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n281), .B2(new_n209), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n210), .B1(G20), .B2(new_n351), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT96), .Z(new_n761));
  OAI21_X1  g0561(.A(new_n745), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n211), .A2(new_n383), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n349), .A2(G200), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G322), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n211), .A2(G190), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n768), .A2(new_n764), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n766), .A2(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n763), .A2(new_n349), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n323), .B(new_n772), .C1(G303), .C2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n383), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n211), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n211), .A2(new_n349), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n779), .A2(new_n383), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n768), .A2(new_n349), .A3(new_n319), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT97), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G329), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n768), .A2(new_n349), .A3(G200), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G283), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n775), .A2(new_n786), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n766), .A2(new_n392), .B1(new_n770), .B2(new_n203), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n777), .A2(new_n505), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n363), .B2(new_n780), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n798), .B(new_n801), .C1(G68), .C2(new_n784), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n773), .A2(new_n548), .ZN(new_n803));
  OR3_X1    g0603(.A1(new_n803), .A2(KEYINPUT98), .A3(new_n428), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n795), .A2(G107), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT98), .B1(new_n803), .B2(new_n428), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n802), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n792), .A2(G159), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n797), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n762), .B1(new_n810), .B2(new_n759), .ZN(new_n811));
  INV_X1    g0611(.A(new_n758), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n675), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n747), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND3_X1  g0615(.A1(new_n348), .A2(new_n354), .A3(new_n673), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n659), .A2(new_n817), .ZN(new_n818));
  AND4_X1   g0618(.A1(new_n352), .A2(new_n350), .A3(new_n353), .A4(new_n673), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n353), .A2(new_n667), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n348), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n821), .B2(new_n354), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n818), .B1(new_n704), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n745), .B1(new_n823), .B2(new_n738), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n738), .B2(new_n823), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n795), .A2(G87), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n771), .B2(new_n791), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT100), .Z(new_n828));
  AOI22_X1  g0628(.A1(G294), .A2(new_n765), .B1(new_n769), .B2(G116), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n428), .C1(new_n325), .C2(new_n773), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n800), .B1(new_n783), .B2(new_n831), .C1(new_n453), .C2(new_n780), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n828), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n323), .B1(new_n773), .B2(new_n363), .C1(new_n392), .C2(new_n777), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n792), .B2(G132), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n795), .A2(G68), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT101), .B(G143), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n765), .A2(new_n837), .B1(new_n769), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n839), .B2(new_n780), .C1(new_n840), .C2(new_n783), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n835), .B(new_n836), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n759), .B1(new_n833), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n745), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n759), .A2(new_n756), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n203), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n845), .B(new_n848), .C1(new_n822), .C2(new_n757), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n825), .A2(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n742), .A2(new_n214), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT39), .ZN(new_n852));
  INV_X1    g0652(.A(new_n665), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT104), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n433), .A2(new_n254), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n431), .A2(new_n432), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT103), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT16), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n404), .A2(KEYINPUT103), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n854), .B1(new_n860), .B2(new_n390), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n857), .B1(new_n407), .B2(new_n397), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(new_n406), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n405), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(KEYINPUT104), .A3(new_n435), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n443), .A2(new_n853), .A3(new_n861), .A4(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n423), .A2(new_n665), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n869), .B2(new_n436), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n440), .A2(new_n853), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n871), .B(new_n436), .C1(new_n409), .C2(new_n423), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  OAI211_X1 g0673(.A(KEYINPUT38), .B(new_n866), .C1(new_n870), .C2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n635), .A2(new_n630), .A3(new_n636), .ZN(new_n876));
  INV_X1    g0676(.A(new_n871), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n872), .B(KEYINPUT37), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n852), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n866), .B1(new_n870), .B2(new_n873), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n874), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n313), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n673), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n819), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n818), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n874), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n276), .A2(new_n667), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n311), .A2(G169), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT14), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n309), .A3(new_n306), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n895), .B1(new_n628), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n313), .A2(new_n322), .A3(new_n894), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(KEYINPUT102), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT102), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n902), .B(new_n895), .C1(new_n628), .C2(new_n898), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n892), .A2(new_n893), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n635), .A2(new_n636), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n665), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n890), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n703), .B(new_n449), .C1(new_n704), .C2(KEYINPUT29), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n639), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT107), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT31), .B1(new_n720), .B2(new_n667), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT105), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n724), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n720), .A2(KEYINPUT105), .A3(KEYINPUT31), .A4(new_n667), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR4_X1   g0718(.A1(new_n500), .A2(new_n626), .A3(new_n533), .A4(new_n667), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n901), .A2(new_n903), .A3(new_n822), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n875), .A2(new_n880), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n901), .A2(new_n822), .A3(new_n903), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n735), .A2(new_n916), .A3(new_n917), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT107), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT106), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT40), .B1(new_n884), .B2(new_n874), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT106), .B1(new_n924), .B2(new_n925), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n927), .A2(KEYINPUT40), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n450), .B2(new_n920), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n875), .A2(new_n880), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n924), .A2(new_n925), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n937), .B2(new_n913), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n935), .B1(new_n938), .B2(new_n926), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n928), .A2(new_n929), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(new_n931), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n449), .B(new_n925), .C1(new_n939), .C2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(G330), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n851), .B1(new_n912), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n912), .B2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(new_n507), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT35), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT35), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(G116), .A4(new_n212), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n208), .A2(new_n203), .A3(new_n394), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n393), .A2(G50), .ZN(new_n952));
  OAI211_X1 g0752(.A(G1), .B(new_n226), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n945), .A2(new_n950), .A3(new_n953), .ZN(G367));
  NAND2_X1  g0754(.A1(new_n602), .A2(new_n667), .ZN(new_n955));
  MUX2_X1   g0755(.A(new_n640), .B(new_n648), .S(new_n955), .Z(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT108), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n758), .ZN(new_n959));
  INV_X1    g0759(.A(new_n761), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n228), .B2(new_n343), .C1(new_n236), .C2(new_n753), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT111), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n846), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n961), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n766), .A2(new_n840), .B1(new_n203), .B2(new_n794), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G58), .B2(new_n774), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n792), .A2(G137), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n323), .B1(new_n770), .B2(new_n363), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G159), .B2(new_n784), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n777), .A2(new_n393), .ZN(new_n970));
  INV_X1    g0770(.A(new_n780), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(new_n971), .B2(new_n837), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n966), .A2(new_n967), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n773), .A2(new_n474), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT46), .ZN(new_n975));
  INV_X1    g0775(.A(new_n777), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(G107), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n792), .A2(G317), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n428), .B1(new_n770), .B2(new_n831), .ZN(new_n979));
  INV_X1    g0779(.A(new_n794), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(G97), .B2(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n974), .A2(KEYINPUT46), .B1(new_n784), .B2(G294), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n977), .A2(new_n978), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n766), .A2(new_n453), .B1(new_n771), .B2(new_n780), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT112), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n973), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n964), .B1(new_n987), .B2(new_n759), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n959), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n528), .A2(new_n532), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n514), .A2(new_n673), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n990), .A2(new_n991), .B1(new_n532), .B2(new_n673), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT110), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n690), .A2(new_n688), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n690), .A2(new_n688), .ZN(new_n999));
  INV_X1    g0799(.A(new_n994), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT44), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1002), .B(new_n994), .C1(new_n690), .C2(new_n688), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n997), .A2(new_n998), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n687), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n994), .B1(new_n690), .B2(new_n688), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT44), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n995), .B(new_n996), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n687), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n689), .A2(new_n673), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n683), .A2(new_n685), .A3(new_n1011), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n1012), .A2(new_n676), .A3(new_n690), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n676), .B1(new_n1012), .B2(new_n690), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n739), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1006), .A2(new_n1010), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n740), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n695), .B(KEYINPUT41), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n744), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n690), .A2(new_n1000), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT42), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n532), .B1(new_n1000), .B2(new_n578), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n673), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n1024), .A3(new_n958), .A4(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1027));
  MUX2_X1   g0827(.A(new_n1025), .B(KEYINPUT43), .S(new_n957), .Z(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n687), .A2(new_n1000), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1030), .B(new_n1026), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n989), .B1(new_n1020), .B2(new_n1034), .ZN(G387));
  INV_X1    g0835(.A(new_n1016), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n739), .A2(new_n1015), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n695), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n686), .A2(new_n812), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n759), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n777), .A2(new_n831), .B1(new_n773), .B2(new_n778), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G317), .A2(new_n765), .B1(new_n769), .B2(G303), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n771), .B2(new_n783), .C1(new_n767), .C2(new_n780), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n428), .B1(new_n474), .B2(new_n794), .C1(new_n791), .C2(new_n781), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n766), .A2(new_n363), .B1(new_n203), .B2(new_n773), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n428), .B(new_n1052), .C1(G68), .C2(new_n769), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n976), .A2(new_n622), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n341), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n783), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G159), .B2(new_n971), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n792), .A2(G150), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n795), .A2(G97), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1053), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1040), .B1(new_n1051), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n341), .A2(new_n363), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT50), .Z(new_n1063));
  AOI21_X1  g0863(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT113), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1064), .C1(new_n1065), .C2(new_n694), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n694), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1067), .A2(KEYINPUT113), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n752), .B1(new_n281), .B2(new_n241), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(G107), .B2(new_n228), .C1(new_n694), .C2(new_n748), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n846), .B(new_n1061), .C1(new_n960), .C2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT114), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1038), .B1(new_n743), .B2(new_n1015), .C1(new_n1039), .C2(new_n1072), .ZN(G393));
  NAND2_X1  g0873(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n1036), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n695), .A3(new_n1017), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n687), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT115), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT115), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1006), .A2(new_n1010), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n744), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n777), .A2(new_n203), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n323), .B1(new_n393), .B2(new_n773), .C1(new_n770), .C2(new_n1055), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(G50), .C2(new_n784), .ZN(new_n1085));
  INV_X1    g0885(.A(G159), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n766), .A2(new_n1086), .B1(new_n840), .B2(new_n780), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n792), .A2(new_n837), .ZN(new_n1089));
  AND4_X1   g0889(.A1(new_n826), .A2(new_n1085), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n428), .B1(new_n770), .B2(new_n778), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G283), .B2(new_n774), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n805), .C1(new_n767), .C2(new_n791), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n777), .A2(new_n474), .B1(new_n783), .B2(new_n453), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT116), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n971), .A2(G317), .B1(new_n765), .B2(G311), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n759), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n761), .B1(G97), .B2(new_n227), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n248), .A2(new_n752), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n846), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1000), .B2(new_n758), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1076), .A2(new_n1082), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT117), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n743), .B1(new_n1074), .B2(KEYINPUT115), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1104), .B1(new_n1109), .B2(new_n1081), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(KEYINPUT117), .A3(new_n1076), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(G390));
  NAND3_X1  g0912(.A1(new_n737), .A2(G330), .A3(new_n822), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT118), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n924), .A2(new_n925), .A3(new_n1115), .A4(G330), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n905), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n821), .A2(new_n354), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n819), .B1(new_n702), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n888), .B(new_n923), .C1(new_n1119), .C2(new_n904), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n889), .B1(new_n892), .B2(new_n905), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1117), .B(new_n1120), .C1(new_n1121), .C2(new_n886), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n925), .A2(G330), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1123), .A2(new_n1115), .A3(new_n921), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n816), .B1(new_n656), .B2(new_n658), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n905), .B1(new_n1125), .B2(new_n819), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1126), .A2(new_n888), .B1(new_n881), .B2(new_n885), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1120), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1122), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n822), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n904), .B1(new_n1123), .B2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1132), .B(new_n1119), .C1(new_n904), .C2(new_n1113), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1123), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n904), .A2(new_n1113), .B1(new_n1134), .B2(new_n924), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n892), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n449), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n910), .A3(new_n639), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1130), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n696), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1122), .A2(new_n1129), .A3(new_n744), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n846), .B1(new_n1055), .B2(new_n847), .ZN(new_n1146));
  INV_X1    g0946(.A(G132), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n766), .A2(new_n1147), .B1(new_n363), .B2(new_n794), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n428), .B(new_n1148), .C1(new_n769), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n773), .A2(new_n840), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT53), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1152), .A2(new_n1153), .B1(new_n1086), .B2(new_n777), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n792), .A2(G125), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G128), .A2(new_n971), .B1(new_n784), .B2(G137), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1151), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n766), .A2(new_n474), .B1(new_n770), .B2(new_n505), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1159), .A2(new_n323), .A3(new_n803), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n780), .A2(new_n831), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1161), .B(new_n1083), .C1(G107), .C2(new_n784), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n792), .A2(G294), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1162), .A3(new_n1163), .A4(new_n836), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1146), .B1(new_n1040), .B2(new_n1165), .C1(new_n886), .C2(new_n757), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1144), .A2(new_n1145), .A3(new_n1166), .ZN(G378));
  OAI21_X1  g0967(.A(new_n1140), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT120), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n446), .B1(new_n386), .B2(new_n387), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n371), .A2(new_n367), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n853), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n446), .B(new_n1172), .C1(new_n386), .C2(new_n387), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1169), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1176), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(KEYINPUT120), .A3(new_n1177), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(G330), .B(new_n1185), .C1(new_n939), .C2(new_n941), .ZN(new_n1186));
  INV_X1    g0986(.A(G330), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n927), .A2(KEYINPUT40), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n930), .A2(new_n932), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1186), .B(new_n909), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1191), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n933), .B2(new_n1187), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n909), .B1(new_n1195), .B2(new_n1186), .ZN(new_n1196));
  OAI211_X1 g0996(.A(KEYINPUT57), .B(new_n1168), .C1(new_n1193), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n695), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n909), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1192), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1168), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1198), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1185), .A2(new_n756), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n847), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n745), .B1(G50), .B2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT119), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n777), .A2(new_n840), .B1(new_n783), .B2(new_n1147), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n774), .A2(new_n1150), .B1(new_n765), .B2(G128), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n769), .A2(G137), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1209), .B(new_n1212), .C1(G125), .C2(new_n971), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n255), .A2(new_n280), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n794), .A2(new_n1086), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(new_n792), .C2(G124), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1215), .A2(new_n1216), .A3(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n980), .A2(G58), .B1(new_n765), .B2(G107), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n343), .B2(new_n770), .C1(new_n791), .C2(new_n831), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n280), .B(new_n428), .C1(new_n773), .C2(new_n203), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n783), .A2(new_n505), .B1(new_n780), .B2(new_n474), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1222), .A2(new_n970), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n363), .B(new_n1217), .C1(new_n323), .C2(G41), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1220), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1208), .B1(new_n1229), .B2(new_n759), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1202), .A2(new_n744), .B1(new_n1205), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1204), .A2(new_n1231), .ZN(G375));
  OAI211_X1 g1032(.A(new_n1133), .B(new_n1139), .C1(new_n1136), .C2(new_n1135), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1141), .A2(new_n1019), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n323), .B1(new_n795), .B2(G77), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT121), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1054), .B1(new_n783), .B2(new_n474), .C1(new_n778), .C2(new_n780), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n791), .A2(new_n453), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n774), .A2(G97), .B1(new_n769), .B2(G107), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n831), .B2(new_n766), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n976), .A2(G50), .B1(G150), .B2(new_n769), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT123), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n323), .B1(new_n794), .B2(new_n392), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n766), .A2(new_n839), .B1(new_n1086), .B2(new_n773), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n784), .C2(new_n1150), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n971), .A2(G132), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT122), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n792), .A2(G128), .ZN(new_n1249));
  AND4_X1   g1049(.A1(new_n1243), .A2(new_n1246), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n759), .B1(new_n1241), .B2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n745), .C1(G68), .C2(new_n1206), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n904), .B2(new_n756), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1137), .B2(new_n744), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1234), .A2(new_n1254), .ZN(G381));
  OR3_X1    g1055(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(G390), .A2(new_n1256), .A3(G387), .A4(G381), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT124), .Z(new_n1258));
  INV_X1    g1058(.A(G375), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1144), .A2(new_n1145), .A3(new_n1166), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1258), .A2(new_n1261), .ZN(G407));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n666), .A3(new_n1260), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1263), .B(G213), .C1(new_n1258), .C2(new_n1261), .ZN(G409));
  XNOR2_X1  g1064(.A(G393), .B(new_n814), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1108), .A2(G387), .A3(new_n1111), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G387), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G387), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT117), .B1(new_n1110), .B2(new_n1076), .ZN(new_n1271));
  AND4_X1   g1071(.A1(KEYINPUT117), .A2(new_n1076), .A3(new_n1082), .A4(new_n1105), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1108), .A2(G387), .A3(new_n1111), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1265), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G378), .B(new_n1231), .C1(new_n1198), .C2(new_n1203), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1019), .B(new_n1168), .C1(new_n1193), .C2(new_n1196), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n744), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1205), .A2(new_n1230), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1260), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  INV_X1    g1084(.A(G213), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1285), .A2(G343), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1233), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(KEYINPUT60), .B2(new_n1141), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1290), .A2(KEYINPUT60), .A3(new_n1139), .A4(new_n1133), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n695), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1254), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(G384), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G384), .B(new_n1254), .C1(new_n1289), .C2(new_n1292), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1283), .A2(new_n1284), .A3(new_n1287), .A4(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1286), .B1(new_n1277), .B2(new_n1282), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1286), .A2(KEYINPUT125), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1295), .A2(new_n1296), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1286), .A2(G2897), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1303), .B(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1299), .B(new_n1300), .C1(new_n1301), .C2(new_n1306), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n1286), .B(new_n1297), .C1(new_n1277), .C2(new_n1282), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1308), .A2(new_n1284), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1276), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1269), .A2(new_n1300), .A3(new_n1275), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(KEYINPUT63), .B2(new_n1308), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1303), .B(new_n1304), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1313), .B2(new_n1297), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT126), .B1(new_n1306), .B2(new_n1301), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1312), .A2(new_n1316), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1310), .A2(new_n1320), .ZN(G405));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1277), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1297), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1277), .A2(new_n1298), .A3(new_n1322), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(new_n1260), .A3(G375), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1276), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G375), .A2(new_n1260), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1324), .A2(new_n1329), .A3(new_n1325), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1327), .A2(new_n1328), .A3(new_n1330), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1324), .A2(new_n1329), .A3(new_n1325), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1329), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1276), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1331), .A2(new_n1334), .ZN(G402));
endmodule


