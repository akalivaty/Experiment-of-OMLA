

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(n817), .A2(n816), .ZN(n827) );
  OR2_X1 U553 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X2 U554 ( .A1(n671), .A2(n670), .ZN(G160) );
  NAND2_X1 U555 ( .A1(n741), .A2(n740), .ZN(n810) );
  NOR2_X1 U556 ( .A1(n686), .A2(n687), .ZN(n679) );
  BUF_X1 U557 ( .A(n890), .Z(n516) );
  XOR2_X1 U558 ( .A(KEYINPUT17), .B(n517), .Z(n890) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n703) );
  NOR2_X1 U560 ( .A1(G1384), .A2(G164), .ZN(n672) );
  XNOR2_X1 U561 ( .A(KEYINPUT66), .B(G2104), .ZN(n520) );
  AND2_X1 U562 ( .A1(n971), .A2(n759), .ZN(n817) );
  NOR2_X1 U563 ( .A1(G651), .A2(n614), .ZN(n634) );
  AND2_X1 U564 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  NAND2_X1 U566 ( .A1(G138), .A2(n890), .ZN(n519) );
  INV_X1 U567 ( .A(G2105), .ZN(n521) );
  NOR2_X2 U568 ( .A1(n521), .A2(n520), .ZN(n897) );
  NAND2_X1 U569 ( .A1(G126), .A2(n897), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n519), .A2(n518), .ZN(n525) );
  AND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n892) );
  NAND2_X1 U572 ( .A1(G102), .A2(n892), .ZN(n523) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n896) );
  NAND2_X1 U574 ( .A1(G114), .A2(n896), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U576 ( .A1(n525), .A2(n524), .ZN(G164) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n626) );
  NAND2_X1 U578 ( .A1(n626), .A2(G85), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n614) );
  XNOR2_X1 U580 ( .A(KEYINPUT67), .B(G651), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n614), .A2(n528), .ZN(n630) );
  NAND2_X1 U582 ( .A1(G72), .A2(n630), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n634), .A2(G47), .ZN(n531) );
  NOR2_X1 U585 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n529), .Z(n627) );
  NAND2_X1 U587 ( .A1(G60), .A2(n627), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n531), .A2(n530), .ZN(n532) );
  OR2_X1 U589 ( .A1(n533), .A2(n532), .ZN(G290) );
  NAND2_X1 U590 ( .A1(G77), .A2(n630), .ZN(n534) );
  XOR2_X1 U591 ( .A(KEYINPUT69), .B(n534), .Z(n536) );
  NAND2_X1 U592 ( .A1(n626), .A2(G90), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U594 ( .A(n537), .B(KEYINPUT9), .ZN(n539) );
  NAND2_X1 U595 ( .A1(G52), .A2(n634), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n627), .A2(G64), .ZN(n540) );
  XOR2_X1 U598 ( .A(KEYINPUT68), .B(n540), .Z(n541) );
  NOR2_X1 U599 ( .A1(n542), .A2(n541), .ZN(G171) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U601 ( .A1(n897), .A2(G123), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n543), .B(KEYINPUT18), .ZN(n545) );
  NAND2_X1 U603 ( .A1(G135), .A2(n516), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U605 ( .A(KEYINPUT78), .B(n546), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G99), .A2(n892), .ZN(n547) );
  XNOR2_X1 U607 ( .A(KEYINPUT79), .B(n547), .ZN(n548) );
  NOR2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n896), .A2(G111), .ZN(n550) );
  NAND2_X1 U610 ( .A1(n551), .A2(n550), .ZN(n927) );
  XNOR2_X1 U611 ( .A(G2096), .B(n927), .ZN(n552) );
  OR2_X1 U612 ( .A1(G2100), .A2(n552), .ZN(G156) );
  INV_X1 U613 ( .A(G120), .ZN(G236) );
  INV_X1 U614 ( .A(G132), .ZN(G219) );
  INV_X1 U615 ( .A(G82), .ZN(G220) );
  NAND2_X1 U616 ( .A1(n634), .A2(G51), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G63), .A2(n627), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT6), .B(n555), .Z(n563) );
  NAND2_X1 U620 ( .A1(G76), .A2(n630), .ZN(n556) );
  XNOR2_X1 U621 ( .A(KEYINPUT75), .B(n556), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n626), .A2(G89), .ZN(n557) );
  XOR2_X1 U623 ( .A(n557), .B(KEYINPUT4), .Z(n558) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT5), .B(n560), .Z(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT76), .B(n561), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U628 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U632 ( .A(G223), .B(KEYINPUT71), .ZN(n829) );
  NAND2_X1 U633 ( .A1(n829), .A2(G567), .ZN(n566) );
  XOR2_X1 U634 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  NAND2_X1 U635 ( .A1(G81), .A2(n626), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n567), .B(KEYINPUT12), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n568), .B(KEYINPUT72), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G68), .A2(n630), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U640 ( .A(KEYINPUT13), .B(n571), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n627), .A2(G56), .ZN(n572) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n572), .Z(n575) );
  NAND2_X1 U643 ( .A1(G43), .A2(n634), .ZN(n573) );
  XNOR2_X1 U644 ( .A(KEYINPUT73), .B(n573), .ZN(n574) );
  NOR2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n984) );
  INV_X1 U647 ( .A(G860), .ZN(n598) );
  OR2_X1 U648 ( .A1(n984), .A2(n598), .ZN(G153) );
  INV_X1 U649 ( .A(G171), .ZN(G301) );
  NAND2_X1 U650 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n634), .A2(G54), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G79), .A2(n630), .ZN(n579) );
  NAND2_X1 U653 ( .A1(G66), .A2(n627), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n626), .A2(G92), .ZN(n580) );
  XOR2_X1 U656 ( .A(KEYINPUT74), .B(n580), .Z(n581) );
  NOR2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U659 ( .A(KEYINPUT15), .B(n585), .ZN(n983) );
  INV_X1 U660 ( .A(n983), .ZN(n686) );
  INV_X1 U661 ( .A(G868), .ZN(n637) );
  NAND2_X1 U662 ( .A1(n686), .A2(n637), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G78), .A2(n630), .ZN(n589) );
  NAND2_X1 U665 ( .A1(G65), .A2(n627), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n626), .A2(G91), .ZN(n590) );
  XOR2_X1 U668 ( .A(KEYINPUT70), .B(n590), .Z(n591) );
  NOR2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n634), .A2(G53), .ZN(n593) );
  NAND2_X1 U671 ( .A1(n594), .A2(n593), .ZN(G299) );
  XOR2_X1 U672 ( .A(KEYINPUT77), .B(n637), .Z(n595) );
  NOR2_X1 U673 ( .A1(G286), .A2(n595), .ZN(n597) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n599), .A2(n983), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n984), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n983), .A2(G868), .ZN(n601) );
  NOR2_X1 U681 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U682 ( .A1(n603), .A2(n602), .ZN(G282) );
  XNOR2_X1 U683 ( .A(KEYINPUT80), .B(n984), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n983), .A2(G559), .ZN(n648) );
  XNOR2_X1 U685 ( .A(n604), .B(n648), .ZN(n605) );
  NOR2_X1 U686 ( .A1(G860), .A2(n605), .ZN(n613) );
  NAND2_X1 U687 ( .A1(G80), .A2(n630), .ZN(n607) );
  NAND2_X1 U688 ( .A1(G67), .A2(n627), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G93), .A2(n626), .ZN(n608) );
  XNOR2_X1 U691 ( .A(KEYINPUT81), .B(n608), .ZN(n609) );
  NOR2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n634), .A2(G55), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n646) );
  XOR2_X1 U695 ( .A(n613), .B(n646), .Z(G145) );
  NAND2_X1 U696 ( .A1(G87), .A2(n614), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G74), .A2(G651), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U699 ( .A1(n627), .A2(n617), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n634), .A2(G49), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(G288) );
  NAND2_X1 U702 ( .A1(n626), .A2(G88), .ZN(n621) );
  NAND2_X1 U703 ( .A1(G75), .A2(n630), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n634), .A2(G50), .ZN(n623) );
  NAND2_X1 U706 ( .A1(G62), .A2(n627), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U708 ( .A1(n625), .A2(n624), .ZN(G166) );
  INV_X1 U709 ( .A(G166), .ZN(G303) );
  NAND2_X1 U710 ( .A1(n626), .A2(G86), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G61), .A2(n627), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n630), .A2(G73), .ZN(n631) );
  XOR2_X1 U714 ( .A(KEYINPUT2), .B(n631), .Z(n632) );
  NOR2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n634), .A2(G48), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U718 ( .A1(n637), .A2(n646), .ZN(n638) );
  XNOR2_X1 U719 ( .A(n638), .B(KEYINPUT84), .ZN(n651) );
  XNOR2_X1 U720 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n640) );
  XNOR2_X1 U721 ( .A(G288), .B(KEYINPUT19), .ZN(n639) );
  XNOR2_X1 U722 ( .A(n640), .B(n639), .ZN(n641) );
  XOR2_X1 U723 ( .A(G299), .B(n641), .Z(n643) );
  XOR2_X1 U724 ( .A(G290), .B(G303), .Z(n642) );
  XNOR2_X1 U725 ( .A(n643), .B(n642), .ZN(n644) );
  XOR2_X1 U726 ( .A(n644), .B(G305), .Z(n645) );
  XNOR2_X1 U727 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U728 ( .A(n984), .B(n647), .ZN(n912) );
  XOR2_X1 U729 ( .A(n912), .B(n648), .Z(n649) );
  NAND2_X1 U730 ( .A1(G868), .A2(n649), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n652) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n652), .Z(n653) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n653), .ZN(n654) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n654), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n655), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U738 ( .A1(G220), .A2(G219), .ZN(n656) );
  XOR2_X1 U739 ( .A(KEYINPUT22), .B(n656), .Z(n657) );
  NOR2_X1 U740 ( .A1(G218), .A2(n657), .ZN(n658) );
  NAND2_X1 U741 ( .A1(G96), .A2(n658), .ZN(n834) );
  NAND2_X1 U742 ( .A1(n834), .A2(G2106), .ZN(n662) );
  NAND2_X1 U743 ( .A1(G69), .A2(G108), .ZN(n659) );
  NOR2_X1 U744 ( .A1(G236), .A2(n659), .ZN(n660) );
  NAND2_X1 U745 ( .A1(G57), .A2(n660), .ZN(n835) );
  NAND2_X1 U746 ( .A1(n835), .A2(G567), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n847) );
  NAND2_X1 U748 ( .A1(G661), .A2(G483), .ZN(n663) );
  XOR2_X1 U749 ( .A(KEYINPUT85), .B(n663), .Z(n664) );
  NOR2_X1 U750 ( .A1(n847), .A2(n664), .ZN(n833) );
  NAND2_X1 U751 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U752 ( .A1(n516), .A2(G137), .ZN(n667) );
  NAND2_X1 U753 ( .A1(G101), .A2(n892), .ZN(n665) );
  XOR2_X1 U754 ( .A(KEYINPUT23), .B(n665), .Z(n666) );
  NAND2_X1 U755 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U756 ( .A1(G113), .A2(n896), .ZN(n669) );
  NAND2_X1 U757 ( .A1(G125), .A2(n897), .ZN(n668) );
  NAND2_X1 U758 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U759 ( .A(G1981), .B(G305), .Z(n971) );
  NAND2_X1 U760 ( .A1(G160), .A2(G40), .ZN(n777) );
  XOR2_X1 U761 ( .A(KEYINPUT64), .B(n672), .Z(n778) );
  NOR2_X2 U762 ( .A1(n777), .A2(n778), .ZN(n705) );
  NAND2_X1 U763 ( .A1(G1996), .A2(n705), .ZN(n673) );
  XNOR2_X1 U764 ( .A(n673), .B(KEYINPUT26), .ZN(n675) );
  INV_X1 U765 ( .A(n705), .ZN(n680) );
  NAND2_X1 U766 ( .A1(G1341), .A2(n680), .ZN(n674) );
  NAND2_X1 U767 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U768 ( .A(n676), .B(KEYINPUT94), .ZN(n677) );
  NOR2_X1 U769 ( .A1(n677), .A2(n984), .ZN(n678) );
  XNOR2_X1 U770 ( .A(n678), .B(KEYINPUT65), .ZN(n687) );
  XNOR2_X1 U771 ( .A(n679), .B(KEYINPUT95), .ZN(n684) );
  NOR2_X1 U772 ( .A1(n705), .A2(G1348), .ZN(n682) );
  NOR2_X1 U773 ( .A1(G2067), .A2(n680), .ZN(n681) );
  NOR2_X1 U774 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U775 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U776 ( .A(n685), .B(KEYINPUT96), .ZN(n695) );
  NAND2_X1 U777 ( .A1(n687), .A2(n686), .ZN(n693) );
  INV_X1 U778 ( .A(G299), .ZN(n698) );
  NAND2_X1 U779 ( .A1(n680), .A2(G1956), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n705), .A2(G2072), .ZN(n688) );
  XOR2_X1 U781 ( .A(KEYINPUT27), .B(n688), .Z(n689) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U783 ( .A(n691), .B(KEYINPUT93), .ZN(n697) );
  NOR2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n692) );
  XOR2_X1 U785 ( .A(n692), .B(KEYINPUT28), .Z(n696) );
  AND2_X1 U786 ( .A1(n693), .A2(n696), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n702) );
  INV_X1 U788 ( .A(n696), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n699) );
  OR2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n704) );
  XNOR2_X1 U792 ( .A(n704), .B(n703), .ZN(n709) );
  NAND2_X1 U793 ( .A1(G1961), .A2(n680), .ZN(n707) );
  XOR2_X1 U794 ( .A(KEYINPUT25), .B(G2078), .Z(n958) );
  NAND2_X1 U795 ( .A1(n705), .A2(n958), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n710) );
  OR2_X1 U797 ( .A1(G301), .A2(n710), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n733) );
  NAND2_X1 U799 ( .A1(G301), .A2(n710), .ZN(n711) );
  XNOR2_X1 U800 ( .A(n711), .B(KEYINPUT97), .ZN(n716) );
  NAND2_X1 U801 ( .A1(G8), .A2(n680), .ZN(n812) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n812), .ZN(n736) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n680), .ZN(n734) );
  NOR2_X1 U804 ( .A1(n736), .A2(n734), .ZN(n712) );
  NAND2_X1 U805 ( .A1(G8), .A2(n712), .ZN(n713) );
  XNOR2_X1 U806 ( .A(KEYINPUT30), .B(n713), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n714), .A2(G168), .ZN(n715) );
  NOR2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U809 ( .A(KEYINPUT31), .B(n717), .Z(n732) );
  INV_X1 U810 ( .A(G8), .ZN(n724) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n812), .ZN(n718) );
  XNOR2_X1 U812 ( .A(n718), .B(KEYINPUT98), .ZN(n720) );
  NOR2_X1 U813 ( .A1(n680), .A2(G2090), .ZN(n719) );
  NOR2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U815 ( .A1(n721), .A2(G303), .ZN(n722) );
  XOR2_X1 U816 ( .A(KEYINPUT99), .B(n722), .Z(n723) );
  OR2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n726) );
  AND2_X1 U818 ( .A1(n732), .A2(n726), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n733), .A2(n725), .ZN(n730) );
  INV_X1 U820 ( .A(n726), .ZN(n728) );
  AND2_X1 U821 ( .A1(G286), .A2(G8), .ZN(n727) );
  OR2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U824 ( .A(n731), .B(KEYINPUT32), .ZN(n741) );
  AND2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n739) );
  NAND2_X1 U826 ( .A1(G8), .A2(n734), .ZN(n735) );
  XOR2_X1 U827 ( .A(KEYINPUT92), .B(n735), .Z(n737) );
  OR2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n742) );
  NOR2_X1 U831 ( .A1(n753), .A2(n742), .ZN(n980) );
  INV_X1 U832 ( .A(KEYINPUT33), .ZN(n743) );
  AND2_X1 U833 ( .A1(n980), .A2(n743), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n810), .A2(n744), .ZN(n750) );
  NAND2_X1 U835 ( .A1(G288), .A2(G1976), .ZN(n745) );
  XOR2_X1 U836 ( .A(KEYINPUT100), .B(n745), .Z(n975) );
  INV_X1 U837 ( .A(n975), .ZN(n747) );
  NOR2_X1 U838 ( .A1(KEYINPUT101), .A2(n812), .ZN(n746) );
  AND2_X1 U839 ( .A1(n747), .A2(n746), .ZN(n748) );
  OR2_X1 U840 ( .A1(KEYINPUT33), .A2(n748), .ZN(n749) );
  NAND2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n758) );
  INV_X1 U842 ( .A(KEYINPUT101), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n753), .A2(KEYINPUT33), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n753), .A2(KEYINPUT101), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U847 ( .A1(n812), .A2(n756), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n892), .A2(G105), .ZN(n760) );
  XNOR2_X1 U850 ( .A(n760), .B(KEYINPUT38), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G129), .A2(n897), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G117), .A2(n896), .ZN(n763) );
  XNOR2_X1 U854 ( .A(KEYINPUT89), .B(n763), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n766), .B(KEYINPUT90), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G141), .A2(n516), .ZN(n767) );
  NAND2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n909) );
  NOR2_X1 U859 ( .A1(G1996), .A2(n909), .ZN(n924) );
  NAND2_X1 U860 ( .A1(G95), .A2(n892), .ZN(n770) );
  NAND2_X1 U861 ( .A1(G131), .A2(n516), .ZN(n769) );
  NAND2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G107), .A2(n896), .ZN(n772) );
  NAND2_X1 U864 ( .A1(G119), .A2(n897), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  OR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n884) );
  AND2_X1 U867 ( .A1(n884), .A2(G1991), .ZN(n776) );
  AND2_X1 U868 ( .A1(G1996), .A2(n909), .ZN(n775) );
  NOR2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n936) );
  INV_X1 U870 ( .A(n777), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n786) );
  NOR2_X1 U872 ( .A1(n936), .A2(n786), .ZN(n818) );
  NOR2_X1 U873 ( .A1(G1986), .A2(G290), .ZN(n780) );
  NOR2_X1 U874 ( .A1(G1991), .A2(n884), .ZN(n930) );
  NOR2_X1 U875 ( .A1(n780), .A2(n930), .ZN(n781) );
  NOR2_X1 U876 ( .A1(n818), .A2(n781), .ZN(n782) );
  XOR2_X1 U877 ( .A(KEYINPUT103), .B(n782), .Z(n783) );
  NOR2_X1 U878 ( .A1(n924), .A2(n783), .ZN(n784) );
  XNOR2_X1 U879 ( .A(KEYINPUT39), .B(n784), .ZN(n785) );
  XNOR2_X1 U880 ( .A(n785), .B(KEYINPUT104), .ZN(n799) );
  INV_X1 U881 ( .A(n786), .ZN(n821) );
  XNOR2_X1 U882 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n790) );
  NAND2_X1 U883 ( .A1(G104), .A2(n892), .ZN(n788) );
  NAND2_X1 U884 ( .A1(G140), .A2(n516), .ZN(n787) );
  NAND2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U886 ( .A(n790), .B(n789), .ZN(n796) );
  XNOR2_X1 U887 ( .A(KEYINPUT35), .B(KEYINPUT87), .ZN(n794) );
  NAND2_X1 U888 ( .A1(G116), .A2(n896), .ZN(n792) );
  NAND2_X1 U889 ( .A1(G128), .A2(n897), .ZN(n791) );
  NAND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U891 ( .A(n794), .B(n793), .ZN(n795) );
  NOR2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U893 ( .A(n797), .B(KEYINPUT36), .ZN(n798) );
  XNOR2_X1 U894 ( .A(n798), .B(KEYINPUT88), .ZN(n905) );
  XNOR2_X1 U895 ( .A(G2067), .B(KEYINPUT37), .ZN(n801) );
  NOR2_X1 U896 ( .A1(n905), .A2(n801), .ZN(n934) );
  NAND2_X1 U897 ( .A1(n821), .A2(n934), .ZN(n820) );
  NAND2_X1 U898 ( .A1(n799), .A2(n820), .ZN(n800) );
  XOR2_X1 U899 ( .A(KEYINPUT105), .B(n800), .Z(n802) );
  NAND2_X1 U900 ( .A1(n905), .A2(n801), .ZN(n938) );
  NAND2_X1 U901 ( .A1(n802), .A2(n938), .ZN(n803) );
  AND2_X1 U902 ( .A1(n803), .A2(n821), .ZN(n825) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n804) );
  XOR2_X1 U904 ( .A(n804), .B(KEYINPUT24), .Z(n805) );
  NOR2_X1 U905 ( .A1(n812), .A2(n805), .ZN(n806) );
  XOR2_X1 U906 ( .A(KEYINPUT91), .B(n806), .Z(n807) );
  NOR2_X1 U907 ( .A1(n825), .A2(n807), .ZN(n815) );
  NOR2_X1 U908 ( .A1(G2090), .A2(G303), .ZN(n808) );
  NAND2_X1 U909 ( .A1(G8), .A2(n808), .ZN(n809) );
  XNOR2_X1 U910 ( .A(n809), .B(KEYINPUT102), .ZN(n811) );
  NAND2_X1 U911 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n815), .A2(n814), .ZN(n816) );
  INV_X1 U914 ( .A(n818), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n823) );
  XNOR2_X1 U916 ( .A(G1986), .B(G290), .ZN(n979) );
  AND2_X1 U917 ( .A1(n979), .A2(n821), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  OR2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(KEYINPUT40), .B(n828), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U923 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n831) );
  XOR2_X1 U925 ( .A(KEYINPUT109), .B(n831), .Z(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U927 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  NOR2_X1 U928 ( .A1(n835), .A2(n834), .ZN(G325) );
  XNOR2_X1 U929 ( .A(KEYINPUT111), .B(G325), .ZN(G261) );
  XNOR2_X1 U930 ( .A(G108), .B(KEYINPUT121), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U933 ( .A(G2454), .B(G2451), .ZN(n844) );
  XNOR2_X1 U934 ( .A(G2430), .B(G2446), .ZN(n842) );
  XOR2_X1 U935 ( .A(G2435), .B(G2427), .Z(n837) );
  XNOR2_X1 U936 ( .A(KEYINPUT106), .B(G2438), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U938 ( .A(n838), .B(G2443), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1341), .B(G1348), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n845) );
  NAND2_X1 U943 ( .A1(n845), .A2(G14), .ZN(n846) );
  XOR2_X1 U944 ( .A(KEYINPUT107), .B(n846), .Z(n916) );
  XOR2_X1 U945 ( .A(KEYINPUT108), .B(n916), .Z(G401) );
  INV_X1 U946 ( .A(n847), .ZN(G319) );
  XNOR2_X1 U947 ( .A(G1981), .B(KEYINPUT41), .ZN(n857) );
  XOR2_X1 U948 ( .A(G1956), .B(G1961), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1966), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(G1971), .B(G1976), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT114), .B(G2474), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(G229) );
  XOR2_X1 U958 ( .A(G2678), .B(KEYINPUT43), .Z(n859) );
  XNOR2_X1 U959 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2090), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(G2096), .B(G2100), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U967 ( .A(G2078), .B(G2084), .Z(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(G227) );
  NAND2_X1 U969 ( .A1(G100), .A2(n892), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G112), .A2(n896), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G124), .A2(n897), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(KEYINPUT44), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G136), .A2(n516), .ZN(n871) );
  XOR2_X1 U975 ( .A(KEYINPUT115), .B(n871), .Z(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G118), .A2(n896), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G130), .A2(n897), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G106), .A2(n892), .ZN(n879) );
  NAND2_X1 U982 ( .A1(G142), .A2(n516), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n880), .Z(n881) );
  NOR2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(n884), .B(n883), .Z(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT116), .B(KEYINPUT119), .Z(n886) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n927), .B(n889), .ZN(n904) );
  NAND2_X1 U992 ( .A1(G139), .A2(n516), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n891), .B(KEYINPUT118), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G103), .A2(n892), .ZN(n893) );
  XOR2_X1 U995 ( .A(KEYINPUT117), .B(n893), .Z(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U997 ( .A1(G115), .A2(n896), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G127), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n940) );
  XNOR2_X1 U1002 ( .A(n940), .B(G162), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G160), .B(G164), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1007 ( .A(n910), .B(n909), .Z(n911) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n911), .ZN(G395) );
  XOR2_X1 U1009 ( .A(G286), .B(n983), .Z(n913) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(n914), .B(G171), .Z(n915) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n915), .ZN(G397) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n917), .B(KEYINPUT49), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT120), .B(n920), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n925), .Z(n932) );
  XNOR2_X1 U1025 ( .A(G160), .B(G2084), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(KEYINPUT122), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n937), .B(KEYINPUT123), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1034 ( .A(G2072), .B(n940), .Z(n942) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n943), .Z(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(KEYINPUT52), .B(n946), .ZN(n948) );
  INV_X1 U1040 ( .A(KEYINPUT55), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(n949), .A2(G29), .ZN(n1024) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n963) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G1991), .B(G25), .ZN(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n957) );
  XOR2_X1 U1047 ( .A(G32), .B(G1996), .Z(n952) );
  NAND2_X1 U1048 ( .A1(n952), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(KEYINPUT124), .B(G2072), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(G33), .B(n953), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(G27), .B(n958), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n964) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n964), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1060 ( .A(KEYINPUT55), .B(n967), .Z(n969) );
  INV_X1 U1061 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n970), .ZN(n1022) );
  INV_X1 U1064 ( .A(G16), .ZN(n1018) );
  XOR2_X1 U1065 ( .A(n1018), .B(KEYINPUT56), .Z(n994) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G168), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n973), .B(KEYINPUT57), .ZN(n992) );
  XOR2_X1 U1069 ( .A(G299), .B(G1956), .Z(n977) );
  AND2_X1 U1070 ( .A1(G303), .A2(G1971), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT125), .ZN(n988) );
  XOR2_X1 U1076 ( .A(G1348), .B(n983), .Z(n986) );
  XNOR2_X1 U1077 ( .A(G1341), .B(n984), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n990) );
  XOR2_X1 U1080 ( .A(G1961), .B(G171), .Z(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n1020) );
  XNOR2_X1 U1084 ( .A(G1348), .B(KEYINPUT59), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(G4), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G1981), .B(G6), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G19), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G20), .B(G1956), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1002), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G1961), .B(G5), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1007), .ZN(n1015) );
  XOR2_X1 U1098 ( .A(G1986), .B(G24), .Z(n1011) );
  XNOR2_X1 U1099 ( .A(G1976), .B(G23), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1012), .Z(n1013) );
  XNOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1025), .ZN(G150) );
  INV_X1 U1112 ( .A(G150), .ZN(G311) );
endmodule

