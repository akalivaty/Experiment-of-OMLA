//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT68), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G219), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n452), .B(new_n453), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n472), .C1(new_n466), .C2(new_n467), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n472), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  INV_X1    g054(.A(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G124), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n485), .A2(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n466), .B2(new_n467), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n499), .B(new_n502), .C1(new_n467), .C2(new_n466), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(G543), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n518), .A2(new_n508), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n510), .A2(new_n511), .A3(new_n517), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n514), .A2(new_n519), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND4_X1  g099(.A1(new_n510), .A2(G51), .A3(G543), .A4(new_n511), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n529), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n517), .A2(new_n526), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n525), .B(new_n531), .C1(new_n520), .C2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n513), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n508), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n521), .A2(G90), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(G171));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n515), .B2(new_n516), .ZN(new_n542));
  AND2_X1   g117(.A1(G68), .A2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(G651), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n510), .A2(G81), .A3(new_n517), .A4(new_n511), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n510), .A2(G43), .A3(G543), .A4(new_n511), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n512), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n507), .A2(new_n509), .B1(new_n506), .B2(G651), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n555), .A2(new_n556), .A3(G53), .A4(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT5), .B(G543), .Z(new_n560));
  XNOR2_X1  g135(.A(KEYINPUT74), .B(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n521), .A2(G91), .B1(new_n562), .B2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(G299));
  NAND3_X1  g139(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(G301));
  NAND3_X1  g140(.A1(new_n555), .A2(G49), .A3(G543), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n510), .A2(G87), .A3(new_n517), .A4(new_n511), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n555), .A2(G86), .A3(new_n517), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n555), .A2(G48), .A3(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n515), .B2(new_n516), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n573), .A3(new_n577), .ZN(G305));
  XOR2_X1   g153(.A(KEYINPUT76), .B(G47), .Z(new_n579));
  NAND2_X1  g154(.A1(new_n513), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n508), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n521), .A2(G85), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n520), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n555), .A2(KEYINPUT10), .A3(G92), .A4(new_n517), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT77), .B(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n560), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n513), .A2(G54), .B1(new_n593), .B2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n585), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n585), .B1(new_n596), .B2(G868), .ZN(G321));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G286), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g175(.A(G299), .B(KEYINPUT78), .Z(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(G297));
  AOI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(G280));
  INV_X1    g178(.A(G860), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n595), .B1(G559), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT79), .Z(G148));
  NAND3_X1  g181(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n599), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n595), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g186(.A(KEYINPUT3), .B(G2104), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n474), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g190(.A(G2100), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n482), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n489), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n472), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n617), .A2(new_n618), .A3(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT81), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  AND2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  OR3_X1    g213(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n638), .B1(new_n634), .B2(new_n635), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT82), .ZN(new_n653));
  XOR2_X1   g228(.A(G2096), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n649), .A2(new_n650), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT83), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n655), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1981), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT84), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G11), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT95), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n684), .A2(G28), .ZN(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n684), .B2(G28), .ZN(new_n687));
  OAI221_X1 g262(.A(new_n683), .B1(new_n685), .B2(new_n687), .C1(new_n623), .C2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(G2084), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n686), .B1(KEYINPUT24), .B2(G34), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(KEYINPUT24), .B2(G34), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n478), .B2(G29), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n688), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(G33), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n482), .A2(G139), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT93), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n612), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(new_n472), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n694), .B1(new_n704), .B2(new_n686), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n693), .B1(new_n689), .B2(new_n692), .C1(new_n705), .C2(G2072), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n686), .A2(G32), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n489), .A2(G129), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT94), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n474), .A2(G105), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT26), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n711), .B(new_n713), .C1(G141), .C2(new_n482), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n707), .B1(new_n716), .B2(new_n686), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT27), .B(G1996), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n686), .A2(G27), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT96), .ZN(new_n723));
  INV_X1    g298(.A(G164), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2078), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n720), .A2(new_n721), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n706), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G21), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G168), .B2(new_n729), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G1966), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n729), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1961), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G19), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n547), .B2(G16), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT90), .B(G1341), .Z(new_n738));
  OAI21_X1  g313(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n732), .B(new_n739), .C1(G2072), .C2(new_n705), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n734), .A2(G1961), .B1(G1966), .B2(new_n731), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n729), .A2(G20), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT23), .Z(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G299), .B2(G16), .ZN(new_n744));
  INV_X1    g319(.A(G1956), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n741), .B(new_n746), .C1(new_n737), .C2(new_n738), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n728), .A2(new_n740), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n596), .A2(G16), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G4), .B2(G16), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(KEYINPUT89), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(KEYINPUT89), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G1348), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n686), .A2(G35), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G162), .B2(new_n686), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n482), .A2(G140), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n489), .A2(G128), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n472), .A2(G116), .ZN(new_n761));
  OAI21_X1  g336(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n759), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G29), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n686), .A2(G26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT91), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(G2067), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(G2067), .ZN(new_n770));
  AOI22_X1  g345(.A1(G2090), .A2(new_n758), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n758), .A2(G2090), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n751), .A2(G1348), .A3(new_n752), .ZN(new_n773));
  AND4_X1   g348(.A1(new_n755), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n748), .A2(new_n774), .A3(KEYINPUT97), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n728), .A2(new_n740), .A3(new_n747), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n755), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n781));
  MUX2_X1   g356(.A(G24), .B(G290), .S(G16), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(KEYINPUT86), .ZN(new_n784));
  INV_X1    g359(.A(G1986), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n782), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT86), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G25), .A2(G29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n482), .A2(G131), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n489), .A2(G119), .ZN(new_n791));
  OR2_X1    g366(.A1(G95), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT85), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT35), .B(G1991), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n784), .A2(new_n788), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G23), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT87), .Z(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n569), .B2(new_n729), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT33), .ZN(new_n803));
  INV_X1    g378(.A(G1976), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n729), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n729), .ZN(new_n807));
  INV_X1    g382(.A(G1971), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G6), .B(G305), .S(G16), .Z(new_n810));
  XOR2_X1   g385(.A(KEYINPUT32), .B(G1981), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n805), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n805), .A2(new_n809), .A3(new_n815), .A4(new_n812), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n799), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n817), .A2(KEYINPUT88), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(KEYINPUT88), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n799), .A2(new_n820), .A3(new_n814), .A4(new_n816), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n818), .A2(KEYINPUT88), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n780), .B(new_n781), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n775), .A2(new_n779), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n823), .B1(new_n819), .B2(new_n821), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT98), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n824), .A2(new_n827), .ZN(G311));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n780), .B(new_n829), .C1(new_n822), .C2(new_n823), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT99), .B1(new_n825), .B2(new_n826), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(G150));
  NAND2_X1  g407(.A1(new_n596), .A2(G559), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT38), .Z(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n515), .B2(new_n516), .ZN(new_n836));
  AND2_X1   g411(.A1(G80), .A2(G543), .ZN(new_n837));
  OAI21_X1  g412(.A(G651), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n510), .A2(G93), .A3(new_n517), .A4(new_n511), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n510), .A2(G55), .A3(G543), .A4(new_n511), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n547), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n607), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n834), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n604), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n843), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(new_n715), .B(new_n763), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(new_n724), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n724), .ZN(new_n855));
  INV_X1    g430(.A(new_n704), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT100), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(KEYINPUT100), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n794), .B(new_n614), .ZN(new_n861));
  AOI22_X1  g436(.A1(G130), .A2(new_n489), .B1(new_n482), .B2(G142), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n472), .A2(KEYINPUT101), .A3(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT101), .B1(new_n472), .B2(G118), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n862), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n861), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n859), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n868), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n860), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n867), .B1(new_n860), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n623), .B(new_n478), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(G162), .Z(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n870), .B2(new_n871), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n842), .A2(new_n880), .A3(new_n844), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n842), .B2(new_n844), .ZN(new_n883));
  OAI22_X1  g458(.A1(new_n882), .A2(new_n883), .B1(G559), .B2(new_n595), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n609), .A3(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(G299), .A2(new_n595), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n558), .A2(new_n590), .A3(new_n563), .A4(new_n594), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(KEYINPUT41), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT41), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n893), .A3(KEYINPUT103), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n889), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT103), .B1(new_n887), .B2(new_n893), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n896), .A2(KEYINPUT105), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT105), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  XNOR2_X1  g474(.A(G303), .B(new_n569), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(G305), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT104), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT42), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n898), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n896), .A2(new_n897), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n907), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  OAI21_X1  g484(.A(G868), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n843), .A2(new_n599), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(G295));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n910), .A2(new_n913), .A3(new_n911), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n910), .B2(new_n911), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  INV_X1    g492(.A(new_n895), .ZN(new_n918));
  INV_X1    g493(.A(new_n844), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n607), .A2(new_n843), .ZN(new_n920));
  OAI21_X1  g495(.A(G171), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n842), .A2(G301), .A3(new_n844), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n921), .A2(G168), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G168), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n842), .A2(G301), .A3(new_n844), .ZN(new_n926));
  AOI21_X1  g501(.A(G301), .B1(new_n842), .B2(new_n844), .ZN(new_n927));
  OAI21_X1  g502(.A(G286), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n895), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n921), .A2(G168), .A3(new_n922), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n890), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n902), .A2(new_n903), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n902), .A2(new_n903), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n925), .A3(new_n932), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT107), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n933), .B2(new_n934), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n936), .B1(new_n942), .B2(new_n939), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI211_X1 g519(.A(KEYINPUT107), .B(new_n936), .C1(new_n942), .C2(new_n939), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n917), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n943), .B2(KEYINPUT108), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n948), .B(new_n936), .C1(new_n942), .C2(new_n939), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT44), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n946), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n946), .B2(new_n950), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(G397));
  INV_X1    g529(.A(KEYINPUT127), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  INV_X1    g531(.A(new_n503), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n502), .B1(new_n612), .B2(new_n499), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(new_n497), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n612), .A2(G125), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n472), .B1(new_n962), .B2(new_n465), .ZN(new_n963));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n963), .A2(new_n964), .A3(new_n476), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G2067), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n763), .B(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n716), .A2(G1996), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n716), .A2(G1996), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n794), .A2(new_n797), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n794), .A2(new_n797), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT110), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(G290), .B(new_n785), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n966), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n471), .A2(new_n477), .A3(G40), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n960), .B2(new_n961), .ZN(new_n981));
  OAI211_X1 g556(.A(KEYINPUT45), .B(new_n956), .C1(new_n959), .C2(new_n497), .ZN(new_n982));
  AOI21_X1  g557(.A(G1971), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n985), .B(new_n956), .C1(new_n959), .C2(new_n497), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT112), .B(G2090), .Z(new_n987));
  NAND4_X1  g562(.A1(new_n984), .A2(new_n986), .A3(new_n965), .A4(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n979), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n501), .A2(new_n503), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n492), .A2(new_n496), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n965), .B1(new_n993), .B2(KEYINPUT45), .ZN(new_n994));
  NOR3_X1   g569(.A1(G164), .A2(new_n961), .A3(G1384), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n808), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(KEYINPUT116), .A3(new_n988), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n990), .A2(G8), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(G303), .A2(G8), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT55), .Z(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n961), .B1(G164), .B2(G1384), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n965), .A3(new_n982), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n988), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(new_n1000), .A3(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G305), .A2(G1981), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n573), .A2(new_n572), .A3(new_n1011), .A4(new_n577), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n965), .B2(new_n993), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1010), .A2(KEYINPUT49), .A3(new_n1012), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n569), .B2(new_n804), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n567), .A2(new_n568), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(KEYINPUT113), .A3(G1976), .A4(new_n566), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1017), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n570), .B2(G1976), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(new_n1024), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n982), .A2(KEYINPUT117), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n993), .A2(new_n1032), .A3(KEYINPUT45), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n981), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1966), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n984), .A2(new_n965), .A3(new_n986), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1034), .A2(new_n1035), .B1(new_n1036), .B2(new_n689), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1037), .A2(new_n1016), .A3(G286), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1002), .A2(new_n1009), .A3(new_n1030), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT63), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1028), .A2(new_n1024), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1042), .A2(KEYINPUT114), .A3(new_n1019), .A4(new_n1025), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1008), .A2(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1001), .ZN(new_n1048));
  NOR4_X1   g623(.A1(new_n1037), .A2(new_n1040), .A3(new_n1016), .A4(G286), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1046), .A2(new_n1009), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1041), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G286), .A2(G8), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT51), .B1(new_n1054), .B2(KEYINPUT124), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1054), .B(new_n1055), .C1(new_n1037), .C2(new_n1016), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1052), .B(KEYINPUT123), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1033), .A2(new_n965), .A3(new_n1005), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n995), .A2(new_n1032), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1035), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1036), .A2(new_n689), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1057), .B1(new_n1062), .B2(G8), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1057), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n1037), .B2(new_n1054), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1056), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1009), .A2(new_n1030), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n996), .A2(new_n988), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1016), .B1(new_n1072), .B2(new_n979), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1000), .B1(new_n1073), .B2(new_n997), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n981), .A2(new_n1031), .A3(new_n1076), .A4(new_n1033), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT125), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(KEYINPUT53), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1006), .B2(G2078), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n984), .A2(new_n965), .A3(new_n986), .ZN(new_n1085));
  INV_X1    g660(.A(G1961), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(G301), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT62), .B(new_n1056), .C1(new_n1063), .C2(new_n1067), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1070), .A2(new_n1075), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1009), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(G288), .B2(G1976), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n570), .A2(KEYINPUT115), .A3(new_n804), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1012), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1093), .B1(new_n1017), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1051), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n477), .A2(KEYINPUT53), .A3(G40), .A4(new_n1076), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n470), .A2(KEYINPUT126), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n472), .B1(new_n470), .B2(KEYINPUT126), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n982), .A3(new_n1005), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1084), .A2(new_n1087), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G171), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1082), .A2(new_n1089), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT54), .B(new_n1108), .C1(new_n1109), .C2(G171), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1068), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1110), .A2(new_n1075), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(G2072), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n981), .A2(new_n982), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1085), .A2(new_n745), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n558), .B(new_n563), .C1(new_n1118), .C2(KEYINPUT57), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n563), .B2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G299), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1119), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1085), .A2(new_n754), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n965), .A2(new_n993), .A3(new_n967), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n596), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(KEYINPUT60), .A3(new_n1126), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n596), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n595), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n1127), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1122), .A2(KEYINPUT121), .A3(new_n1124), .A4(KEYINPUT61), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(G1341), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n960), .B2(new_n980), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1006), .B2(G1996), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT59), .B1(new_n1142), .B2(new_n547), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1123), .B1(new_n1116), .B2(new_n1115), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(KEYINPUT59), .A3(new_n547), .ZN(new_n1147));
  NAND2_X1  g722(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1123), .A2(new_n1116), .A3(new_n1115), .A4(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1138), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1122), .B(new_n1128), .C1(new_n1137), .C2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1107), .A2(G171), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1090), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1112), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n978), .B1(new_n1101), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n976), .A2(new_n966), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT48), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n763), .A2(G2067), .ZN(new_n1160));
  INV_X1    g735(.A(new_n971), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(new_n972), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n1157), .A2(new_n1159), .B1(new_n1162), .B2(new_n966), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n966), .A2(G1996), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT46), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n966), .B1(new_n716), .B2(new_n968), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT47), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n955), .B1(new_n1156), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1128), .A2(new_n1122), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1127), .A2(new_n1136), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1150), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1172), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1154), .A2(new_n1110), .A3(new_n1075), .A4(new_n1111), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1051), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(KEYINPUT127), .B(new_n1169), .C1(new_n1181), .C2(new_n978), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1171), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g758(.A1(new_n463), .A2(G227), .ZN(new_n1185));
  NAND3_X1  g759(.A1(new_n680), .A2(new_n646), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1186), .B1(new_n875), .B2(new_n877), .ZN(new_n1187));
  INV_X1    g761(.A(new_n945), .ZN(new_n1188));
  INV_X1    g762(.A(new_n944), .ZN(new_n1189));
  AND3_X1   g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(G308));
  NAND3_X1  g764(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(G225));
endmodule


