

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U321 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n378) );
  XNOR2_X1 U322 ( .A(n379), .B(n378), .ZN(n402) );
  XOR2_X1 U323 ( .A(G99GAT), .B(G85GAT), .Z(n346) );
  NOR2_X1 U324 ( .A1(n407), .A2(n405), .ZN(n406) );
  XNOR2_X1 U325 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U326 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U327 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U328 ( .A(n345), .B(n344), .ZN(n407) );
  NOR2_X1 U329 ( .A1(n539), .A2(n451), .ZN(n566) );
  XOR2_X1 U330 ( .A(n324), .B(n323), .Z(n534) );
  XNOR2_X1 U331 ( .A(n452), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U332 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(G120GAT), .B(G71GAT), .Z(n357) );
  XOR2_X1 U334 ( .A(G127GAT), .B(KEYINPUT0), .Z(n290) );
  XNOR2_X1 U335 ( .A(G113GAT), .B(G134GAT), .ZN(n289) );
  XNOR2_X1 U336 ( .A(n290), .B(n289), .ZN(n314) );
  XOR2_X1 U337 ( .A(n357), .B(n314), .Z(n292) );
  NAND2_X1 U338 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U339 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U340 ( .A(n293), .B(G176GAT), .Z(n297) );
  XOR2_X1 U341 ( .A(G183GAT), .B(KEYINPUT17), .Z(n295) );
  XNOR2_X1 U342 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n424) );
  XNOR2_X1 U344 ( .A(n424), .B(KEYINPUT85), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n305) );
  XOR2_X1 U346 ( .A(G190GAT), .B(G99GAT), .Z(n299) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(G43GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U349 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n301) );
  XNOR2_X1 U350 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U352 ( .A(n303), .B(n302), .Z(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n539) );
  XOR2_X1 U354 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n324) );
  XOR2_X1 U357 ( .A(KEYINPUT90), .B(G148GAT), .Z(n309) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(G120GAT), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U360 ( .A(G29GAT), .B(G85GAT), .Z(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n320) );
  XOR2_X1 U362 ( .A(G155GAT), .B(KEYINPUT2), .Z(n313) );
  XNOR2_X1 U363 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n433) );
  XNOR2_X1 U365 ( .A(n314), .B(n433), .ZN(n318) );
  XOR2_X1 U366 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n316) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(G57GAT), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n322) );
  NAND2_X1 U371 ( .A1(G225GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  INV_X1 U373 ( .A(KEYINPUT76), .ZN(n325) );
  NAND2_X1 U374 ( .A1(G190GAT), .A2(n325), .ZN(n328) );
  INV_X1 U375 ( .A(G190GAT), .ZN(n326) );
  NAND2_X1 U376 ( .A1(n326), .A2(KEYINPUT76), .ZN(n327) );
  NAND2_X1 U377 ( .A1(n328), .A2(n327), .ZN(n417) );
  XOR2_X1 U378 ( .A(KEYINPUT9), .B(n417), .Z(n330) );
  XNOR2_X1 U379 ( .A(G218GAT), .B(n346), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n336) );
  XOR2_X1 U381 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n332) );
  XNOR2_X1 U382 ( .A(G36GAT), .B(KEYINPUT10), .ZN(n331) );
  XOR2_X1 U383 ( .A(n332), .B(n331), .Z(n334) );
  NAND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  XOR2_X1 U385 ( .A(n337), .B(G92GAT), .Z(n345) );
  XOR2_X1 U386 ( .A(G29GAT), .B(G43GAT), .Z(n339) );
  XNOR2_X1 U387 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n338) );
  XNOR2_X1 U388 ( .A(n339), .B(n338), .ZN(n366) );
  XNOR2_X1 U389 ( .A(n366), .B(G106GAT), .ZN(n343) );
  XOR2_X1 U390 ( .A(KEYINPUT65), .B(G162GAT), .Z(n341) );
  XNOR2_X1 U391 ( .A(G50GAT), .B(G134GAT), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT13), .Z(n383) );
  XNOR2_X1 U394 ( .A(n346), .B(n383), .ZN(n348) );
  AND2_X1 U395 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U396 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U397 ( .A(KEYINPUT69), .B(KEYINPUT33), .Z(n350) );
  XNOR2_X1 U398 ( .A(KEYINPUT31), .B(KEYINPUT70), .ZN(n349) );
  XNOR2_X1 U399 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U400 ( .A(n352), .B(n351), .Z(n359) );
  INV_X1 U401 ( .A(G204GAT), .ZN(n356) );
  XOR2_X1 U402 ( .A(G92GAT), .B(G64GAT), .Z(n354) );
  XNOR2_X1 U403 ( .A(G176GAT), .B(KEYINPUT72), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U405 ( .A(n356), .B(n355), .ZN(n416) );
  XNOR2_X1 U406 ( .A(n357), .B(n416), .ZN(n358) );
  XNOR2_X1 U407 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U408 ( .A(n360), .B(KEYINPUT32), .ZN(n364) );
  XOR2_X1 U409 ( .A(G78GAT), .B(G148GAT), .Z(n362) );
  XNOR2_X1 U410 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n361) );
  XNOR2_X1 U411 ( .A(n362), .B(n361), .ZN(n442) );
  XOR2_X1 U412 ( .A(n442), .B(KEYINPUT73), .Z(n363) );
  XNOR2_X1 U413 ( .A(n364), .B(n363), .ZN(n575) );
  XNOR2_X1 U414 ( .A(n575), .B(KEYINPUT41), .ZN(n455) );
  XNOR2_X1 U415 ( .A(G15GAT), .B(G1GAT), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n365), .B(KEYINPUT67), .ZN(n387) );
  XOR2_X1 U417 ( .A(n366), .B(KEYINPUT29), .Z(n368) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U420 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n370) );
  XNOR2_X1 U421 ( .A(G113GAT), .B(G197GAT), .ZN(n369) );
  XNOR2_X1 U422 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U423 ( .A(n372), .B(n371), .Z(n376) );
  XNOR2_X1 U424 ( .A(G50GAT), .B(G22GAT), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n373), .B(G141GAT), .ZN(n445) );
  XNOR2_X1 U426 ( .A(G169GAT), .B(G36GAT), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n374), .B(G8GAT), .ZN(n425) );
  XNOR2_X1 U428 ( .A(n445), .B(n425), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n387), .B(n377), .ZN(n570) );
  NAND2_X1 U431 ( .A1(n455), .A2(n570), .ZN(n379) );
  XOR2_X1 U432 ( .A(G211GAT), .B(G127GAT), .Z(n381) );
  XNOR2_X1 U433 ( .A(G183GAT), .B(G71GAT), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U435 ( .A(n383), .B(n382), .Z(n385) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U438 ( .A(n386), .B(KEYINPUT82), .Z(n389) );
  XNOR2_X1 U439 ( .A(n387), .B(KEYINPUT81), .ZN(n388) );
  XNOR2_X1 U440 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U441 ( .A(G64GAT), .B(G155GAT), .Z(n391) );
  XNOR2_X1 U442 ( .A(G22GAT), .B(G78GAT), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U444 ( .A(n393), .B(n392), .Z(n401) );
  XOR2_X1 U445 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n395) );
  XNOR2_X1 U446 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U448 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n397) );
  XNOR2_X1 U449 ( .A(G8GAT), .B(KEYINPUT78), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n544) );
  NAND2_X1 U453 ( .A1(n402), .A2(n544), .ZN(n404) );
  INV_X1 U454 ( .A(KEYINPUT113), .ZN(n403) );
  XNOR2_X1 U455 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U456 ( .A(n406), .B(KEYINPUT47), .ZN(n413) );
  XOR2_X1 U457 ( .A(KEYINPUT36), .B(n407), .Z(n583) );
  NOR2_X1 U458 ( .A1(n544), .A2(n583), .ZN(n408) );
  XNOR2_X1 U459 ( .A(KEYINPUT45), .B(n408), .ZN(n409) );
  AND2_X1 U460 ( .A1(n409), .A2(n575), .ZN(n410) );
  XNOR2_X1 U461 ( .A(n410), .B(KEYINPUT114), .ZN(n411) );
  XOR2_X1 U462 ( .A(KEYINPUT68), .B(n570), .Z(n463) );
  NAND2_X1 U463 ( .A1(n411), .A2(n463), .ZN(n412) );
  NAND2_X1 U464 ( .A1(n413), .A2(n412), .ZN(n415) );
  XOR2_X1 U465 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n414) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n536) );
  XOR2_X1 U467 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U469 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U470 ( .A(KEYINPUT88), .B(G218GAT), .Z(n421) );
  XNOR2_X1 U471 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n420) );
  XNOR2_X1 U472 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U473 ( .A(G197GAT), .B(n422), .Z(n444) );
  XOR2_X1 U474 ( .A(n423), .B(n444), .Z(n427) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n427), .B(n426), .ZN(n525) );
  XNOR2_X1 U477 ( .A(n525), .B(KEYINPUT119), .ZN(n428) );
  NOR2_X1 U478 ( .A1(n536), .A2(n428), .ZN(n431) );
  XNOR2_X1 U479 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n429) );
  XNOR2_X1 U480 ( .A(n429), .B(KEYINPUT54), .ZN(n430) );
  XNOR2_X1 U481 ( .A(n431), .B(n430), .ZN(n432) );
  NOR2_X1 U482 ( .A1(n534), .A2(n432), .ZN(n569) );
  XOR2_X1 U483 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n435) );
  XNOR2_X1 U484 ( .A(KEYINPUT86), .B(n433), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U486 ( .A(n436), .B(KEYINPUT23), .Z(n441) );
  XOR2_X1 U487 ( .A(KEYINPUT89), .B(KEYINPUT87), .Z(n438) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(G204GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U492 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U493 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U494 ( .A(n447), .B(n446), .ZN(n472) );
  NAND2_X1 U495 ( .A1(n569), .A2(n472), .ZN(n449) );
  XOR2_X1 U496 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n448) );
  XNOR2_X1 U497 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT55), .B(n450), .Z(n451) );
  NAND2_X1 U499 ( .A1(n566), .A2(n407), .ZN(n454) );
  XOR2_X1 U500 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n452) );
  BUF_X1 U501 ( .A(n455), .Z(n558) );
  NAND2_X1 U502 ( .A1(n566), .A2(n558), .ZN(n459) );
  XOR2_X1 U503 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n457) );
  XNOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n456) );
  XNOR2_X1 U505 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U506 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  XOR2_X1 U507 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n461) );
  XNOR2_X1 U508 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n460) );
  XNOR2_X1 U509 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U510 ( .A(KEYINPUT97), .B(n462), .Z(n484) );
  INV_X1 U511 ( .A(n463), .ZN(n564) );
  NAND2_X1 U512 ( .A1(n575), .A2(n564), .ZN(n464) );
  XNOR2_X1 U513 ( .A(n464), .B(KEYINPUT74), .ZN(n494) );
  NOR2_X1 U514 ( .A1(n544), .A2(n407), .ZN(n465) );
  XNOR2_X1 U515 ( .A(KEYINPUT16), .B(n465), .ZN(n482) );
  XNOR2_X1 U516 ( .A(n525), .B(KEYINPUT93), .ZN(n466) );
  XNOR2_X1 U517 ( .A(n466), .B(KEYINPUT27), .ZN(n474) );
  XOR2_X1 U518 ( .A(n472), .B(KEYINPUT28), .Z(n529) );
  NOR2_X1 U519 ( .A1(n474), .A2(n529), .ZN(n537) );
  NAND2_X1 U520 ( .A1(n539), .A2(n537), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n467), .A2(n534), .ZN(n480) );
  XOR2_X1 U522 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n471) );
  INV_X1 U523 ( .A(n539), .ZN(n527) );
  NAND2_X1 U524 ( .A1(n527), .A2(n525), .ZN(n468) );
  XOR2_X1 U525 ( .A(KEYINPUT95), .B(n468), .Z(n469) );
  NAND2_X1 U526 ( .A1(n469), .A2(n472), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n471), .B(n470), .ZN(n478) );
  NOR2_X1 U528 ( .A1(n472), .A2(n527), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n473), .B(KEYINPUT26), .ZN(n568) );
  INV_X1 U530 ( .A(n474), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n568), .A2(n475), .ZN(n552) );
  XOR2_X1 U532 ( .A(KEYINPUT94), .B(n552), .Z(n476) );
  NOR2_X1 U533 ( .A1(n534), .A2(n476), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U535 ( .A1(n480), .A2(n479), .ZN(n490) );
  INV_X1 U536 ( .A(n490), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n482), .A2(n481), .ZN(n508) );
  NOR2_X1 U538 ( .A1(n494), .A2(n508), .ZN(n488) );
  NAND2_X1 U539 ( .A1(n488), .A2(n534), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n484), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n488), .A2(n525), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U544 ( .A1(n488), .A2(n527), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NAND2_X1 U546 ( .A1(n488), .A2(n529), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U548 ( .A1(n583), .A2(n490), .ZN(n491) );
  NAND2_X1 U549 ( .A1(n544), .A2(n491), .ZN(n493) );
  XOR2_X1 U550 ( .A(KEYINPUT37), .B(KEYINPUT100), .Z(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n522) );
  NOR2_X1 U552 ( .A1(n494), .A2(n522), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT38), .ZN(n504) );
  NAND2_X1 U554 ( .A1(n534), .A2(n504), .ZN(n497) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n499) );
  NAND2_X1 U558 ( .A1(n525), .A2(n504), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n502) );
  NAND2_X1 U562 ( .A1(n527), .A2(n504), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n529), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(KEYINPUT104), .ZN(n506) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n510) );
  INV_X1 U569 ( .A(n570), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n507), .A2(n558), .ZN(n521) );
  NOR2_X1 U571 ( .A1(n521), .A2(n508), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n517), .A2(n534), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n517), .A2(n525), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n515) );
  NAND2_X1 U579 ( .A1(n517), .A2(n527), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U583 ( .A1(n517), .A2(n529), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U585 ( .A(G78GAT), .B(n520), .Z(G1335GAT) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n524) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n534), .A2(n530), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n530), .A2(n525), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n532) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  INV_X1 U598 ( .A(n534), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n550) );
  NAND2_X1 U600 ( .A1(n537), .A2(n550), .ZN(n538) );
  NOR2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n547), .A2(n564), .ZN(n540) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(n540), .Z(n541) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U606 ( .A1(n547), .A2(n558), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  INV_X1 U608 ( .A(n544), .ZN(n578) );
  NAND2_X1 U609 ( .A1(n578), .A2(n547), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U613 ( .A1(n547), .A2(n407), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  INV_X1 U615 ( .A(n550), .ZN(n551) );
  NOR2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n562), .A2(n570), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT116), .B(n553), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(KEYINPUT117), .B(n557), .Z(n560) );
  NAND2_X1 U624 ( .A1(n562), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n578), .A2(n562), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n407), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n566), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n578), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(KEYINPUT126), .B(KEYINPUT59), .ZN(n574) );
  XOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT60), .Z(n572) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n582) );
  INV_X1 U637 ( .A(n582), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n579), .A2(n570), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  OR2_X1 U642 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

