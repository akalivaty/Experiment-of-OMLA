//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n229), .B(new_n232), .C1(new_n220), .C2(new_n221), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n223), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n215), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G45), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n217), .B1(new_n257), .B2(KEYINPUT71), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(KEYINPUT71), .B2(new_n257), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n262), .A3(new_n251), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n215), .A2(G1698), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G226), .B2(G1698), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  OAI22_X1  g0072(.A1(new_n268), .A2(new_n271), .B1(new_n272), .B2(new_n202), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n274));
  INV_X1    g0074(.A(new_n226), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT67), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(new_n255), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n259), .A2(new_n266), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n281));
  XOR2_X1   g0081(.A(new_n281), .B(KEYINPUT72), .Z(new_n282));
  OR2_X1    g0082(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G179), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n281), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G169), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT14), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT14), .B1(new_n285), .B2(G169), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n284), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n275), .B1(KEYINPUT68), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT68), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n293), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT73), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n227), .A2(G33), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n299), .A2(new_n208), .B1(new_n227), .B2(G68), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n295), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT11), .ZN(new_n302));
  INV_X1    g0102(.A(G13), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G1), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G68), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT12), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n291), .A2(KEYINPUT68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n253), .A2(G20), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n308), .A2(new_n294), .A3(new_n226), .A4(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n216), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n307), .A2(KEYINPUT74), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT74), .B1(new_n307), .B2(new_n311), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n302), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n290), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n282), .A2(G190), .A3(new_n283), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n314), .B1(new_n285), .B2(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G226), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n272), .ZN(new_n321));
  NAND2_X1  g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G222), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G223), .A2(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(G77), .B2(new_n323), .ZN(new_n328));
  INV_X1    g0128(.A(new_n278), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n266), .B1(new_n319), .B2(new_n257), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G179), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n330), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n303), .A2(new_n227), .A3(G1), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(G50), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(G50), .B2(new_n310), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT69), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT8), .B(G58), .ZN(new_n338));
  INV_X1    g0138(.A(G150), .ZN(new_n339));
  INV_X1    g0139(.A(new_n296), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n338), .A2(new_n299), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G50), .A2(G58), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n227), .B1(new_n342), .B2(new_n216), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n295), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n333), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G179), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n271), .A2(new_n203), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G238), .A2(G1698), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n349), .B1(new_n215), .B2(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n278), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n275), .A2(new_n255), .B1(new_n252), .B2(new_n253), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(G244), .B1(new_n263), .B2(new_n265), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT70), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT70), .B1(new_n351), .B2(new_n353), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n347), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n351), .A2(new_n353), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT70), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n332), .A3(new_n354), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n362), .A2(new_n299), .B1(new_n227), .B2(new_n208), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n338), .A2(new_n340), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n295), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n310), .A2(new_n208), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n334), .A2(new_n208), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n357), .A2(new_n361), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(G190), .B1(new_n355), .B2(new_n356), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n360), .A2(G200), .A3(new_n354), .ZN(new_n372));
  INV_X1    g0172(.A(new_n368), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n346), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n315), .A2(new_n318), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT79), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n338), .A2(new_n334), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n310), .B2(new_n338), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT76), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n352), .A2(G232), .B1(new_n263), .B2(new_n265), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n319), .A2(G1698), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n384), .B1(G223), .B2(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G87), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n382), .B(new_n383), .C1(new_n387), .C2(new_n329), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n385), .A2(new_n386), .B1(new_n277), .B2(new_n274), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n266), .B1(new_n257), .B2(new_n215), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n214), .A2(new_n216), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n296), .A2(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n271), .B2(new_n227), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n216), .B1(new_n400), .B2(KEYINPUT75), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n321), .A2(new_n227), .A3(new_n322), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n321), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n322), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI211_X1 g0207(.A(new_n394), .B(new_n399), .C1(new_n401), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n216), .B1(new_n404), .B2(new_n406), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n394), .B1(new_n409), .B2(new_n399), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n295), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n381), .B(new_n393), .C1(new_n408), .C2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n378), .B1(new_n412), .B2(KEYINPUT17), .ZN(new_n413));
  INV_X1    g0213(.A(new_n412), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT79), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(KEYINPUT78), .ZN(new_n417));
  INV_X1    g0217(.A(new_n399), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n402), .A2(KEYINPUT75), .A3(new_n403), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G68), .ZN(new_n421));
  OAI211_X1 g0221(.A(KEYINPUT16), .B(new_n418), .C1(new_n419), .C2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(new_n295), .A3(new_n410), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT78), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n381), .A4(new_n393), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n413), .B(new_n416), .C1(new_n415), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n381), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT77), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT76), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n380), .B(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n295), .ZN(new_n433));
  INV_X1    g0233(.A(new_n406), .ZN(new_n434));
  OAI21_X1  g0234(.A(G68), .B1(new_n400), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n418), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n436), .B2(new_n394), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n432), .B1(new_n437), .B2(new_n422), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT77), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n390), .A2(new_n391), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(new_n332), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n441), .B2(G179), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT18), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  AND4_X1   g0245(.A1(KEYINPUT18), .A2(new_n430), .A3(new_n439), .A4(new_n444), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n427), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n345), .B(KEYINPUT9), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT10), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n330), .A2(G200), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n382), .B2(new_n330), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n448), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n449), .B1(new_n448), .B2(new_n452), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n377), .A2(new_n447), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(G107), .B1(new_n400), .B2(new_n434), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n204), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT80), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(KEYINPUT6), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n204), .A2(KEYINPUT80), .A3(new_n462), .A4(new_n458), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n202), .A2(KEYINPUT6), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n461), .A2(G20), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n296), .A2(G77), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n457), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n295), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n334), .B1(new_n253), .B2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(G97), .A3(new_n294), .A4(new_n292), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n334), .A2(new_n202), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n324), .A2(KEYINPUT4), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n323), .A2(G244), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n271), .A2(new_n209), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(KEYINPUT4), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n323), .A2(G250), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n324), .B1(new_n480), .B2(KEYINPUT4), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n278), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n253), .B(G45), .C1(new_n483), .C2(G41), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n260), .A2(new_n262), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n483), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n264), .B1(new_n275), .B2(new_n255), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT5), .B1(new_n260), .B2(new_n262), .ZN(new_n489));
  OAI211_X1 g0289(.A(G257), .B(new_n256), .C1(new_n489), .C2(new_n484), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n482), .A2(new_n347), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n482), .A2(new_n491), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n474), .B(new_n492), .C1(new_n493), .C2(G169), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n482), .A2(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G200), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n472), .B1(new_n467), .B2(new_n295), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n482), .A2(G190), .A3(new_n491), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT81), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n494), .A2(new_n499), .A3(KEYINPUT81), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  AOI21_X1  g0305(.A(G20), .B1(G33), .B2(G283), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n272), .A2(G97), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n506), .A2(new_n507), .B1(G20), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n295), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT20), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n305), .A2(G116), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n469), .A2(new_n294), .A3(new_n292), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G303), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n321), .A2(new_n518), .A3(new_n322), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n324), .A2(G257), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G264), .A2(G1698), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n269), .C2(new_n270), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n278), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G270), .B(new_n256), .C1(new_n489), .C2(new_n484), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n523), .A2(new_n488), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G169), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n505), .B1(new_n517), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(G200), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(G190), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n517), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n516), .A2(G179), .A3(new_n525), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n516), .A2(KEYINPUT21), .A3(G169), .A4(new_n526), .ZN(new_n533));
  AND4_X1   g0333(.A1(new_n528), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  XOR2_X1   g0334(.A(KEYINPUT85), .B(KEYINPUT22), .Z(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(new_n227), .A3(G87), .A4(new_n323), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n227), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n537));
  XNOR2_X1  g0337(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n227), .B2(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n272), .A2(new_n508), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n227), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n536), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT24), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n536), .A2(new_n547), .A3(new_n539), .A4(new_n544), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n433), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n305), .A2(G107), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT25), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n433), .A2(new_n469), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n203), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G250), .B(new_n324), .C1(new_n269), .C2(new_n270), .ZN(new_n555));
  OAI211_X1 g0355(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n556));
  INV_X1    g0356(.A(G294), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n556), .C1(new_n272), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n278), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT86), .ZN(new_n560));
  OAI211_X1 g0360(.A(G264), .B(new_n256), .C1(new_n489), .C2(new_n484), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n488), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT86), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n563), .A3(new_n278), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n560), .A2(new_n562), .A3(new_n382), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n559), .A2(new_n488), .A3(new_n561), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n389), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n554), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n566), .A2(new_n347), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(G169), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(new_n554), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT84), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n211), .B1(new_n251), .B2(G1), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n253), .A2(new_n264), .A3(G45), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n256), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G238), .A2(G1698), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n209), .B2(G1698), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n543), .B1(new_n579), .B2(new_n323), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n329), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n332), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G179), .B2(new_n581), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n323), .A2(new_n227), .A3(G68), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n299), .A2(new_n202), .ZN(new_n585));
  NAND3_X1  g0385(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n227), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT82), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n210), .A2(new_n202), .A3(new_n203), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n587), .A2(KEYINPUT82), .ZN(new_n591));
  OAI221_X1 g0391(.A(new_n584), .B1(KEYINPUT19), .B2(new_n585), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n295), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n362), .A2(new_n334), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n552), .B2(new_n362), .ZN(new_n597));
  INV_X1    g0397(.A(new_n362), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n514), .A2(KEYINPUT83), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n583), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n514), .A2(G87), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n593), .A2(new_n594), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n577), .ZN(new_n604));
  INV_X1    g0404(.A(new_n580), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n278), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G190), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n581), .A2(G200), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n574), .B1(new_n601), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n552), .A2(new_n596), .A3(new_n362), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT83), .B1(new_n514), .B2(new_n598), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n594), .B(new_n593), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n583), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n603), .A2(new_n609), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT84), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n573), .B1(new_n611), .B2(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n456), .A2(new_n504), .A3(new_n534), .A4(new_n619), .ZN(G372));
  NAND2_X1  g0420(.A1(new_n444), .A2(new_n428), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT18), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n318), .A2(new_n370), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n315), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n622), .B1(new_n624), .B2(new_n427), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n455), .B(KEYINPUT87), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n346), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n617), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n528), .A2(new_n532), .A3(new_n533), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n572), .A2(new_n554), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n499), .B(new_n569), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n630), .B1(new_n633), .B2(new_n494), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n494), .B1(new_n611), .B2(new_n618), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n616), .B1(new_n635), .B2(new_n629), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n456), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n628), .A2(new_n638), .ZN(G369));
  NAND2_X1  g0439(.A1(new_n304), .A2(new_n227), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(G213), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n516), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n534), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n631), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n646), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n573), .ZN(new_n651));
  INV_X1    g0451(.A(new_n645), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n554), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n632), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n652), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n648), .A2(new_n645), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n651), .B1(new_n632), .B2(new_n652), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(G399));
  OR2_X1    g0459(.A1(new_n589), .A2(G116), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT88), .ZN(new_n661));
  INV_X1    g0461(.A(new_n230), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n485), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G1), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n661), .A2(new_n665), .B1(new_n224), .B2(new_n664), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT29), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n668), .B(new_n652), .C1(new_n634), .C2(new_n636), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n569), .A2(new_n499), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n648), .B2(new_n654), .ZN(new_n671));
  INV_X1    g0471(.A(new_n494), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n672), .A2(new_n601), .A3(new_n610), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n601), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n601), .A2(new_n610), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .A3(new_n672), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n645), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n669), .B1(new_n678), .B2(new_n668), .ZN(new_n679));
  XOR2_X1   g0479(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n680));
  NOR2_X1   g0480(.A1(new_n652), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n559), .A2(new_n561), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT90), .B1(new_n682), .B2(new_n581), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT90), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n606), .A2(new_n684), .A3(new_n559), .A4(new_n561), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n523), .A2(new_n488), .A3(G179), .A4(new_n524), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT91), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n522), .A2(new_n519), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n689), .A2(new_n278), .B1(new_n486), .B2(new_n487), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT91), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(G179), .A4(new_n524), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n686), .A2(new_n493), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT92), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n686), .A2(new_n697), .A3(new_n493), .A4(new_n693), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n686), .A2(KEYINPUT30), .A3(new_n493), .A4(new_n693), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n606), .A2(G179), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n495), .A2(new_n526), .A3(new_n701), .A4(new_n566), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n681), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n619), .A2(new_n504), .A3(new_n534), .A4(new_n652), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n525), .A2(new_n606), .A3(G179), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(KEYINPUT93), .A3(new_n495), .A4(new_n566), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n700), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT30), .B1(new_n694), .B2(KEYINPUT92), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n698), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n652), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n704), .B(new_n705), .C1(new_n713), .C2(KEYINPUT31), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n679), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n667), .B1(new_n716), .B2(G1), .ZN(G364));
  NAND3_X1  g0517(.A1(new_n227), .A2(G13), .A3(G45), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n253), .B1(new_n718), .B2(KEYINPUT94), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n663), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n650), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n649), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n662), .A2(new_n271), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G355), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G116), .B2(new_n230), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n245), .A2(G45), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n662), .A2(new_n323), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n251), .B2(new_n225), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n727), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n226), .B1(G20), .B2(new_n332), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(KEYINPUT95), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n722), .B1(new_n732), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n227), .A2(new_n347), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n389), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n271), .B1(new_n746), .B2(G68), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n382), .A2(G179), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n227), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G97), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n227), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G107), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n382), .A2(new_n389), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n752), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G87), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n747), .A2(new_n751), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n743), .A2(new_n756), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n743), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G50), .A2(new_n762), .B1(new_n765), .B2(G77), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n743), .A2(G190), .A3(new_n389), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n214), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT32), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n752), .A2(new_n763), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n770), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(KEYINPUT32), .A3(G159), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n760), .B(new_n768), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT96), .Z(new_n776));
  OR2_X1    g0576(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G329), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n764), .A2(new_n782), .B1(new_n753), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n767), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n323), .B(new_n784), .C1(G322), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n750), .A2(G294), .ZN(new_n787));
  INV_X1    g0587(.A(G326), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n761), .A2(new_n788), .B1(new_n757), .B2(new_n518), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n746), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n781), .A2(new_n786), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n776), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n794));
  INV_X1    g0594(.A(new_n736), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n793), .B2(KEYINPUT98), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n742), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n739), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n649), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n724), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n637), .A2(new_n652), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n368), .A2(new_n645), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n369), .A2(new_n374), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT99), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n369), .A2(new_n374), .A3(KEYINPUT99), .A4(new_n803), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT101), .ZN(new_n809));
  OR3_X1    g0609(.A1(new_n369), .A2(KEYINPUT100), .A3(new_n652), .ZN(new_n810));
  OAI21_X1  g0610(.A(KEYINPUT100), .B1(new_n369), .B2(new_n652), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n809), .B1(new_n808), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n802), .B(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n715), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n722), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n780), .A2(G311), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n761), .A2(new_n518), .B1(new_n764), .B2(new_n508), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n323), .B(new_n821), .C1(G283), .C2(new_n746), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n767), .A2(new_n557), .B1(new_n753), .B2(new_n210), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G107), .B2(new_n758), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n820), .A2(new_n822), .A3(new_n751), .A4(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G137), .A2(new_n762), .B1(new_n746), .B2(G150), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n827), .B2(new_n767), .C1(new_n771), .C2(new_n764), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  INV_X1    g0629(.A(G50), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n757), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n323), .B1(new_n753), .B2(new_n216), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(G58), .C2(new_n750), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n779), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n825), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n736), .ZN(new_n837));
  INV_X1    g0637(.A(new_n722), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n736), .A2(new_n737), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n839), .B2(new_n208), .ZN(new_n840));
  INV_X1    g0640(.A(new_n815), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n837), .B(new_n840), .C1(new_n841), .C2(new_n738), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n819), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G384));
  NAND3_X1  g0644(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT35), .ZN(new_n846));
  OAI211_X1 g0646(.A(G116), .B(new_n228), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n846), .B2(new_n845), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT36), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n225), .B(G77), .C1(new_n214), .C2(new_n216), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n830), .A2(G68), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n253), .B(G13), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n622), .A2(new_n643), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  INV_X1    g0655(.A(new_n380), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n399), .B1(new_n401), .B2(new_n407), .ZN(new_n857));
  OAI211_X1 g0657(.A(KEYINPUT102), .B(new_n295), .C1(new_n857), .C2(KEYINPUT16), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n422), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n394), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT102), .B1(new_n861), .B2(new_n295), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n856), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n643), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n855), .B1(new_n447), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT104), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n444), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n424), .B1(new_n438), .B2(new_n393), .ZN(new_n870));
  INV_X1    g0670(.A(new_n425), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT103), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT102), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n407), .A2(G68), .A3(new_n420), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT16), .B1(new_n876), .B2(new_n418), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n877), .B2(new_n433), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(new_n422), .A3(new_n858), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n443), .B1(new_n879), .B2(new_n856), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT103), .B1(new_n880), .B2(new_n426), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n874), .A2(new_n881), .A3(new_n865), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n430), .B(new_n439), .C1(new_n444), .C2(new_n864), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n872), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n868), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  AOI211_X1 g0688(.A(KEYINPUT104), .B(new_n886), .C1(new_n882), .C2(KEYINPUT37), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n867), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT105), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT105), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n867), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n447), .A2(new_n866), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n888), .B2(new_n889), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n891), .A2(new_n893), .B1(new_n855), .B2(new_n895), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n802), .A2(new_n815), .B1(new_n369), .B2(new_n645), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n314), .A2(new_n645), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n315), .A2(new_n318), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n290), .A2(new_n314), .A3(new_n645), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n854), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n890), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n622), .B1(new_n427), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n427), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n440), .A2(new_n864), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n621), .A2(new_n412), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n887), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n904), .A2(new_n913), .A3(KEYINPUT39), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n896), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n315), .A2(new_n645), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n903), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n456), .ZN(new_n919));
  INV_X1    g0719(.A(new_n679), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n628), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n918), .B(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n680), .B1(new_n712), .B2(new_n652), .ZN(new_n924));
  OAI211_X1 g0724(.A(KEYINPUT31), .B(new_n645), .C1(new_n699), .C2(new_n710), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n925), .A3(new_n705), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT107), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT107), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n924), .A2(new_n925), .A3(new_n705), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n815), .B1(new_n899), .B2(new_n900), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n923), .B1(new_n896), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n932), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(KEYINPUT40), .C1(new_n904), .C2(new_n913), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n930), .A2(new_n456), .ZN(new_n937));
  OAI21_X1  g0737(.A(G330), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n922), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(KEYINPUT108), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n253), .B1(G13), .B2(new_n227), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n922), .B2(new_n939), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT108), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n944), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n853), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT109), .ZN(G367));
  OAI21_X1  g0748(.A(new_n740), .B1(new_n230), .B2(new_n362), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n241), .A2(new_n729), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n722), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n761), .A2(new_n782), .B1(new_n745), .B2(new_n557), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n323), .B(new_n952), .C1(G303), .C2(new_n785), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n757), .A2(new_n508), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT46), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G107), .A2(new_n750), .B1(new_n954), .B2(KEYINPUT46), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n764), .A2(new_n783), .B1(new_n753), .B2(new_n202), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G317), .B2(new_n773), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n953), .A2(new_n955), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n749), .A2(new_n216), .ZN(new_n960));
  INV_X1    g0760(.A(G137), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n745), .A2(new_n771), .B1(new_n770), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n323), .B1(new_n761), .B2(new_n827), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n785), .A2(G150), .B1(new_n758), .B2(G58), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n753), .A2(new_n208), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G50), .B2(new_n765), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT47), .B1(new_n959), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n795), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n959), .A2(KEYINPUT47), .A3(new_n968), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n951), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n603), .A2(new_n645), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n616), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n675), .A2(new_n973), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT110), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n972), .B1(new_n978), .B2(new_n798), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n672), .A2(new_n645), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n494), .B(new_n499), .C1(new_n497), .C2(new_n652), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n658), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT45), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n658), .A2(new_n982), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n656), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n657), .A2(new_n651), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n655), .B2(new_n657), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n650), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n716), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n716), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n663), .B(KEYINPUT41), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n721), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n988), .A2(new_n982), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT112), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT111), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1000), .B(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n990), .B1(new_n981), .B2(new_n980), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n494), .B1(new_n981), .B2(new_n654), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1005), .A2(KEYINPUT42), .B1(new_n652), .B2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1006), .A2(new_n1008), .B1(KEYINPUT43), .B2(new_n978), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1003), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n979), .B1(new_n998), .B2(new_n1010), .ZN(G387));
  OR2_X1    g0811(.A1(new_n655), .A2(new_n798), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n745), .A2(new_n782), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n767), .A2(new_n1014), .B1(new_n764), .B2(new_n518), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G322), .C2(new_n762), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT48), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(KEYINPUT48), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n749), .A2(new_n783), .B1(new_n757), .B2(new_n557), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1020), .A2(KEYINPUT49), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n271), .B1(new_n770), .B2(new_n788), .C1(new_n508), .C2(new_n753), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(KEYINPUT49), .B2(new_n1020), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n216), .A2(new_n764), .B1(new_n745), .B2(new_n338), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n271), .B(new_n1025), .C1(G97), .C2(new_n754), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n757), .A2(new_n208), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n761), .A2(new_n771), .B1(new_n770), .B2(new_n339), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G50), .C2(new_n785), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1026), .B(new_n1029), .C1(new_n362), .C2(new_n749), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n795), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n238), .A2(G45), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n661), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n338), .A2(G50), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT113), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1036), .B(new_n1037), .C1(new_n661), .C2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1032), .B(new_n729), .C1(new_n1034), .C2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n661), .A2(new_n725), .B1(new_n203), .B2(new_n662), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n741), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1031), .A2(new_n838), .A3(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n992), .A2(new_n721), .B1(new_n1012), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n663), .B(KEYINPUT114), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n993), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n716), .A2(new_n992), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(G393));
  OAI21_X1  g0848(.A(new_n740), .B1(new_n202), .B2(new_n230), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n248), .A2(new_n730), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n722), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G68), .A2(new_n758), .B1(new_n773), .B2(G143), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n323), .C1(new_n210), .C2(new_n753), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT115), .Z(new_n1054));
  OAI22_X1  g0854(.A1(new_n767), .A2(new_n771), .B1(new_n761), .B2(new_n339), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT51), .Z(new_n1056));
  NOR2_X1   g0856(.A1(new_n749), .A2(new_n208), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n830), .A2(new_n745), .B1(new_n764), .B2(new_n338), .ZN(new_n1058));
  OR4_X1    g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G283), .A2(new_n758), .B1(new_n773), .B2(G322), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n271), .A3(new_n755), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT116), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n767), .A2(new_n782), .B1(new_n761), .B2(new_n1014), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n557), .A2(new_n764), .B1(new_n745), .B2(new_n518), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G116), .B2(new_n750), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT117), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1068), .A2(new_n795), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1059), .A2(KEYINPUT117), .A3(new_n1067), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1051), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n798), .B2(new_n982), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n721), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n994), .A2(new_n1045), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n989), .A2(new_n993), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1072), .B1(new_n1073), .B2(new_n989), .C1(new_n1074), .C2(new_n1075), .ZN(G390));
  INV_X1    g0876(.A(new_n917), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n902), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n914), .B(new_n1078), .C1(new_n915), .C2(new_n896), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n678), .A2(new_n841), .B1(new_n370), .B2(new_n652), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n901), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .C1(new_n904), .C2(new_n913), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n901), .A2(new_n841), .A3(G330), .A4(new_n714), .ZN(new_n1083));
  INV_X1    g0883(.A(G330), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n927), .B2(new_n929), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n931), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT118), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1083), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1079), .A2(new_n1082), .A3(new_n1089), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1084), .B(new_n815), .C1(new_n927), .C2(new_n929), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT119), .B1(new_n1091), .B2(new_n901), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n930), .A2(G330), .A3(new_n841), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT119), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n1081), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1092), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n901), .B1(new_n715), .B2(new_n841), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n897), .B1(new_n1087), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1085), .A2(new_n456), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n628), .B(new_n1102), .C1(new_n919), .C2(new_n920), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1090), .B(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1105), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1079), .A2(new_n1082), .A3(new_n1089), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1112), .A3(new_n1045), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n916), .A2(new_n738), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n838), .B1(new_n839), .B2(new_n338), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n785), .A2(G116), .B1(new_n754), .B2(G68), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n271), .A3(new_n759), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1057), .B(new_n1117), .C1(G294), .C2(new_n780), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G283), .A2(new_n762), .B1(new_n765), .B2(G97), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n203), .B2(new_n745), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n271), .B1(new_n762), .B2(G128), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n771), .B2(new_n749), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n745), .A2(new_n961), .B1(new_n753), .B2(new_n830), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n767), .A2(new_n834), .B1(new_n764), .B2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n758), .A2(G150), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G125), .B2(new_n780), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1118), .A2(new_n1121), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1115), .B1(new_n1131), .B2(new_n795), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1114), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1090), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n721), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1113), .A2(new_n1135), .A3(KEYINPUT121), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT121), .B1(new_n1113), .B2(new_n1135), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(G378));
  NAND2_X1  g0938(.A1(new_n891), .A2(new_n893), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n895), .A2(new_n855), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n932), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(G330), .B(new_n935), .C1(new_n1141), .C2(KEYINPUT40), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1143));
  OR3_X1    g0943(.A1(new_n626), .A2(new_n346), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n626), .B2(new_n346), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n345), .A2(new_n864), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1142), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n933), .A2(new_n1148), .A3(G330), .A4(new_n935), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n918), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT123), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1150), .A2(new_n918), .A3(new_n1151), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1101), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1104), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1152), .A2(KEYINPUT123), .A3(new_n1153), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1045), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n1158), .B2(new_n1104), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1157), .A2(new_n721), .A3(new_n1160), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1148), .A2(new_n738), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n764), .A2(new_n362), .B1(new_n753), .B2(new_n214), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n761), .A2(new_n508), .B1(new_n745), .B2(new_n202), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n780), .C2(G283), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n271), .A2(new_n260), .A3(new_n262), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n960), .A2(new_n1027), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n785), .A2(G107), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT122), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1173), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT58), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1174), .B(new_n830), .C1(G33), .C2(G41), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n765), .A2(G137), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n757), .B2(new_n1125), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n785), .A2(G128), .B1(new_n762), .B2(G125), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n834), .B2(new_n745), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G150), .C2(new_n750), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n754), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n773), .C2(G124), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1182), .B1(new_n1179), .B2(new_n1178), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n736), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n838), .B1(new_n839), .B2(new_n830), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1170), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1169), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1168), .A2(new_n1201), .ZN(G375));
  NAND3_X1  g1002(.A1(new_n1098), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1105), .A2(new_n997), .A3(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT124), .Z(new_n1205));
  AOI21_X1  g1005(.A(new_n838), .B1(new_n839), .B2(new_n216), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n761), .A2(new_n557), .B1(new_n745), .B2(new_n508), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n749), .A2(new_n362), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n323), .A4(new_n966), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n785), .A2(G283), .B1(new_n758), .B2(G97), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n203), .B2(new_n764), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G303), .B2(new_n780), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n785), .A2(G137), .B1(new_n758), .B2(G159), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n339), .B2(new_n764), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G128), .B2(new_n780), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n323), .B1(new_n753), .B2(new_n214), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n761), .A2(new_n834), .B1(new_n745), .B2(new_n1125), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G50), .C2(new_n750), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1209), .A2(new_n1212), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1206), .B1(new_n795), .B2(new_n1219), .C1(new_n901), .C2(new_n738), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1093), .A2(new_n1081), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1096), .B1(new_n1221), .B2(KEYINPUT119), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1099), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1086), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1222), .A2(new_n1095), .B1(new_n1224), .B2(new_n897), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1220), .B1(new_n1225), .B2(new_n1073), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1205), .A2(new_n1227), .ZN(G381));
  NAND2_X1  g1028(.A1(new_n1113), .A2(new_n1135), .ZN(new_n1229));
  OR2_X1    g1029(.A1(G387), .A2(G390), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G396), .A2(new_n1230), .A3(G384), .A4(G393), .ZN(new_n1231));
  OR4_X1    g1031(.A1(new_n1229), .A2(new_n1231), .A3(G375), .A4(G381), .ZN(G407));
  AOI21_X1  g1032(.A(new_n1200), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1229), .ZN(new_n1234));
  INV_X1    g1034(.A(G213), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(G343), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(G407), .A2(G213), .A3(new_n1237), .ZN(G409));
  NAND2_X1  g1038(.A1(new_n1236), .A2(G2897), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1098), .A2(KEYINPUT60), .A3(new_n1100), .A4(new_n1103), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT125), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1164), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1203), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT126), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1225), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1103), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1240), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT126), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1244), .A4(new_n1242), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1246), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1227), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n843), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(G384), .A3(new_n1227), .ZN(new_n1256));
  AOI211_X1 g1056(.A(KEYINPUT127), .B(new_n1239), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1255), .A2(KEYINPUT127), .A3(new_n1256), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1239), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1257), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1168), .A2(G378), .A3(new_n1201), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1157), .A2(new_n997), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1198), .B1(new_n1166), .B2(new_n721), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1229), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1236), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1272), .B2(new_n1258), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G387), .B(G390), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(G393), .B(new_n800), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1276), .B(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1236), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G384), .B1(new_n1253), .B2(new_n1227), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n843), .B(new_n1226), .C1(new_n1246), .C2(new_n1252), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1273), .A2(new_n1275), .A3(new_n1279), .A4(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1258), .A2(new_n1259), .A3(new_n1262), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1239), .B1(new_n1283), .B2(KEYINPUT127), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1283), .A2(KEYINPUT127), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1286), .B1(new_n1290), .B2(new_n1280), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1268), .B1(new_n1233), .B2(G378), .ZN(new_n1292));
  NOR4_X1   g1092(.A1(new_n1292), .A2(KEYINPUT62), .A3(new_n1236), .A4(new_n1258), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1291), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1285), .B1(new_n1296), .B2(new_n1279), .ZN(G405));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1234), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1265), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1279), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1278), .A2(new_n1265), .A3(new_n1298), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1258), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1283), .A3(new_n1301), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(G402));
endmodule


