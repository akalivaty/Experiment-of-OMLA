

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584;

  AND2_X1 U324 ( .A1(n560), .A2(n549), .ZN(n399) );
  XNOR2_X1 U325 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n402) );
  XNOR2_X1 U326 ( .A(n403), .B(n402), .ZN(n409) );
  XNOR2_X1 U327 ( .A(n443), .B(KEYINPUT121), .ZN(n444) );
  XNOR2_X1 U328 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U329 ( .A(n572), .B(KEYINPUT41), .Z(n549) );
  XNOR2_X1 U330 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U331 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n293) );
  XNOR2_X1 U333 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n305) );
  XOR2_X1 U335 ( .A(G134GAT), .B(G190GAT), .Z(n295) );
  XOR2_X1 U336 ( .A(G120GAT), .B(G71GAT), .Z(n396) );
  XOR2_X1 U337 ( .A(G15GAT), .B(G127GAT), .Z(n358) );
  XNOR2_X1 U338 ( .A(n396), .B(n358), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U340 ( .A(n296), .B(G99GAT), .Z(n303) );
  XOR2_X1 U341 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n298) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n311) );
  XOR2_X1 U344 ( .A(n311), .B(KEYINPUT83), .Z(n300) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U350 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n307) );
  XNOR2_X1 U351 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U353 ( .A(G169GAT), .B(n308), .Z(n416) );
  XOR2_X1 U354 ( .A(n309), .B(n416), .Z(n509) );
  XNOR2_X1 U355 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n310), .B(KEYINPUT2), .ZN(n430) );
  XNOR2_X1 U357 ( .A(n311), .B(n430), .ZN(n330) );
  XOR2_X1 U358 ( .A(KEYINPUT4), .B(G148GAT), .Z(n313) );
  XNOR2_X1 U359 ( .A(G120GAT), .B(G127GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U361 ( .A(G57GAT), .B(KEYINPUT90), .Z(n315) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(KEYINPUT91), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U364 ( .A(n317), .B(n316), .Z(n328) );
  XOR2_X1 U365 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n319) );
  XNOR2_X1 U366 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n326) );
  XOR2_X1 U368 ( .A(G134GAT), .B(KEYINPUT75), .Z(n333) );
  XOR2_X1 U369 ( .A(G85GAT), .B(G162GAT), .Z(n321) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(G141GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U372 ( .A(n333), .B(n322), .Z(n324) );
  NAND2_X1 U373 ( .A1(G225GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U376 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U377 ( .A(n330), .B(n329), .Z(n502) );
  INV_X1 U378 ( .A(n502), .ZN(n518) );
  XOR2_X1 U379 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n332) );
  XNOR2_X1 U380 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n344) );
  XOR2_X1 U382 ( .A(KEYINPUT74), .B(KEYINPUT64), .Z(n335) );
  XOR2_X1 U383 ( .A(G50GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U384 ( .A(n437), .B(n333), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .Z(n411) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n336), .B(KEYINPUT71), .ZN(n388) );
  XOR2_X1 U389 ( .A(n411), .B(n388), .Z(n338) );
  NAND2_X1 U390 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n342) );
  XOR2_X1 U393 ( .A(G218GAT), .B(G106GAT), .Z(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U396 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n346) );
  XNOR2_X1 U397 ( .A(G43GAT), .B(G29GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U399 ( .A(KEYINPUT69), .B(n347), .ZN(n379) );
  XNOR2_X1 U400 ( .A(n348), .B(n379), .ZN(n404) );
  XOR2_X1 U401 ( .A(G64GAT), .B(KEYINPUT79), .Z(n350) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U404 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n352) );
  XNOR2_X1 U405 ( .A(KEYINPUT76), .B(KEYINPUT78), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U407 ( .A(n354), .B(n353), .Z(n360) );
  XOR2_X1 U408 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n356) );
  XNOR2_X1 U409 ( .A(G183GAT), .B(G71GAT), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U413 ( .A(G57GAT), .B(KEYINPUT13), .Z(n391) );
  XOR2_X1 U414 ( .A(n391), .B(G78GAT), .Z(n362) );
  XOR2_X1 U415 ( .A(G1GAT), .B(G8GAT), .Z(n372) );
  XNOR2_X1 U416 ( .A(n372), .B(G211GAT), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U418 ( .A(n364), .B(n363), .Z(n366) );
  XNOR2_X1 U419 ( .A(G22GAT), .B(G155GAT), .ZN(n365) );
  XOR2_X1 U420 ( .A(n366), .B(n365), .Z(n454) );
  INV_X1 U421 ( .A(n454), .ZN(n576) );
  XOR2_X1 U422 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n368) );
  XNOR2_X1 U423 ( .A(KEYINPUT70), .B(KEYINPUT68), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n383) );
  XOR2_X1 U425 ( .A(G113GAT), .B(G197GAT), .Z(n370) );
  XNOR2_X1 U426 ( .A(G36GAT), .B(G50GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U428 ( .A(n371), .B(G15GAT), .Z(n374) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(n372), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U431 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n376) );
  NAND2_X1 U432 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U434 ( .A(n378), .B(n377), .Z(n381) );
  XOR2_X1 U435 ( .A(G141GAT), .B(G22GAT), .Z(n438) );
  XOR2_X1 U436 ( .A(n379), .B(n438), .Z(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n560) );
  XOR2_X1 U439 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n385) );
  NAND2_X1 U440 ( .A1(G230GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U442 ( .A(n386), .B(KEYINPUT31), .Z(n390) );
  XNOR2_X1 U443 ( .A(G106GAT), .B(G78GAT), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n387), .B(G148GAT), .ZN(n429) );
  XNOR2_X1 U445 ( .A(n429), .B(n388), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n392) );
  XOR2_X1 U447 ( .A(n392), .B(n391), .Z(n398) );
  XOR2_X1 U448 ( .A(G92GAT), .B(KEYINPUT72), .Z(n394) );
  XNOR2_X1 U449 ( .A(G204GAT), .B(G64GAT), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U451 ( .A(G176GAT), .B(n395), .Z(n414) );
  XNOR2_X1 U452 ( .A(n396), .B(n414), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n572) );
  XNOR2_X1 U454 ( .A(n399), .B(KEYINPUT46), .ZN(n400) );
  NOR2_X1 U455 ( .A1(n576), .A2(n400), .ZN(n401) );
  NAND2_X1 U456 ( .A1(n404), .A2(n401), .ZN(n403) );
  INV_X1 U457 ( .A(n404), .ZN(n557) );
  XOR2_X1 U458 ( .A(KEYINPUT36), .B(n557), .Z(n581) );
  NOR2_X1 U459 ( .A1(n581), .A2(n454), .ZN(n405) );
  XNOR2_X1 U460 ( .A(KEYINPUT45), .B(n405), .ZN(n406) );
  INV_X1 U461 ( .A(n560), .ZN(n567) );
  NAND2_X1 U462 ( .A1(n406), .A2(n567), .ZN(n407) );
  NOR2_X1 U463 ( .A1(n407), .A2(n572), .ZN(n408) );
  NOR2_X1 U464 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n410), .B(KEYINPUT48), .ZN(n529) );
  XOR2_X1 U466 ( .A(n411), .B(G8GAT), .Z(n413) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U469 ( .A(n415), .B(n414), .Z(n422) );
  INV_X1 U470 ( .A(n416), .ZN(n420) );
  XOR2_X1 U471 ( .A(KEYINPUT21), .B(G218GAT), .Z(n418) );
  XNOR2_X1 U472 ( .A(KEYINPUT85), .B(G211GAT), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U474 ( .A(G197GAT), .B(n419), .Z(n441) );
  XOR2_X1 U475 ( .A(n420), .B(n441), .Z(n421) );
  XOR2_X1 U476 ( .A(n422), .B(n421), .Z(n506) );
  XNOR2_X1 U477 ( .A(KEYINPUT120), .B(n506), .ZN(n423) );
  NOR2_X1 U478 ( .A1(n529), .A2(n423), .ZN(n424) );
  XOR2_X1 U479 ( .A(KEYINPUT54), .B(n424), .Z(n425) );
  NOR2_X1 U480 ( .A1(n518), .A2(n425), .ZN(n566) );
  XOR2_X1 U481 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n427) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n428), .B(KEYINPUT87), .Z(n432) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U487 ( .A(G204GAT), .B(KEYINPUT22), .Z(n434) );
  XNOR2_X1 U488 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U493 ( .A(n442), .B(n441), .Z(n463) );
  AND2_X1 U494 ( .A1(n566), .A2(n463), .ZN(n445) );
  INV_X1 U495 ( .A(KEYINPUT55), .ZN(n443) );
  NOR2_X1 U496 ( .A1(n509), .A2(n446), .ZN(n562) );
  NAND2_X1 U497 ( .A1(n562), .A2(n549), .ZN(n449) );
  XOR2_X1 U498 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n447) );
  XNOR2_X1 U499 ( .A(n447), .B(G176GAT), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  NAND2_X1 U501 ( .A1(n562), .A2(n557), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n450) );
  NOR2_X1 U503 ( .A1(n572), .A2(n567), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT73), .ZN(n487) );
  NOR2_X1 U505 ( .A1(n557), .A2(n454), .ZN(n455) );
  XNOR2_X1 U506 ( .A(n455), .B(KEYINPUT16), .ZN(n469) );
  INV_X1 U507 ( .A(n509), .ZN(n530) );
  INV_X1 U508 ( .A(n506), .ZN(n521) );
  NAND2_X1 U509 ( .A1(n530), .A2(n521), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n463), .A2(n456), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT25), .B(n457), .Z(n461) );
  XNOR2_X1 U512 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n530), .A2(n463), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n565) );
  XOR2_X1 U515 ( .A(n506), .B(KEYINPUT27), .Z(n465) );
  NAND2_X1 U516 ( .A1(n565), .A2(n465), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U518 ( .A1(n462), .A2(n502), .ZN(n468) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT65), .ZN(n464) );
  XOR2_X1 U520 ( .A(n464), .B(KEYINPUT28), .Z(n512) );
  INV_X1 U521 ( .A(n512), .ZN(n533) );
  NAND2_X1 U522 ( .A1(n518), .A2(n465), .ZN(n528) );
  NOR2_X1 U523 ( .A1(n533), .A2(n528), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n466), .A2(n509), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n484) );
  NAND2_X1 U526 ( .A1(n469), .A2(n484), .ZN(n500) );
  NOR2_X1 U527 ( .A1(n487), .A2(n500), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT93), .B(n470), .Z(n480) );
  NAND2_X1 U529 ( .A1(n480), .A2(n518), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n472) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n480), .A2(n521), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(KEYINPUT96), .ZN(n476) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n476), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U538 ( .A1(n480), .A2(n530), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U540 ( .A(G15GAT), .B(n479), .Z(G1326GAT) );
  NAND2_X1 U541 ( .A1(n480), .A2(n533), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT98), .ZN(n482) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n491) );
  NOR2_X1 U545 ( .A1(n581), .A2(n576), .ZN(n483) );
  NAND2_X1 U546 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n485), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT100), .B(n486), .Z(n517) );
  NOR2_X1 U549 ( .A1(n517), .A2(n487), .ZN(n489) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(KEYINPUT101), .Z(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(n498) );
  NAND2_X1 U552 ( .A1(n518), .A2(n498), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U554 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NAND2_X1 U555 ( .A1(n498), .A2(n521), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n493), .B(KEYINPUT102), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n496) );
  NAND2_X1 U559 ( .A1(n530), .A2(n498), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n498), .A2(n533), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U564 ( .A1(n567), .A2(n549), .ZN(n516) );
  NOR2_X1 U565 ( .A1(n500), .A2(n516), .ZN(n501) );
  XOR2_X1 U566 ( .A(KEYINPUT104), .B(n501), .Z(n513) );
  NOR2_X1 U567 ( .A1(n513), .A2(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n513), .A2(n506), .ZN(n507) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(n507), .Z(n508) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n513), .A2(n509), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n518), .A2(n524), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n524), .A2(n521), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n530), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U589 ( .A1(n524), .A2(n533), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n545) );
  NAND2_X1 U593 ( .A1(n530), .A2(n545), .ZN(n531) );
  XOR2_X1 U594 ( .A(KEYINPUT111), .B(n531), .Z(n532) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n560), .A2(n541), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U599 ( .A1(n541), .A2(n549), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(KEYINPUT112), .ZN(n540) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n538) );
  NAND2_X1 U603 ( .A1(n541), .A2(n576), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n543) );
  NAND2_X1 U607 ( .A1(n541), .A2(n557), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n565), .A2(n545), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT115), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n558), .A2(n560), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n551) );
  NAND2_X1 U616 ( .A1(n558), .A2(n549), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT53), .Z(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U621 ( .A1(n558), .A2(n576), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n562), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(n561), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n576), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT122), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G183GAT), .B(n564), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n580) );
  NOR2_X1 U633 ( .A1(n567), .A2(n580), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U638 ( .A(n580), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n577), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

