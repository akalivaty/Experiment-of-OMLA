//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT16), .ZN(new_n200));
  OR3_X1    g014(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G128), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G110), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n211), .A2(KEYINPUT73), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT24), .B(G110), .Z(new_n213));
  XNOR2_X1  g027(.A(G119), .B(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(new_n211), .B2(KEYINPUT73), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n203), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(G110), .A2(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n218));
  INV_X1    g032(.A(new_n202), .ZN(new_n219));
  AOI21_X1  g033(.A(G146), .B1(new_n200), .B2(new_n201), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n191), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n217), .A2(new_n222), .A3(new_n191), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(G234), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G902), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT76), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n224), .A2(new_n225), .A3(G902), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT74), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(KEYINPUT75), .B2(KEYINPUT25), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n229), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n217), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n221), .A3(new_n190), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n238), .A2(new_n223), .A3(KEYINPUT74), .A4(new_n228), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n239), .B2(KEYINPUT75), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n232), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n244), .B(G146), .C1(new_n208), .C2(KEYINPUT1), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n208), .A2(new_n198), .A3(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n198), .A2(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n244), .A2(G146), .ZN(new_n254));
  AND4_X1   g068(.A1(new_n249), .A2(new_n251), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n248), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n257), .A2(G137), .ZN(new_n260));
  OAI21_X1  g074(.A(G131), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n257), .B2(G137), .ZN(new_n263));
  INV_X1    g077(.A(G137), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT11), .A3(G134), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .A4(new_n258), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n253), .A2(new_n254), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT64), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n250), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n253), .A2(new_n254), .ZN(new_n275));
  OR2_X1    g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n272), .A2(new_n274), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n263), .A2(new_n258), .A3(new_n265), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G131), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n267), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n256), .A2(new_n269), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n205), .A2(G116), .ZN(new_n284));
  INV_X1    g098(.A(G116), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G119), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT2), .B(G113), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n281), .A2(new_n267), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n275), .A2(new_n277), .A3(new_n276), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n273), .B1(new_n250), .B2(new_n270), .ZN(new_n294));
  AND4_X1   g108(.A1(new_n273), .A2(new_n253), .A3(new_n254), .A4(new_n270), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n250), .A2(new_n249), .A3(new_n251), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n247), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI22_X1  g114(.A1(new_n292), .A2(new_n296), .B1(new_n300), .B2(new_n268), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n289), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n243), .B1(new_n291), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT71), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n289), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT28), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT26), .B(G101), .Z(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G210), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n304), .A2(new_n309), .A3(new_n310), .A4(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n308), .ZN(new_n321));
  INV_X1    g135(.A(new_n303), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n317), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n289), .B1(new_n301), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n283), .B2(KEYINPUT30), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n301), .A2(KEYINPUT66), .A3(new_n324), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n301), .A2(new_n289), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n329), .A2(new_n330), .A3(new_n316), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n318), .B1(new_n323), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n320), .A2(new_n332), .A3(new_n228), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G472), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n291), .A2(new_n316), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT31), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n290), .B1(new_n283), .B2(KEYINPUT30), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n283), .A2(new_n326), .A3(KEYINPUT30), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT66), .B1(new_n301), .B2(new_n324), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT31), .ZN(new_n341));
  INV_X1    g155(.A(new_n335), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n317), .B1(new_n308), .B2(new_n303), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n336), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT69), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n336), .A2(new_n343), .A3(new_n344), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G472), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n228), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n334), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n356));
  AOI21_X1  g170(.A(G902), .B1(new_n346), .B2(new_n348), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n350), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n242), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n312), .A2(G214), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n244), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n312), .A2(G143), .A3(G214), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G131), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT17), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n266), .A3(new_n362), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT92), .B1(new_n219), .B2(new_n220), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n363), .A2(KEYINPUT17), .A3(G131), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n200), .A2(new_n201), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n198), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n202), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G113), .B(G122), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT89), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n196), .B2(G146), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n196), .A2(G146), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n196), .A2(new_n378), .A3(G146), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT18), .A2(G131), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT90), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n361), .A3(new_n362), .ZN(new_n386));
  INV_X1    g200(.A(new_n384), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n363), .A2(KEYINPUT88), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT88), .B1(new_n363), .B2(new_n387), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n383), .B(new_n386), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n374), .A2(new_n377), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n377), .B1(new_n374), .B2(new_n390), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n228), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(KEYINPUT93), .ZN(new_n394));
  INV_X1    g208(.A(G475), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n393), .B2(KEYINPUT93), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(G475), .A2(G902), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n219), .B1(new_n364), .B2(new_n366), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n197), .A2(KEYINPUT91), .A3(KEYINPUT19), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT19), .B1(new_n197), .B2(KEYINPUT91), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n399), .B1(new_n402), .B2(G146), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n377), .B1(new_n403), .B2(new_n390), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n398), .B1(new_n391), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT20), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n390), .ZN(new_n407));
  INV_X1    g221(.A(new_n377), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n374), .A2(new_n377), .A3(new_n390), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n398), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n397), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G478), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(KEYINPUT15), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G122), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT94), .B1(new_n419), .B2(G116), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT94), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n285), .A3(G122), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G107), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(G116), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT95), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n244), .B2(G128), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n208), .A2(KEYINPUT95), .A3(G143), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n428), .A2(new_n429), .B1(G128), .B2(new_n244), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n430), .A2(new_n257), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n257), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n423), .A2(KEYINPUT14), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n423), .A2(KEYINPUT14), .B1(G116), .B2(new_n419), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n424), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT13), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n430), .B1(new_n437), .B2(new_n257), .ZN(new_n438));
  INV_X1    g252(.A(new_n426), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT13), .B1(new_n428), .B2(new_n429), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n430), .A2(new_n442), .A3(new_n257), .ZN(new_n443));
  OAI22_X1  g257(.A1(new_n433), .A2(new_n436), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT9), .B(G234), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n445), .A2(new_n227), .A3(G953), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  OAI221_X1 g262(.A(new_n446), .B1(new_n441), .B2(new_n443), .C1(new_n436), .C2(new_n433), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n418), .B1(new_n450), .B2(new_n228), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI211_X1 g266(.A(G902), .B(new_n417), .C1(new_n448), .C2(new_n449), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT96), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT96), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n451), .B2(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(G234), .A2(G237), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(G952), .A3(new_n188), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT97), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(G898), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n459), .A2(G902), .A3(G953), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n415), .A2(new_n458), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G221), .B1(new_n445), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G469), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n188), .A2(G227), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT77), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G140), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT3), .B1(new_n376), .B2(G107), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n424), .A3(G104), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n376), .A2(G107), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G101), .ZN(new_n480));
  INV_X1    g294(.A(G101), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n475), .A2(new_n477), .A3(new_n481), .A4(new_n478), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(KEYINPUT4), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT4), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(new_n484), .A3(G101), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n279), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT78), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n279), .A2(new_n483), .A3(KEYINPUT78), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n376), .A2(G107), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n424), .A2(G104), .ZN(new_n492));
  OAI21_X1  g306(.A(G101), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT10), .B1(new_n300), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT10), .ZN(new_n496));
  INV_X1    g310(.A(new_n494), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n256), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n490), .A2(new_n292), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n292), .B1(new_n490), .B2(new_n499), .ZN(new_n501));
  OAI211_X1 g315(.A(KEYINPUT79), .B(new_n474), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n488), .A2(new_n489), .B1(new_n495), .B2(new_n498), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n474), .B1(new_n503), .B2(new_n292), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n256), .A2(new_n497), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n300), .A2(new_n494), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n282), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n490), .A2(new_n499), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n282), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n292), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT79), .B1(new_n515), .B2(new_n474), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n469), .B(new_n228), .C1(new_n511), .C2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n469), .A2(new_n228), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n509), .A2(new_n514), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n519), .A2(new_n474), .B1(new_n513), .B2(new_n504), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n520), .B2(G469), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n468), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n483), .A2(new_n289), .A3(new_n485), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n287), .A2(new_n288), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT80), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n284), .B2(KEYINPUT5), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT5), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n528), .A2(new_n205), .A3(KEYINPUT80), .A4(G116), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n526), .A2(new_n527), .A3(G113), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n497), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G122), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n523), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT6), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n523), .A2(new_n531), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n532), .B(KEYINPUT81), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT6), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(new_n537), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n245), .A2(new_n194), .A3(new_n246), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n252), .B2(new_n255), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n296), .A2(G125), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT82), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n545), .B(new_n541), .C1(new_n252), .C2(new_n255), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G224), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G953), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n549), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n543), .A2(new_n544), .A3(new_n546), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n540), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G210), .B1(G237), .B2(G902), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n555), .B(KEYINPUT86), .Z(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n532), .B(KEYINPUT8), .Z(new_n558));
  NAND2_X1  g372(.A1(new_n530), .A2(new_n524), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n494), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n531), .B2(new_n560), .ZN(new_n561));
  AND4_X1   g375(.A1(new_n543), .A2(new_n544), .A3(new_n546), .A4(new_n551), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(KEYINPUT7), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT83), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n549), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n564), .B2(new_n565), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT84), .B1(new_n547), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n547), .A2(KEYINPUT84), .A3(new_n567), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n563), .B(KEYINPUT85), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n533), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n547), .A2(new_n567), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT84), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n547), .A2(KEYINPUT84), .A3(new_n567), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT85), .B1(new_n576), .B2(new_n563), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n554), .B(new_n557), .C1(new_n571), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT87), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n554), .B1(new_n571), .B2(new_n577), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n556), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT85), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n569), .A2(new_n568), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n531), .A2(new_n560), .ZN(new_n584));
  OAI22_X1  g398(.A1(new_n584), .A2(new_n558), .B1(new_n552), .B2(new_n565), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n533), .A3(new_n570), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT87), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n554), .A4(new_n557), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n579), .A2(new_n581), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G214), .B1(G237), .B2(G902), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n466), .A2(new_n522), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n359), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n481), .ZN(G3));
  AOI211_X1 g408(.A(new_n241), .B(new_n468), .C1(new_n517), .C2(new_n521), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n349), .A2(new_n350), .A3(new_n228), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n349), .A2(new_n228), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n595), .A2(KEYINPUT98), .A3(new_n596), .A4(new_n598), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n581), .A2(new_n578), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n591), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n450), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n606), .A2(new_n607), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n448), .B(new_n449), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n608), .A2(G478), .A3(new_n228), .A4(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n450), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n416), .B1(new_n613), .B2(G902), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n415), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n605), .A2(new_n465), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n603), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT100), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT34), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n414), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n406), .A2(new_n413), .A3(KEYINPUT101), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n465), .B(KEYINPUT102), .Z(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(new_n458), .A3(new_n397), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT103), .ZN(new_n628));
  INV_X1    g442(.A(new_n591), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n581), .B2(new_n578), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n623), .A2(new_n624), .B1(new_n394), .B2(new_n396), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n458), .A4(new_n626), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n628), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n603), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT104), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n236), .A2(new_n240), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n237), .A2(new_n221), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n639), .B1(new_n231), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n598), .A2(new_n644), .A3(new_n596), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n592), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT37), .B(G110), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  INV_X1    g462(.A(new_n356), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n596), .A2(new_n649), .ZN(new_n650));
  AOI22_X1  g464(.A1(G472), .A2(new_n333), .B1(new_n349), .B2(new_n353), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(KEYINPUT105), .A2(G900), .ZN(new_n653));
  NAND2_X1  g467(.A1(KEYINPUT105), .A2(G900), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n464), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n461), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n625), .A2(new_n458), .A3(new_n397), .A4(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n517), .A2(new_n521), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n467), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n605), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n652), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(new_n656), .B(KEYINPUT39), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n522), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT40), .Z(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n590), .B(KEYINPUT38), .Z(new_n669));
  AOI21_X1  g483(.A(new_n317), .B1(new_n340), .B2(new_n291), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n291), .A2(new_n302), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n228), .B1(new_n671), .B2(new_n316), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n650), .A2(new_n354), .A3(new_n673), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n394), .A2(new_n396), .B1(new_n406), .B2(new_n413), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n455), .B2(new_n457), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n591), .A3(new_n643), .A4(new_n676), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n667), .A2(new_n668), .A3(new_n669), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n244), .ZN(G45));
  NAND3_X1  g493(.A1(new_n415), .A2(new_n615), .A3(new_n656), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n652), .A2(new_n661), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  AOI21_X1  g497(.A(new_n241), .B1(new_n650), .B2(new_n651), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n474), .B1(new_n500), .B2(new_n501), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT79), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n510), .A3(new_n502), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n469), .B1(new_n688), .B2(new_n228), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n517), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n468), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n684), .A2(new_n617), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT41), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G113), .ZN(G15));
  NAND3_X1  g509(.A1(new_n634), .A2(new_n684), .A3(new_n692), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  OAI21_X1  g511(.A(new_n644), .B1(new_n355), .B2(new_n358), .ZN(new_n698));
  INV_X1    g512(.A(new_n517), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n689), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n466), .A3(new_n467), .A4(new_n630), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n205), .ZN(G21));
  NAND4_X1  g517(.A1(new_n690), .A2(new_n467), .A3(new_n517), .A4(new_n626), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n630), .A2(new_n676), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n304), .A2(new_n309), .A3(new_n310), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n317), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n336), .A2(new_n343), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n351), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n350), .B1(new_n349), .B2(new_n228), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT107), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n713), .B1(new_n357), .B2(new_n350), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n710), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n706), .A2(new_n715), .A3(new_n242), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  NOR3_X1   g531(.A1(new_n691), .A2(new_n605), .A3(new_n468), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n715), .A3(new_n644), .A4(new_n681), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  AND2_X1   g534(.A1(new_n579), .A2(new_n589), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n629), .B1(new_n580), .B2(new_n556), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n681), .A3(new_n522), .A4(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT108), .B1(new_n359), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n579), .A2(new_n581), .A3(new_n591), .A4(new_n589), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n660), .A2(new_n725), .A3(new_n680), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n684), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n724), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n596), .A2(new_n352), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n241), .B1(new_n731), .B2(new_n651), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n726), .A3(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT109), .B(G131), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G33));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n657), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n660), .A2(new_n725), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n684), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  NAND2_X1  g555(.A1(new_n520), .A2(KEYINPUT45), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT111), .ZN(new_n743));
  OAI21_X1  g557(.A(G469), .B1(new_n520), .B2(KEYINPUT45), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n518), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n699), .B1(new_n746), .B2(KEYINPUT46), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(KEYINPUT112), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n746), .A2(KEYINPUT46), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n748), .B2(KEYINPUT112), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n467), .A3(new_n664), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT113), .B1(new_n675), .B2(new_n615), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT43), .Z(new_n755));
  INV_X1    g569(.A(new_n596), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n755), .B(new_n644), .C1(new_n756), .C2(new_n711), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n725), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n264), .ZN(G39));
  INV_X1    g576(.A(new_n725), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n241), .A3(new_n681), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n358), .A3(new_n355), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n467), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT47), .B1(new_n752), .B2(new_n467), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  NAND4_X1  g583(.A1(new_n755), .A2(new_n462), .A3(new_n692), .A4(new_n763), .ZN(new_n770));
  INV_X1    g584(.A(new_n732), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT48), .Z(new_n773));
  AND4_X1   g587(.A1(new_n242), .A2(new_n715), .A3(new_n755), .A4(new_n462), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n718), .ZN(new_n775));
  INV_X1    g589(.A(G952), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n692), .A2(new_n763), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n777), .A2(new_n674), .A3(new_n241), .A4(new_n461), .ZN(new_n778));
  INV_X1    g592(.A(new_n616), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n776), .B(G953), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n773), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n766), .ZN(new_n782));
  INV_X1    g596(.A(new_n767), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n700), .A2(KEYINPUT117), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n700), .A2(KEYINPUT117), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n468), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n763), .A3(new_n774), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n715), .A2(new_n644), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n770), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n774), .A2(new_n629), .A3(new_n669), .A4(new_n692), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT50), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n415), .A2(new_n615), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n790), .B(new_n792), .C1(new_n778), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n781), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n643), .A2(new_n656), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n674), .A2(new_n661), .A3(new_n676), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n719), .A2(new_n662), .A3(new_n800), .A4(new_n682), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT52), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n715), .A2(new_n644), .A3(new_n681), .A4(new_n739), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n625), .A2(new_n397), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n451), .A2(new_n453), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n451), .B2(new_n453), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n656), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n763), .A2(KEYINPUT115), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n631), .A2(new_n656), .A3(new_n807), .A4(new_n808), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n813), .B2(new_n725), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n652), .A2(new_n811), .A3(new_n814), .A4(new_n522), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n803), .A2(new_n815), .A3(new_n740), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n734), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n592), .B1(new_n359), .B2(new_n645), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n702), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n684), .B(new_n692), .C1(new_n634), .C2(new_n617), .ZN(new_n820));
  INV_X1    g634(.A(new_n808), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n675), .B1(new_n821), .B2(new_n806), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n616), .A2(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n591), .A2(new_n823), .A3(new_n590), .A4(new_n626), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n601), .A2(new_n602), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n819), .A2(new_n716), .A3(new_n820), .A4(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT116), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n702), .ZN(new_n828));
  INV_X1    g642(.A(new_n592), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n756), .A2(new_n711), .A3(new_n643), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n829), .B1(new_n684), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n825), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n696), .A2(new_n716), .A3(new_n693), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n734), .A4(new_n816), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n802), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n719), .A2(new_n662), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n838), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n837), .A2(KEYINPUT53), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n817), .A2(new_n826), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n801), .B(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n846), .A2(new_n848), .A3(KEYINPUT53), .A4(new_n841), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n845), .B(new_n849), .C1(new_n837), .C2(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n788), .A2(KEYINPUT51), .A3(new_n794), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n797), .A2(new_n844), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(G952), .B2(G953), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n675), .A2(new_n615), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n242), .A2(new_n591), .A3(new_n467), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n674), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n700), .B(KEYINPUT49), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n669), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n859), .ZN(G75));
  OAI21_X1  g674(.A(new_n849), .B1(new_n837), .B2(KEYINPUT53), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n228), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n556), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n540), .B(KEYINPUT118), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT55), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(new_n553), .Z(new_n868));
  AND3_X1   g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n776), .A2(G953), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT119), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(G51));
  NAND2_X1  g688(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n850), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n861), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n518), .B(KEYINPUT57), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n688), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n861), .A2(G902), .A3(new_n745), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(KEYINPUT121), .A3(new_n872), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n880), .B2(new_n688), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n887), .B2(new_n873), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(G54));
  NAND2_X1  g703(.A1(KEYINPUT58), .A2(G475), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT122), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n863), .A2(new_n411), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n411), .B1(new_n863), .B2(new_n891), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n873), .ZN(G60));
  NAND2_X1  g708(.A1(G478), .A2(G902), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT59), .Z(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n844), .B2(new_n850), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n608), .A2(new_n611), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n872), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n877), .A2(new_n878), .ZN(new_n900));
  INV_X1    g714(.A(new_n896), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(G63));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n861), .A2(new_n642), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n862), .A2(new_n905), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n872), .B(new_n907), .C1(new_n908), .C2(new_n226), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT123), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g725(.A(G953), .B1(new_n463), .B2(new_n548), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n834), .B2(G953), .ZN(new_n913));
  INV_X1    g727(.A(new_n866), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(G898), .B2(new_n188), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n913), .B(new_n915), .ZN(G69));
  NAND3_X1  g730(.A1(new_n719), .A2(new_n662), .A3(new_n682), .ZN(new_n917));
  INV_X1    g731(.A(new_n753), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n760), .B1(new_n705), .B2(new_n771), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n734), .A2(new_n740), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n768), .A3(new_n188), .A4(new_n921), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n327), .A2(new_n328), .B1(KEYINPUT30), .B2(new_n283), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n402), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(G900), .B2(G953), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n665), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n684), .A2(new_n930), .A3(new_n763), .A4(new_n823), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n753), .B2(new_n760), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n678), .A2(new_n917), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT62), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n938), .A3(KEYINPUT62), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n935), .A2(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n782), .A2(new_n783), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n765), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n934), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n188), .ZN(new_n945));
  AOI221_X4 g759(.A(new_n927), .B1(KEYINPUT126), .B2(new_n929), .C1(new_n945), .C2(new_n924), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n929), .B1(new_n927), .B2(KEYINPUT126), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n924), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n926), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n946), .A2(new_n949), .ZN(G72));
  INV_X1    g764(.A(new_n670), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n934), .A2(new_n940), .A3(new_n943), .A4(new_n834), .ZN(new_n952));
  NAND2_X1  g766(.A1(G472), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT63), .Z(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n920), .A2(new_n768), .A3(new_n921), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(new_n826), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n331), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n842), .A2(new_n843), .ZN(new_n959));
  INV_X1    g773(.A(new_n331), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n951), .A3(new_n954), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT127), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NOR4_X1   g777(.A1(new_n955), .A2(new_n958), .A3(new_n873), .A4(new_n963), .ZN(G57));
endmodule


