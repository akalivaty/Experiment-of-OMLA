//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997;
  XNOR2_X1  g000(.A(KEYINPUT69), .B(G71gat), .ZN(new_n202));
  INV_X1    g001(.A(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G15gat), .B(G43gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G183gat), .B2(G190gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT23), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT25), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n208), .B1(new_n212), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n223), .B(new_n209), .C1(G183gat), .C2(G190gat), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n215), .A2(new_n218), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n217), .A2(KEYINPUT25), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(KEYINPUT66), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(new_n221), .B2(new_n222), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n210), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n229), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n220), .B(new_n227), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n239), .A3(new_n237), .ZN(new_n242));
  NOR2_X1   g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(KEYINPUT26), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n218), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n243), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n241), .A2(new_n242), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n235), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(KEYINPUT1), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n252));
  INV_X1    g051(.A(G127gat), .ZN(new_n253));
  INV_X1    g052(.A(G120gat), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n254), .A2(G113gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(G113gat), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n252), .B(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G134gat), .ZN(new_n259));
  INV_X1    g058(.A(G134gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n251), .A2(new_n260), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n248), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n251), .A2(new_n260), .A3(new_n257), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n260), .B1(new_n251), .B2(new_n257), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(new_n235), .A3(new_n247), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G227gat), .A2(G233gat), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT33), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n207), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(KEYINPUT32), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n266), .A2(new_n235), .A3(new_n247), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n235), .A2(new_n247), .B1(new_n259), .B2(new_n261), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT71), .A3(new_n267), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n269), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(KEYINPUT72), .A3(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT34), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n287), .A3(new_n269), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT73), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n280), .A2(KEYINPUT72), .A3(new_n281), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT72), .B1(new_n280), .B2(new_n281), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT73), .B(new_n288), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n274), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n272), .B(new_n273), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n292), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n298), .A2(new_n299), .A3(new_n292), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT74), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT36), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n305), .B1(new_n294), .B2(new_n300), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT88), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT37), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT22), .ZN(new_n312));
  INV_X1    g111(.A(G211gat), .ZN(new_n313));
  INV_X1    g112(.A(G218gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n311), .A3(new_n315), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT29), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n248), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n235), .A2(KEYINPUT75), .A3(new_n247), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n235), .A2(new_n247), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n322), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n321), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(new_n322), .A3(new_n327), .ZN(new_n333));
  INV_X1    g132(.A(new_n321), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n248), .A2(new_n323), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n310), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G8gat), .B(G36gat), .Z(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT76), .ZN(new_n339));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  OAI21_X1  g140(.A(new_n309), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n336), .ZN(new_n343));
  INV_X1    g142(.A(new_n327), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT75), .B1(new_n235), .B2(new_n247), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n323), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n334), .B1(new_n346), .B2(new_n330), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT37), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n341), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT88), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n310), .A3(new_n336), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT38), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n354));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  INV_X1    g154(.A(G155gat), .ZN(new_n356));
  INV_X1    g155(.A(G162gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(KEYINPUT2), .ZN(new_n359));
  INV_X1    g158(.A(G141gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT77), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G141gat), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n361), .A2(new_n363), .A3(KEYINPUT78), .A4(G148gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n365));
  OR3_X1    g164(.A1(new_n365), .A2(new_n360), .A3(G148gat), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n365), .B1(new_n360), .B2(G148gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT77), .B(G141gat), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT78), .B1(new_n369), .B2(G148gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n359), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n358), .A2(new_n355), .ZN(new_n372));
  XOR2_X1   g171(.A(G141gat), .B(G148gat), .Z(new_n373));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT80), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n363), .A3(G148gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n381), .A2(new_n364), .A3(new_n367), .A4(new_n366), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n375), .B1(new_n382), .B2(new_n359), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n378), .A2(new_n385), .A3(new_n266), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n262), .A2(new_n383), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n354), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n378), .A2(new_n385), .A3(KEYINPUT3), .ZN(new_n392));
  AOI211_X1 g191(.A(KEYINPUT3), .B(new_n375), .C1(new_n382), .C2(new_n359), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n262), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n262), .A2(new_n383), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n262), .A2(new_n383), .A3(KEYINPUT81), .A4(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n391), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G1gat), .B(G29gat), .Z(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT5), .B1(new_n401), .B2(new_n397), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT83), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n404), .A2(new_n412), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n409), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n391), .A2(new_n403), .B1(new_n395), .B2(new_n411), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n410), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n414), .A2(new_n416), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n410), .B1(new_n404), .B2(new_n412), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT87), .B1(new_n422), .B2(KEYINPUT6), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n424));
  NOR4_X1   g223(.A1(new_n417), .A2(new_n424), .A3(new_n420), .A4(new_n410), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n334), .B1(new_n328), .B2(new_n331), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n333), .A2(new_n321), .A3(new_n335), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT37), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n341), .A2(KEYINPUT38), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n351), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n332), .A2(new_n336), .A3(new_n341), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n353), .A2(new_n421), .A3(new_n426), .A4(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n392), .A2(new_n394), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n401), .A2(new_n397), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT39), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n390), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n410), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT39), .B1(new_n388), .B2(new_n390), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n389), .B1(new_n436), .B2(new_n437), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n435), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n409), .B1(new_n443), .B2(new_n439), .ZN(new_n446));
  INV_X1    g245(.A(new_n435), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n446), .B(new_n447), .C1(new_n443), .C2(new_n442), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n445), .A2(new_n448), .A3(new_n416), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n349), .B1(new_n343), .B2(new_n347), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n332), .A2(new_n336), .A3(new_n452), .A4(new_n341), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457));
  INV_X1    g256(.A(G50gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n371), .A2(new_n461), .A3(new_n376), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n321), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G228gat), .ZN(new_n465));
  INV_X1    g264(.A(G233gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT3), .B1(new_n321), .B2(new_n463), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n383), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n469), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n378), .A2(new_n385), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n334), .B1(new_n393), .B2(KEYINPUT29), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n475), .B2(new_n467), .ZN(new_n476));
  INV_X1    g275(.A(G22gat), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT85), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n479));
  OAI21_X1  g278(.A(G22gat), .B1(new_n479), .B2(new_n471), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n460), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n464), .A2(new_n470), .ZN(new_n483));
  AOI211_X1 g282(.A(KEYINPUT80), .B(new_n375), .C1(new_n382), .C2(new_n359), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n384), .B1(new_n371), .B2(new_n376), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n464), .B1(new_n486), .B2(new_n472), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n483), .B(new_n477), .C1(new_n487), .C2(new_n468), .ZN(new_n488));
  AND4_X1   g287(.A1(new_n482), .A2(new_n480), .A3(new_n460), .A4(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n456), .B1(new_n481), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n480), .A2(new_n488), .A3(new_n482), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n459), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n478), .A2(new_n460), .A3(new_n480), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n455), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n449), .A2(new_n454), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n422), .A2(KEYINPUT6), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n421), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n454), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n490), .A2(new_n494), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n434), .A2(new_n495), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n306), .A2(new_n308), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n426), .A2(new_n421), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n454), .A2(KEYINPUT35), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n504), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n304), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n454), .B1(new_n421), .B2(new_n496), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n508), .A2(new_n300), .A3(new_n294), .A4(new_n500), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n503), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT16), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(G1gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(G1gat), .B2(new_n513), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n516), .B(G8gat), .Z(new_n517));
  INV_X1    g316(.A(KEYINPUT21), .ZN(new_n518));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(G71gat), .A2(G78gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT9), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n522), .B(new_n521), .C1(new_n519), .C2(new_n524), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n517), .B1(new_n518), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT95), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n518), .ZN(new_n531));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT94), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G183gat), .B(G211gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n535), .A2(new_n536), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n535), .B2(new_n536), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G190gat), .B(G218gat), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(G29gat), .A2(G36gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(KEYINPUT90), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT90), .B(KEYINPUT14), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(new_n548), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n552), .A2(KEYINPUT91), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n554), .B(new_n550), .C1(new_n551), .C2(new_n548), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n458), .A2(G43gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT15), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n458), .A2(G43gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n557), .A2(KEYINPUT92), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(KEYINPUT92), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n558), .ZN(new_n566));
  NAND2_X1  g365(.A1(G29gat), .A2(G36gat), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n552), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n556), .A2(new_n562), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT17), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n566), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n561), .B1(new_n553), .B2(new_n555), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(KEYINPUT8), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(KEYINPUT97), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G106gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n203), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n577), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n577), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n578), .A2(new_n587), .A3(new_n579), .A4(new_n582), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT98), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(KEYINPUT98), .A3(new_n588), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n575), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n591), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n556), .A2(new_n562), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n572), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n595), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n547), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT96), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n593), .A2(new_n599), .A3(new_n547), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n605), .ZN(new_n608));
  INV_X1    g407(.A(new_n606), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(new_n600), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n545), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n516), .B(G8gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n517), .B1(new_n569), .B2(KEYINPUT17), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n573), .A2(new_n574), .A3(new_n571), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n614), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT18), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n570), .A2(new_n575), .A3(new_n517), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n622), .A2(KEYINPUT18), .A3(new_n614), .A4(new_n616), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n517), .A2(new_n569), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n614), .B(KEYINPUT13), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT89), .B(G197gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT11), .B(G169gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n621), .A2(new_n623), .A3(new_n627), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n619), .A2(new_n620), .B1(new_n625), .B2(new_n626), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n637), .A2(KEYINPUT93), .A3(new_n623), .A4(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n623), .ZN(new_n639));
  INV_X1    g438(.A(new_n633), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n636), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G230gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n466), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n586), .A2(new_n588), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n526), .A2(new_n527), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n528), .A2(new_n586), .A3(new_n588), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n645), .A4(new_n591), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n648), .A2(new_n642), .A3(new_n466), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OR3_X1    g456(.A1(new_n652), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n657), .B1(new_n652), .B2(new_n653), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n613), .A2(new_n641), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n512), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n497), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n454), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT16), .B(G8gat), .ZN(new_n669));
  OR3_X1    g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n667), .A2(G8gat), .ZN(new_n674));
  OAI22_X1  g473(.A1(new_n674), .A2(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(G1325gat));
  AOI21_X1  g475(.A(G15gat), .B1(new_n663), .B2(new_n304), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n307), .B1(new_n304), .B2(new_n305), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G15gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT100), .Z(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n663), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n662), .A2(new_n500), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  AOI21_X1  g484(.A(new_n612), .B1(new_n503), .B2(new_n511), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n545), .A2(new_n641), .A3(new_n660), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689));
  INV_X1    g488(.A(G29gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n664), .A2(new_n690), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n688), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n426), .A2(new_n421), .A3(new_n433), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n352), .A2(KEYINPUT38), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n495), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n499), .A2(new_n501), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT36), .B1(new_n301), .B2(new_n303), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(new_n702), .A3(new_n307), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n304), .A2(new_n506), .B1(new_n509), .B2(KEYINPUT35), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n503), .A2(new_n706), .A3(new_n511), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n612), .A2(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n512), .A2(new_n611), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT44), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n705), .A2(new_n713), .A3(new_n707), .A4(new_n708), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n664), .A3(new_n687), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n696), .B1(new_n690), .B2(new_n717), .ZN(G1328gat));
  NOR3_X1   g517(.A1(new_n688), .A2(G36gat), .A3(new_n498), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT46), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n715), .A2(new_n454), .A3(new_n687), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT105), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G36gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(KEYINPUT105), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(G1329gat));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n503), .A2(new_n706), .A3(new_n511), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n706), .B1(new_n503), .B2(new_n511), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n713), .B1(new_n732), .B2(new_n708), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n712), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n679), .B(new_n687), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n688), .ZN(new_n737));
  INV_X1    g536(.A(new_n304), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(G43gat), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n737), .A2(new_n739), .B1(new_n726), .B2(new_n727), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n729), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n740), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n728), .B(new_n742), .C1(new_n735), .C2(G43gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(new_n743), .ZN(G1330gat));
  NAND4_X1  g543(.A1(new_n715), .A2(G50gat), .A3(new_n501), .A4(new_n687), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n500), .B1(new_n688), .B2(KEYINPUT107), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(KEYINPUT107), .B2(new_n688), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n458), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT48), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n745), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1331gat));
  NAND2_X1  g552(.A1(new_n636), .A2(new_n638), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n639), .A2(new_n640), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n660), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n613), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n705), .A2(new_n707), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n497), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT108), .B(G57gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1332gat));
  OR2_X1    g561(.A1(new_n759), .A2(KEYINPUT109), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(KEYINPUT109), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n454), .B(KEYINPUT110), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n763), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n768), .B(new_n769), .Z(G1333gat));
  NAND4_X1  g569(.A1(new_n763), .A2(G71gat), .A3(new_n679), .A4(new_n764), .ZN(new_n771));
  INV_X1    g570(.A(G71gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n759), .B2(new_n738), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g574(.A1(new_n763), .A2(new_n501), .A3(new_n764), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n545), .A2(new_n756), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n757), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n715), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n664), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G85gat), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT51), .B1(new_n711), .B2(new_n779), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n686), .A2(new_n785), .A3(new_n778), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n660), .A3(new_n786), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n787), .A2(G85gat), .A3(new_n497), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n788), .ZN(G1336gat));
  NOR3_X1   g588(.A1(new_n787), .A2(G92gat), .A3(new_n766), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n715), .A2(new_n765), .A3(new_n780), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G92gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n715), .A2(new_n454), .A3(new_n780), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n790), .B1(new_n795), .B2(G92gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(G1337gat));
  NOR2_X1   g597(.A1(new_n678), .A2(new_n203), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n787), .A2(new_n738), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n781), .A2(new_n799), .B1(new_n800), .B2(new_n203), .ZN(G1338gat));
  NAND4_X1  g600(.A1(new_n715), .A2(G106gat), .A3(new_n501), .A4(new_n780), .ZN(new_n802));
  NAND2_X1  g601(.A1(KEYINPUT111), .A2(KEYINPUT53), .ZN(new_n803));
  NOR2_X1   g602(.A1(KEYINPUT111), .A2(KEYINPUT53), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n784), .A2(new_n501), .A3(new_n660), .A4(new_n786), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n584), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n802), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n803), .B1(new_n802), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(G1339gat));
  NAND4_X1  g608(.A1(new_n545), .A2(new_n641), .A3(new_n612), .A4(new_n757), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n656), .B1(new_n652), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n645), .A2(KEYINPUT10), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n594), .A2(new_n814), .A3(new_n589), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT10), .B1(new_n646), .B2(new_n647), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n815), .A2(new_n816), .B1(new_n642), .B2(new_n466), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n650), .A2(new_n643), .A3(new_n651), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT54), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n813), .A2(new_n819), .A3(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n658), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n813), .A2(new_n819), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(new_n813), .B2(new_n819), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n821), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n622), .A2(new_n616), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n830), .A2(new_n614), .B1(new_n625), .B2(new_n626), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n636), .A2(new_n638), .B1(new_n632), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n832), .A3(new_n611), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n756), .A2(new_n829), .B1(new_n832), .B2(new_n660), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n611), .ZN(new_n835));
  INV_X1    g634(.A(new_n545), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n811), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n294), .A2(new_n300), .A3(new_n500), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n837), .A2(new_n497), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n766), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT113), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n641), .A2(G113gat), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n304), .A2(new_n500), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n765), .A2(new_n497), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n641), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n849), .ZN(G1340gat));
  NAND3_X1  g649(.A1(new_n841), .A2(new_n254), .A3(new_n660), .ZN(new_n851));
  OAI21_X1  g650(.A(G120gat), .B1(new_n848), .B2(new_n757), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1341gat));
  NOR3_X1   g652(.A1(new_n848), .A2(new_n253), .A3(new_n836), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n840), .A2(new_n836), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(KEYINPUT115), .ZN(new_n856));
  AOI21_X1  g655(.A(G127gat), .B1(new_n855), .B2(KEYINPUT115), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(G1342gat));
  OAI21_X1  g657(.A(G134gat), .B1(new_n848), .B2(new_n612), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n454), .A2(new_n612), .ZN(new_n860));
  XOR2_X1   g659(.A(KEYINPUT68), .B(G134gat), .Z(new_n861));
  NAND3_X1  g660(.A1(new_n839), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(KEYINPUT116), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(KEYINPUT116), .ZN(new_n865));
  OAI221_X1 g664(.A(new_n859), .B1(KEYINPUT56), .B2(new_n862), .C1(new_n864), .C2(new_n865), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n835), .A2(new_n836), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n497), .B1(new_n867), .B2(new_n810), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n702), .A2(new_n307), .A3(new_n500), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT120), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n756), .A2(new_n360), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(KEYINPUT120), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n871), .A2(new_n766), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n678), .A2(new_n847), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n831), .A2(new_n632), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n754), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n820), .A2(new_n658), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n825), .B(KEYINPUT55), .C1(new_n813), .C2(new_n819), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n880), .B(new_n611), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n754), .A2(new_n660), .A3(new_n878), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n641), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n884), .B1(new_n887), .B2(new_n612), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n810), .B1(new_n888), .B2(new_n545), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n889), .B2(new_n501), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n501), .A2(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n821), .B2(new_n827), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n880), .A2(KEYINPUT117), .A3(new_n824), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n756), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n611), .B1(new_n895), .B2(new_n885), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n836), .B1(new_n896), .B2(new_n884), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n891), .B1(new_n897), .B2(new_n810), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n756), .B(new_n877), .C1(new_n890), .C2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n369), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n875), .A2(new_n876), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n678), .A2(new_n847), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n897), .A2(new_n810), .ZN(new_n904));
  INV_X1    g703(.A(new_n891), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n837), .B2(new_n500), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n369), .B1(new_n909), .B2(new_n756), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n765), .A2(new_n872), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n868), .A2(new_n869), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT118), .A4(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT119), .B(KEYINPUT58), .C1(new_n910), .C2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n914), .A3(new_n915), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT119), .B1(new_n919), .B2(KEYINPUT58), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n902), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT121), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n923), .B(new_n902), .C1(new_n918), .C2(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1344gat));
  AOI21_X1  g724(.A(new_n500), .B1(new_n897), .B2(new_n810), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n926), .A2(KEYINPUT57), .B1(new_n837), .B2(new_n891), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n660), .A3(new_n877), .ZN(new_n928));
  AND2_X1   g727(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n906), .A2(new_n908), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n903), .A2(KEYINPUT59), .A3(new_n757), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n928), .A2(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n871), .A2(new_n874), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n934), .A2(new_n766), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n935), .B2(new_n660), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n936), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n356), .A3(new_n545), .ZN(new_n938));
  INV_X1    g737(.A(new_n909), .ZN(new_n939));
  OAI21_X1  g738(.A(G155gat), .B1(new_n939), .B2(new_n836), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1346gat));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n357), .A3(new_n860), .ZN(new_n942));
  OAI21_X1  g741(.A(G162gat), .B1(new_n939), .B2(new_n612), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1347gat));
  NOR2_X1   g743(.A1(new_n837), .A2(new_n664), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n766), .A2(new_n838), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n756), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n664), .A2(new_n498), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n837), .A2(new_n845), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n641), .A2(new_n213), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(G1348gat));
  NAND3_X1  g754(.A1(new_n953), .A2(G176gat), .A3(new_n660), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n948), .A2(new_n660), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT123), .A3(new_n214), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT123), .B1(new_n957), .B2(new_n214), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT124), .ZN(G1349gat));
  NAND2_X1  g760(.A1(new_n953), .A2(new_n545), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G183gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n236), .A3(new_n545), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g765(.A(new_n237), .B1(new_n953), .B2(new_n611), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(KEYINPUT61), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n948), .A2(new_n237), .A3(new_n611), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n971), .B(new_n972), .C1(KEYINPUT61), .C2(new_n969), .ZN(G1351gat));
  NAND3_X1  g772(.A1(new_n945), .A2(new_n869), .A3(new_n765), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G197gat), .B1(new_n975), .B2(new_n756), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n679), .A2(new_n951), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n927), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n756), .A2(G197gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1352gat));
  NOR3_X1   g779(.A1(new_n974), .A2(G204gat), .A3(new_n757), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n978), .A2(new_n660), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G204gat), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1353gat));
  NAND3_X1  g784(.A1(new_n975), .A2(new_n313), .A3(new_n545), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n978), .A2(new_n545), .ZN(new_n987));
  AND2_X1   g786(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n988));
  OAI21_X1  g787(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n988), .B1(new_n987), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  NAND3_X1  g792(.A1(new_n975), .A2(new_n314), .A3(new_n611), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n611), .ZN(new_n995));
  INV_X1    g794(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n994), .B1(new_n996), .B2(new_n314), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


