//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n441, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  AND2_X1   g014(.A1(KEYINPUT65), .A2(G57), .ZN(new_n440));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(G57), .ZN(new_n441));
  NOR2_X1   g016(.A1(new_n440), .A2(new_n441), .ZN(G237));
  XOR2_X1   g017(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(new_n454), .B2(G2106), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n471), .B1(new_n465), .B2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n463), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G137), .A4(new_n466), .ZN(new_n474));
  NAND2_X1  g049(.A1(G101), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n470), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI211_X1 g053(.A(KEYINPUT69), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(G160));
  AND3_X1   g055(.A1(new_n472), .A2(new_n466), .A3(new_n473), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(KEYINPUT70), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n481), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n494), .B2(G124), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n489), .A2(new_n495), .ZN(G162));
  AND2_X1   g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n472), .A2(new_n473), .A3(new_n466), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G102), .A2(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(G2105), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n472), .A2(new_n473), .A3(G126), .A4(new_n466), .ZN(new_n501));
  NAND2_X1  g076(.A1(G114), .A2(G2104), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n482), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n482), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n500), .A2(new_n503), .A3(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT73), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n508), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n516), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n515), .B1(new_n523), .B2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n516), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT74), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n517), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AOI22_X1  g114(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n508), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n517), .A2(new_n542), .B1(new_n528), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n517), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n508), .ZN(new_n549));
  AOI211_X1 g124(.A(new_n547), .B(new_n549), .C1(G43), .C2(new_n520), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND3_X1  g130(.A1(new_n520), .A2(KEYINPUT9), .A3(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n528), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n556), .A2(KEYINPUT75), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n511), .A2(G65), .ZN(new_n564));
  INV_X1    g139(.A(G78), .ZN(new_n565));
  INV_X1    g140(.A(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT76), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT76), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n518), .B2(G91), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n562), .A2(new_n563), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  NAND2_X1  g147(.A1(new_n523), .A2(new_n525), .ZN(new_n573));
  INV_X1    g148(.A(new_n515), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G303));
  NAND2_X1  g150(.A1(new_n518), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n520), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n576), .A2(KEYINPUT77), .A3(new_n578), .A4(new_n577), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G288));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n509), .B2(new_n510), .ZN(new_n586));
  AND2_X1   g161(.A1(G73), .A2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n517), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n508), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT78), .B(G85), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n517), .A2(new_n597), .B1(new_n528), .B2(new_n598), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n596), .A2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n511), .A2(new_n516), .A3(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n511), .A2(G66), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n605), .B2(new_n566), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n605), .A2(new_n566), .A3(KEYINPUT79), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n601), .B1(new_n610), .B2(G868), .ZN(G321));
  XNOR2_X1  g186(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  XNOR2_X1  g191(.A(KEYINPUT81), .B(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(G860), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g194(.A1(new_n610), .A2(new_n617), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g198(.A1(new_n482), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2100), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  NOR3_X1   g207(.A1(new_n482), .A2(KEYINPUT84), .A3(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT84), .B1(new_n482), .B2(G111), .ZN(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(G2104), .A3(new_n635), .ZN(new_n636));
  OAI22_X1  g211(.A1(new_n493), .A2(new_n632), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n487), .B2(G135), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n629), .A2(new_n630), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  OAI221_X1 g214(.A(new_n639), .B1(new_n631), .B2(new_n638), .C1(new_n626), .C2(new_n630), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT85), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT86), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n644), .B2(new_n645), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n652), .B2(new_n655), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT87), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n665), .B(new_n662), .C1(new_n659), .C2(new_n661), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n661), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n667), .A2(new_n662), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n631), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(G2096), .ZN(new_n673));
  INV_X1    g248(.A(G2100), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n678), .A2(new_n679), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n682), .A3(new_n680), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n682), .C2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  INV_X1    g264(.A(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n688), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT89), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NOR2_X1   g272(.A1(G168), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n697), .B2(G21), .ZN(new_n699));
  INV_X1    g274(.A(G1966), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT99), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G2084), .ZN(new_n704));
  NAND2_X1  g279(.A1(G160), .A2(G29), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT24), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G34), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(KEYINPUT96), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(G34), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n708), .B2(KEYINPUT96), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n703), .B1(new_n704), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n697), .A2(G20), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G299), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1956), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n713), .B(new_n718), .C1(new_n704), .C2(new_n712), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n706), .A2(G35), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G162), .B2(new_n706), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT29), .Z(new_n722));
  INV_X1    g297(.A(G2090), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n610), .A2(new_n697), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G4), .B2(new_n697), .ZN(new_n726));
  INV_X1    g301(.A(G1348), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n697), .A2(G19), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n550), .B2(new_n697), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1341), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n706), .A2(G33), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  INV_X1    g309(.A(new_n467), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n735), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(new_n736), .B2(new_n482), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n487), .B2(G139), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(new_n706), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G2072), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(new_n727), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n728), .A2(new_n731), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n638), .A2(G29), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT98), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G28), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n706), .B1(new_n746), .B2(G28), .ZN(new_n748));
  AND2_X1   g323(.A1(KEYINPUT31), .A2(G11), .ZN(new_n749));
  NOR2_X1   g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n697), .A2(G5), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G171), .B2(new_n697), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n751), .B1(new_n753), .B2(G1961), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n745), .B(new_n754), .C1(G1961), .C2(new_n753), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n699), .A2(new_n700), .B1(new_n744), .B2(new_n743), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n742), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n739), .A2(G2072), .ZN(new_n758));
  NAND2_X1  g333(.A1(G164), .A2(G29), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G27), .B2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n758), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n706), .A2(G32), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND3_X1  g342(.A1(new_n482), .A2(G105), .A3(G2104), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n767), .B(new_n768), .C1(new_n493), .C2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n485), .A2(new_n486), .ZN(new_n771));
  INV_X1    g346(.A(G141), .ZN(new_n772));
  OAI21_X1  g347(.A(KEYINPUT97), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n487), .A2(new_n774), .A3(G141), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n770), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n765), .B1(new_n776), .B2(new_n706), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT27), .B(G1996), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n757), .A2(new_n764), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n706), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT28), .ZN(new_n783));
  INV_X1    g358(.A(G128), .ZN(new_n784));
  NOR2_X1   g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(new_n482), .B2(G116), .ZN(new_n786));
  OAI22_X1  g361(.A1(new_n493), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n487), .B2(G140), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(new_n706), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT95), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n719), .A2(new_n724), .A3(new_n780), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n697), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(new_n579), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n697), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT92), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(G166), .A2(G16), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G16), .B2(G22), .ZN(new_n800));
  INV_X1    g375(.A(G1971), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n796), .A2(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  NOR2_X1   g378(.A1(G6), .A2(G16), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n593), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT32), .B(G1981), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n796), .B2(new_n798), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n706), .A2(G25), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n481), .A2(G119), .A3(G2105), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT90), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(G107), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n463), .B1(new_n816), .B2(G2105), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n487), .A2(G131), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n812), .B1(new_n821), .B2(new_n706), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n822), .A2(new_n824), .ZN(new_n826));
  NOR2_X1   g401(.A1(G16), .A2(G24), .ZN(new_n827));
  XNOR2_X1  g402(.A(G290), .B(KEYINPUT91), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(G16), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1986), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n810), .A2(new_n811), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT93), .B(KEYINPUT36), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n722), .A2(new_n723), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n722), .A2(KEYINPUT100), .A3(new_n723), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n832), .A2(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(KEYINPUT93), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n810), .A2(new_n840), .A3(new_n811), .A4(new_n831), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n792), .A2(new_n838), .A3(new_n841), .ZN(G150));
  INV_X1    g417(.A(G150), .ZN(G311));
  AOI22_X1  g418(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n508), .ZN(new_n845));
  INV_X1    g420(.A(G93), .ZN(new_n846));
  INV_X1    g421(.A(G55), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n517), .A2(new_n846), .B1(new_n528), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n550), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n550), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT38), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n610), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  INV_X1    g431(.A(G860), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n849), .A2(new_n857), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G145));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n487), .A2(G140), .ZN(new_n864));
  OAI21_X1  g439(.A(G164), .B1(new_n864), .B2(new_n787), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n498), .A2(new_n499), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n482), .ZN(new_n867));
  INV_X1    g442(.A(new_n506), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n501), .A2(new_n502), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G2105), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n788), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n873), .A2(new_n776), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n776), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n738), .A2(KEYINPUT102), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n776), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n865), .A3(new_n872), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n873), .A2(new_n776), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(G118), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n883), .A2(KEYINPUT104), .B1(new_n884), .B2(G2105), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(KEYINPUT104), .B2(new_n883), .ZN(new_n886));
  INV_X1    g461(.A(G130), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n493), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  INV_X1    g464(.A(G142), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n771), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n487), .A2(KEYINPUT103), .A3(G142), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n625), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n896), .A2(new_n820), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n891), .A2(new_n892), .ZN(new_n899));
  INV_X1    g474(.A(new_n888), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n625), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n821), .B1(new_n902), .B2(new_n895), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n878), .A2(new_n882), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n877), .B1(new_n874), .B2(new_n875), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n820), .B1(new_n896), .B2(new_n897), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n880), .A2(new_n881), .A3(new_n876), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n821), .A3(new_n895), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G162), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n638), .B(G160), .ZN(new_n913));
  INV_X1    g488(.A(G162), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n904), .A2(new_n909), .A3(new_n910), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n913), .B1(new_n912), .B2(new_n915), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n863), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n915), .ZN(new_n921));
  INV_X1    g496(.A(new_n913), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(KEYINPUT40), .A3(new_n917), .A4(new_n916), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n920), .A2(new_n924), .ZN(G395));
  INV_X1    g500(.A(G290), .ZN(new_n926));
  XNOR2_X1  g501(.A(G166), .B(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n579), .B(new_n593), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n929), .B(KEYINPUT42), .Z(new_n930));
  XNOR2_X1  g505(.A(new_n620), .B(KEYINPUT106), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(new_n852), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n610), .A2(G299), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n610), .A2(G299), .A3(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n610), .A2(G299), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(KEYINPUT41), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  INV_X1    g516(.A(new_n933), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n941), .B1(new_n942), .B2(new_n938), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n932), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n938), .B1(new_n935), .B2(new_n936), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n946), .B2(new_n932), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n930), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(G868), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(G868), .B2(new_n849), .ZN(G295));
  OAI21_X1  g525(.A(new_n949), .B1(G868), .B2(new_n849), .ZN(G331));
  NAND2_X1  g526(.A1(G168), .A2(G301), .ZN(new_n952));
  NAND2_X1  g527(.A1(G286), .A2(G171), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n850), .A2(new_n952), .A3(new_n851), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n852), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n946), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n954), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n944), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n960), .B2(new_n929), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n937), .A2(new_n939), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n941), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n939), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n946), .B2(KEYINPUT41), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n957), .B1(new_n968), .B2(new_n959), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n961), .B(new_n962), .C1(new_n929), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n929), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n968), .A2(new_n959), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n957), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(KEYINPUT109), .A3(new_n962), .A4(new_n961), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n961), .B1(new_n929), .B2(new_n960), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n975), .A2(KEYINPUT43), .A3(new_n961), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n962), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT44), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n985), .ZN(G397));
  OAI21_X1  g561(.A(KEYINPUT115), .B1(G164), .B2(G1384), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n871), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G40), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n478), .A2(new_n991), .A3(new_n479), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n987), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT116), .B(G8), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n794), .A2(G1976), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT52), .ZN(new_n998));
  INV_X1    g573(.A(G1976), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n581), .A2(new_n999), .A3(new_n582), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1002), .A2(new_n995), .A3(new_n993), .A4(new_n996), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n592), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n690), .A3(new_n588), .ZN(new_n1006));
  OAI21_X1  g581(.A(G1981), .B1(new_n589), .B2(new_n592), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT49), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(new_n995), .A3(new_n993), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1012), .A2(new_n993), .A3(KEYINPUT117), .A4(new_n995), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1004), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(G303), .B2(G8), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  NOR3_X1   g597(.A1(G166), .A2(KEYINPUT55), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n476), .A2(new_n477), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n476), .A2(new_n477), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(G40), .A3(new_n1026), .A4(new_n470), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n871), .A2(new_n989), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(KEYINPUT50), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n987), .A2(new_n1030), .A3(new_n990), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G2090), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n869), .A2(G2105), .B1(new_n505), .B2(new_n504), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n1035), .B2(new_n867), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT114), .B(new_n1037), .C1(G164), .C2(G1384), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n1042));
  NOR3_X1   g617(.A1(G164), .A2(new_n1042), .A3(G1384), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n1027), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1971), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1024), .B(G8), .C1(new_n1033), .C2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G288), .A2(G1976), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1017), .A2(new_n1047), .B1(new_n690), .B2(new_n593), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n993), .A2(new_n995), .ZN(new_n1049));
  XOR2_X1   g624(.A(new_n1049), .B(KEYINPUT118), .Z(new_n1050));
  OAI22_X1  g625(.A1(new_n1019), .A2(new_n1046), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1037), .A2(G1384), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NOR3_X1   g629(.A1(G164), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT119), .B1(new_n871), .B2(new_n1053), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n992), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT45), .B1(new_n987), .B2(new_n990), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G2078), .ZN(new_n1061));
  INV_X1    g636(.A(G1961), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1059), .A2(new_n1061), .B1(new_n1032), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1041), .A2(new_n1044), .A3(new_n761), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1060), .ZN(new_n1065));
  AOI21_X1  g640(.A(G301), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1030), .B1(new_n987), .B2(new_n990), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n992), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1067), .A2(new_n1068), .A3(G2090), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n995), .B1(new_n1069), .B2(new_n1045), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1024), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1018), .A2(new_n1066), .A3(new_n1072), .A4(new_n1046), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n700), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT120), .B(new_n700), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1029), .A2(new_n1031), .A3(new_n704), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G286), .A2(new_n995), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1074), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1084));
  NOR3_X1   g659(.A1(G164), .A2(KEYINPUT115), .A3(G1384), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n988), .B1(new_n871), .B2(new_n989), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1042), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1052), .B1(G164), .B2(new_n1054), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n871), .A2(KEYINPUT119), .A3(new_n1053), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1027), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1966), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1079), .B1(new_n1091), .B2(KEYINPUT120), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1078), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n995), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT51), .B1(G286), .B2(new_n995), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1083), .A2(new_n1084), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1073), .B1(new_n1096), .B2(KEYINPUT62), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1082), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(KEYINPUT51), .A3(new_n1084), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1051), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1956), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1041), .A2(new_n1044), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n570), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(new_n560), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1106), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1112), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1106), .A2(new_n1108), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1114), .B(new_n1115), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n610), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n993), .A2(KEYINPUT122), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n987), .A2(new_n990), .A3(new_n992), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G2067), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1120), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1119), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1041), .A2(new_n1044), .A3(new_n1107), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT50), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1027), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1956), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT123), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1106), .A2(new_n1108), .A3(new_n1116), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1114), .B1(new_n1138), .B2(new_n1115), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1113), .B1(new_n1131), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1115), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT125), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT58), .B(G1341), .Z(new_n1144));
  NAND3_X1  g719(.A1(new_n1121), .A2(new_n1123), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G1996), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1041), .A2(new_n1044), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n550), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1142), .A2(new_n1143), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(KEYINPUT59), .A3(new_n550), .ZN(new_n1152));
  AOI21_X1  g727(.A(G2067), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1153), .A2(new_n610), .A3(new_n1127), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT60), .B1(new_n1129), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1113), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1156), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1106), .A2(new_n1108), .A3(new_n1112), .A4(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1153), .A2(new_n1127), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1120), .A2(KEYINPUT60), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1157), .A2(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1151), .A2(new_n1152), .A3(new_n1155), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1140), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1032), .A2(new_n1062), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1028), .A2(new_n1037), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1044), .A2(new_n1167), .A3(new_n1061), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1064), .A2(new_n1060), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1169), .A2(new_n1170), .A3(G171), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1165), .B1(new_n1171), .B2(new_n1066), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT126), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1174), .B(new_n1165), .C1(new_n1171), .C2(new_n1066), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(G171), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1063), .A2(G301), .A3(new_n1065), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(KEYINPUT54), .A3(new_n1178), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1046), .A2(new_n1004), .A3(new_n1017), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(new_n1180), .A3(new_n1072), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1181), .A2(new_n1101), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1164), .A2(new_n1176), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1072), .A2(new_n1046), .A3(new_n1004), .A4(new_n1017), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1080), .A2(G168), .A3(new_n995), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g764(.A(KEYINPUT121), .B(new_n1184), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1186), .ZN(new_n1191));
  OAI21_X1  g766(.A(G8), .B1(new_n1033), .B2(new_n1045), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1184), .B1(new_n1192), .B2(new_n1071), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1191), .A2(new_n1180), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1189), .A2(new_n1190), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1104), .A2(new_n1183), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n992), .A2(new_n1028), .A3(new_n1037), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(KEYINPUT112), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT112), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1202), .A2(G1996), .A3(new_n879), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT113), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1203), .B(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1198), .A2(new_n1146), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n879), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n788), .B(new_n1125), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1207), .B1(new_n1202), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1202), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n820), .B(new_n823), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1205), .B(new_n1209), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  AND2_X1   g787(.A1(G290), .A2(G1986), .ZN(new_n1213));
  NOR2_X1   g788(.A1(G290), .A2(G1986), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1198), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  XOR2_X1   g790(.A(new_n1215), .B(KEYINPUT111), .Z(new_n1216));
  NOR2_X1   g791(.A1(new_n1212), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1196), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1202), .B1(new_n879), .B2(new_n1208), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1206), .B(KEYINPUT46), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT47), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1198), .A2(new_n1214), .ZN(new_n1223));
  XOR2_X1   g798(.A(new_n1223), .B(KEYINPUT48), .Z(new_n1224));
  OAI21_X1  g799(.A(new_n1222), .B1(new_n1212), .B2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1205), .A2(new_n823), .A3(new_n821), .A4(new_n1209), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n788), .A2(new_n1125), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1210), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1218), .A2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g805(.A1(new_n672), .A2(new_n675), .A3(G319), .ZN(new_n1232));
  NOR2_X1   g806(.A1(G229), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g807(.A(new_n1233), .B1(new_n657), .B2(new_n656), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n1234), .A2(KEYINPUT127), .ZN(new_n1235));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1236));
  OAI211_X1 g810(.A(new_n1233), .B(new_n1236), .C1(new_n657), .C2(new_n656), .ZN(new_n1237));
  NAND2_X1  g811(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n923), .A2(new_n917), .A3(new_n916), .ZN(new_n1239));
  AND3_X1   g813(.A1(new_n1238), .A2(new_n1239), .A3(new_n979), .ZN(G308));
  NAND3_X1  g814(.A1(new_n1238), .A2(new_n1239), .A3(new_n979), .ZN(G225));
endmodule


