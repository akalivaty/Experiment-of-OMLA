

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(n743), .ZN(n759) );
  NOR2_X1 U555 ( .A1(n772), .A2(n771), .ZN(n775) );
  BUF_X1 U556 ( .A(n635), .Z(n636) );
  XNOR2_X1 U557 ( .A(n531), .B(n530), .ZN(n629) );
  NOR2_X2 U558 ( .A1(G2104), .A2(n537), .ZN(n916) );
  INV_X1 U559 ( .A(KEYINPUT65), .ZN(n783) );
  NAND2_X1 U560 ( .A1(n629), .A2(G113), .ZN(n532) );
  NOR2_X1 U561 ( .A1(n753), .A2(n752), .ZN(n754) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n735) );
  XNOR2_X1 U563 ( .A(n798), .B(KEYINPUT105), .ZN(n801) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n820) );
  INV_X1 U565 ( .A(KEYINPUT68), .ZN(n530) );
  XOR2_X1 U566 ( .A(KEYINPUT17), .B(n529), .Z(n635) );
  NOR2_X1 U567 ( .A1(G651), .A2(n671), .ZN(n676) );
  NOR2_X2 U568 ( .A1(n541), .A2(n540), .ZN(G160) );
  AND2_X1 U569 ( .A1(n744), .A2(G8), .ZN(n522) );
  AND2_X1 U570 ( .A1(n527), .A2(n999), .ZN(n523) );
  AND2_X1 U571 ( .A1(n831), .A2(n840), .ZN(n524) );
  XOR2_X1 U572 ( .A(KEYINPUT31), .B(KEYINPUT102), .Z(n525) );
  AND2_X1 U573 ( .A1(n743), .A2(G1341), .ZN(n526) );
  OR2_X1 U574 ( .A1(n788), .A2(n777), .ZN(n527) );
  OR2_X1 U575 ( .A1(n777), .A2(n800), .ZN(n528) );
  NOR2_X1 U576 ( .A1(n743), .A2(n963), .ZN(n713) );
  AND2_X1 U577 ( .A1(n715), .A2(n714), .ZN(n721) );
  BUF_X1 U578 ( .A(n743), .Z(n757) );
  INV_X1 U579 ( .A(KEYINPUT30), .ZN(n748) );
  NOR2_X1 U580 ( .A1(n759), .A2(n745), .ZN(n772) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  NAND2_X1 U582 ( .A1(G160), .A2(G40), .ZN(n819) );
  INV_X1 U583 ( .A(G651), .ZN(n567) );
  INV_X1 U584 ( .A(G2105), .ZN(n537) );
  BUF_X1 U585 ( .A(n629), .Z(n917) );
  NOR2_X1 U586 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U587 ( .A(n551), .B(n550), .ZN(G164) );
  NAND2_X1 U588 ( .A1(n635), .A2(G137), .ZN(n533) );
  NAND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U591 ( .A(n534), .B(KEYINPUT69), .ZN(n536) );
  NAND2_X1 U592 ( .A1(G125), .A2(n916), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n537), .A2(G2104), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n538), .B(KEYINPUT67), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G101), .A2(n920), .ZN(n539) );
  XNOR2_X1 U597 ( .A(KEYINPUT23), .B(n539), .ZN(n540) );
  INV_X1 U598 ( .A(KEYINPUT93), .ZN(n551) );
  NAND2_X1 U599 ( .A1(G126), .A2(n916), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G114), .A2(n629), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n544), .B(KEYINPUT92), .ZN(n549) );
  BUF_X2 U603 ( .A(n545), .Z(n920) );
  NAND2_X1 U604 ( .A1(G102), .A2(n920), .ZN(n547) );
  NAND2_X1 U605 ( .A1(G138), .A2(n635), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U607 ( .A(G2446), .B(G2430), .Z(n553) );
  XNOR2_X1 U608 ( .A(G2451), .B(G2454), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U610 ( .A(n554), .B(G2427), .Z(n556) );
  XNOR2_X1 U611 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n556), .B(n555), .ZN(n560) );
  XOR2_X1 U613 ( .A(G2443), .B(KEYINPUT108), .Z(n558) );
  XNOR2_X1 U614 ( .A(G2438), .B(G2435), .ZN(n557) );
  XNOR2_X1 U615 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U616 ( .A(n560), .B(n559), .Z(n561) );
  AND2_X1 U617 ( .A1(G14), .A2(n561), .ZN(G401) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U619 ( .A(G543), .B(KEYINPUT0), .Z(n562) );
  XNOR2_X1 U620 ( .A(KEYINPUT70), .B(n562), .ZN(n671) );
  NAND2_X1 U621 ( .A1(n676), .A2(G53), .ZN(n566) );
  NOR2_X1 U622 ( .A1(G543), .A2(n567), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT1), .B(n563), .Z(n564) );
  XNOR2_X2 U624 ( .A(KEYINPUT72), .B(n564), .ZN(n675) );
  NAND2_X1 U625 ( .A1(G65), .A2(n675), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n571) );
  NOR2_X1 U627 ( .A1(n567), .A2(n671), .ZN(n664) );
  NAND2_X1 U628 ( .A1(G78), .A2(n664), .ZN(n569) );
  NOR2_X1 U629 ( .A1(G651), .A2(G543), .ZN(n661) );
  NAND2_X1 U630 ( .A1(G91), .A2(n661), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n731) );
  INV_X1 U633 ( .A(n731), .ZN(G299) );
  INV_X1 U634 ( .A(G108), .ZN(G238) );
  INV_X1 U635 ( .A(G120), .ZN(G236) );
  INV_X1 U636 ( .A(G57), .ZN(G237) );
  INV_X1 U637 ( .A(G132), .ZN(G219) );
  INV_X1 U638 ( .A(G82), .ZN(G220) );
  NAND2_X1 U639 ( .A1(n661), .A2(G88), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G50), .A2(n676), .ZN(n572) );
  XOR2_X1 U641 ( .A(KEYINPUT85), .B(n572), .Z(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G75), .A2(n664), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G62), .A2(n675), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U646 ( .A1(n578), .A2(n577), .ZN(G166) );
  NAND2_X1 U647 ( .A1(n676), .A2(G51), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G63), .A2(n675), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U650 ( .A(KEYINPUT6), .B(n581), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n661), .A2(G89), .ZN(n582) );
  XNOR2_X1 U652 ( .A(n582), .B(KEYINPUT4), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G76), .A2(n664), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U655 ( .A(n585), .B(KEYINPUT5), .Z(n586) );
  NOR2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U657 ( .A(KEYINPUT7), .B(n588), .Z(n589) );
  XOR2_X1 U658 ( .A(KEYINPUT77), .B(n589), .Z(G168) );
  XOR2_X1 U659 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U660 ( .A1(G7), .A2(G661), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U662 ( .A(G567), .ZN(n706) );
  NOR2_X1 U663 ( .A1(n706), .A2(G223), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U665 ( .A1(n661), .A2(G81), .ZN(n592) );
  XNOR2_X1 U666 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G68), .A2(n664), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n595) );
  XNOR2_X1 U670 ( .A(n596), .B(n595), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G56), .A2(n675), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n597), .Z(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n676), .A2(G43), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n998) );
  INV_X1 U676 ( .A(G860), .ZN(n651) );
  OR2_X1 U677 ( .A1(n998), .A2(n651), .ZN(G153) );
  NAND2_X1 U678 ( .A1(n675), .A2(G64), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n602), .B(KEYINPUT73), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G77), .A2(n664), .ZN(n604) );
  NAND2_X1 U681 ( .A1(G90), .A2(n661), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U683 ( .A(KEYINPUT9), .B(n605), .Z(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n676), .A2(G52), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(G301) );
  NAND2_X1 U687 ( .A1(G54), .A2(n676), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G79), .A2(n664), .ZN(n611) );
  NAND2_X1 U689 ( .A1(G92), .A2(n661), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G66), .A2(n675), .ZN(n612) );
  XNOR2_X1 U692 ( .A(KEYINPUT75), .B(n612), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U695 ( .A(n617), .B(KEYINPUT15), .ZN(n618) );
  XNOR2_X2 U696 ( .A(KEYINPUT76), .B(n618), .ZN(n992) );
  INV_X1 U697 ( .A(n992), .ZN(n881) );
  NOR2_X1 U698 ( .A1(n881), .A2(G868), .ZN(n620) );
  INV_X1 U699 ( .A(G868), .ZN(n689) );
  NOR2_X1 U700 ( .A1(n689), .A2(G301), .ZN(n619) );
  NOR2_X1 U701 ( .A1(n620), .A2(n619), .ZN(G284) );
  NOR2_X1 U702 ( .A1(G286), .A2(n689), .ZN(n622) );
  NOR2_X1 U703 ( .A1(G868), .A2(G299), .ZN(n621) );
  NOR2_X1 U704 ( .A1(n622), .A2(n621), .ZN(G297) );
  NAND2_X1 U705 ( .A1(n651), .A2(G559), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n623), .A2(n992), .ZN(n624) );
  XNOR2_X1 U707 ( .A(n624), .B(KEYINPUT78), .ZN(n625) );
  XNOR2_X1 U708 ( .A(KEYINPUT16), .B(n625), .ZN(G148) );
  NOR2_X1 U709 ( .A1(G868), .A2(n998), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n992), .A2(G868), .ZN(n626) );
  NOR2_X1 U711 ( .A1(G559), .A2(n626), .ZN(n627) );
  NOR2_X1 U712 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U713 ( .A1(n917), .A2(G111), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n630), .B(KEYINPUT80), .ZN(n634) );
  XOR2_X1 U715 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n632) );
  NAND2_X1 U716 ( .A1(G123), .A2(n916), .ZN(n631) );
  XNOR2_X1 U717 ( .A(n632), .B(n631), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G99), .A2(n920), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G135), .A2(n636), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n943) );
  XNOR2_X1 U723 ( .A(n943), .B(G2096), .ZN(n642) );
  INV_X1 U724 ( .A(G2100), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(G156) );
  NAND2_X1 U726 ( .A1(n676), .A2(G55), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G67), .A2(n675), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G80), .A2(n664), .ZN(n646) );
  NAND2_X1 U730 ( .A1(G93), .A2(n661), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n690) );
  XOR2_X1 U733 ( .A(n690), .B(KEYINPUT82), .Z(n653) );
  XNOR2_X1 U734 ( .A(n998), .B(KEYINPUT81), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n992), .A2(G559), .ZN(n649) );
  XNOR2_X1 U736 ( .A(n650), .B(n649), .ZN(n687) );
  NAND2_X1 U737 ( .A1(n687), .A2(n651), .ZN(n652) );
  XNOR2_X1 U738 ( .A(n653), .B(n652), .ZN(G145) );
  NAND2_X1 U739 ( .A1(G85), .A2(n661), .ZN(n655) );
  NAND2_X1 U740 ( .A1(G60), .A2(n675), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U742 ( .A1(G72), .A2(n664), .ZN(n656) );
  XNOR2_X1 U743 ( .A(KEYINPUT71), .B(n656), .ZN(n657) );
  NOR2_X1 U744 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U745 ( .A1(n676), .A2(G47), .ZN(n659) );
  NAND2_X1 U746 ( .A1(n660), .A2(n659), .ZN(G290) );
  NAND2_X1 U747 ( .A1(G48), .A2(n676), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G86), .A2(n661), .ZN(n663) );
  NAND2_X1 U749 ( .A1(G61), .A2(n675), .ZN(n662) );
  NAND2_X1 U750 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n664), .A2(G73), .ZN(n665) );
  XOR2_X1 U752 ( .A(KEYINPUT2), .B(n665), .Z(n666) );
  NOR2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U755 ( .A(n670), .B(KEYINPUT84), .ZN(G305) );
  NAND2_X1 U756 ( .A1(G651), .A2(G74), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G87), .A2(n671), .ZN(n672) );
  NAND2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U760 ( .A1(G49), .A2(n676), .ZN(n677) );
  XOR2_X1 U761 ( .A(KEYINPUT83), .B(n677), .Z(n678) );
  NAND2_X1 U762 ( .A1(n679), .A2(n678), .ZN(G288) );
  XOR2_X1 U763 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n681) );
  XNOR2_X1 U764 ( .A(n731), .B(KEYINPUT87), .ZN(n680) );
  XNOR2_X1 U765 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U766 ( .A(n690), .B(n682), .ZN(n684) );
  XNOR2_X1 U767 ( .A(G290), .B(G305), .ZN(n683) );
  XNOR2_X1 U768 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U769 ( .A(G166), .B(n685), .ZN(n686) );
  XNOR2_X1 U770 ( .A(n686), .B(G288), .ZN(n884) );
  XNOR2_X1 U771 ( .A(n884), .B(n687), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n688), .A2(G868), .ZN(n692) );
  NAND2_X1 U773 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U774 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U775 ( .A(KEYINPUT88), .B(n693), .Z(G295) );
  NAND2_X1 U776 ( .A1(G2084), .A2(G2078), .ZN(n694) );
  XNOR2_X1 U777 ( .A(n694), .B(KEYINPUT89), .ZN(n695) );
  XNOR2_X1 U778 ( .A(n695), .B(KEYINPUT20), .ZN(n696) );
  NAND2_X1 U779 ( .A1(n696), .A2(G2090), .ZN(n697) );
  XNOR2_X1 U780 ( .A(KEYINPUT21), .B(n697), .ZN(n698) );
  NAND2_X1 U781 ( .A1(n698), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U782 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U783 ( .A1(G220), .A2(G219), .ZN(n699) );
  XOR2_X1 U784 ( .A(KEYINPUT22), .B(n699), .Z(n700) );
  NOR2_X1 U785 ( .A1(G218), .A2(n700), .ZN(n701) );
  XNOR2_X1 U786 ( .A(KEYINPUT90), .B(n701), .ZN(n702) );
  NAND2_X1 U787 ( .A1(n702), .A2(G96), .ZN(n858) );
  NAND2_X1 U788 ( .A1(G2106), .A2(n858), .ZN(n703) );
  XNOR2_X1 U789 ( .A(n703), .B(KEYINPUT91), .ZN(n708) );
  NOR2_X1 U790 ( .A1(G236), .A2(G238), .ZN(n704) );
  NAND2_X1 U791 ( .A1(G69), .A2(n704), .ZN(n705) );
  NOR2_X1 U792 ( .A1(G237), .A2(n705), .ZN(n857) );
  NOR2_X1 U793 ( .A1(n706), .A2(n857), .ZN(n707) );
  NOR2_X1 U794 ( .A1(n708), .A2(n707), .ZN(G319) );
  INV_X1 U795 ( .A(G319), .ZN(n932) );
  NAND2_X1 U796 ( .A1(G483), .A2(G661), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n932), .A2(n709), .ZN(n856) );
  NAND2_X1 U798 ( .A1(n856), .A2(G36), .ZN(G176) );
  INV_X1 U799 ( .A(G166), .ZN(G303) );
  INV_X1 U800 ( .A(G301), .ZN(G171) );
  INV_X1 U801 ( .A(n819), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n710), .A2(n820), .ZN(n711) );
  XNOR2_X2 U803 ( .A(n711), .B(KEYINPUT64), .ZN(n743) );
  NOR2_X1 U804 ( .A1(n526), .A2(n998), .ZN(n715) );
  INV_X1 U805 ( .A(G1996), .ZN(n963) );
  XOR2_X1 U806 ( .A(KEYINPUT66), .B(KEYINPUT26), .Z(n712) );
  XNOR2_X1 U807 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n721), .A2(n992), .ZN(n719) );
  NOR2_X1 U809 ( .A1(G2067), .A2(n757), .ZN(n717) );
  NOR2_X1 U810 ( .A1(G1348), .A2(n759), .ZN(n716) );
  NOR2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U813 ( .A(n720), .B(KEYINPUT100), .ZN(n723) );
  OR2_X1 U814 ( .A1(n992), .A2(n721), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n729) );
  XOR2_X1 U816 ( .A(KEYINPUT27), .B(KEYINPUT99), .Z(n725) );
  NAND2_X1 U817 ( .A1(G2072), .A2(n759), .ZN(n724) );
  XNOR2_X1 U818 ( .A(n725), .B(n724), .ZN(n727) );
  AND2_X1 U819 ( .A1(n757), .A2(G1956), .ZN(n726) );
  NOR2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n728) );
  NAND2_X1 U822 ( .A1(n729), .A2(n728), .ZN(n734) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U824 ( .A(n732), .B(KEYINPUT28), .Z(n733) );
  NAND2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n736) );
  XNOR2_X1 U826 ( .A(n736), .B(n735), .ZN(n742) );
  NOR2_X1 U827 ( .A1(G1961), .A2(n759), .ZN(n738) );
  XOR2_X1 U828 ( .A(G2078), .B(KEYINPUT25), .Z(n968) );
  NOR2_X1 U829 ( .A1(n757), .A2(n968), .ZN(n737) );
  NOR2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U831 ( .A(n739), .B(KEYINPUT97), .ZN(n751) );
  NAND2_X1 U832 ( .A1(G171), .A2(n751), .ZN(n740) );
  XNOR2_X1 U833 ( .A(n740), .B(KEYINPUT98), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n756) );
  NOR2_X1 U835 ( .A1(n743), .A2(G2084), .ZN(n773) );
  INV_X1 U836 ( .A(n773), .ZN(n744) );
  INV_X1 U837 ( .A(G8), .ZN(n758) );
  OR2_X1 U838 ( .A1(G1966), .A2(n758), .ZN(n745) );
  INV_X1 U839 ( .A(n772), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n522), .A2(n746), .ZN(n747) );
  XNOR2_X1 U841 ( .A(n747), .B(KEYINPUT101), .ZN(n749) );
  XNOR2_X1 U842 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U843 ( .A1(G168), .A2(n750), .ZN(n753) );
  NOR2_X1 U844 ( .A1(G171), .A2(n751), .ZN(n752) );
  XNOR2_X1 U845 ( .A(n754), .B(n525), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n770) );
  NAND2_X1 U847 ( .A1(n770), .A2(G286), .ZN(n767) );
  NOR2_X1 U848 ( .A1(n757), .A2(G2090), .ZN(n761) );
  OR2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n777) );
  NOR2_X1 U850 ( .A1(G1971), .A2(n777), .ZN(n760) );
  NOR2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U852 ( .A(n762), .B(KEYINPUT103), .ZN(n763) );
  NOR2_X1 U853 ( .A1(G166), .A2(n763), .ZN(n764) );
  XOR2_X1 U854 ( .A(KEYINPUT104), .B(n764), .Z(n765) );
  OR2_X1 U855 ( .A1(n758), .A2(n765), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n769) );
  INV_X1 U857 ( .A(KEYINPUT32), .ZN(n768) );
  XNOR2_X1 U858 ( .A(n769), .B(n768), .ZN(n790) );
  INV_X1 U859 ( .A(n770), .ZN(n771) );
  NAND2_X1 U860 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n791) );
  NAND2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n986) );
  AND2_X1 U863 ( .A1(n791), .A2(n986), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n790), .A2(n776), .ZN(n782) );
  INV_X1 U865 ( .A(n986), .ZN(n779) );
  NOR2_X1 U866 ( .A1(G1976), .A2(G288), .ZN(n787) );
  NOR2_X1 U867 ( .A1(G1971), .A2(G303), .ZN(n778) );
  NOR2_X1 U868 ( .A1(n787), .A2(n778), .ZN(n987) );
  OR2_X1 U869 ( .A1(n779), .A2(n987), .ZN(n780) );
  OR2_X1 U870 ( .A1(n777), .A2(n780), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(n783), .ZN(n785) );
  NOR2_X1 U873 ( .A1(KEYINPUT33), .A2(n785), .ZN(n786) );
  INV_X1 U874 ( .A(n786), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n787), .A2(KEYINPUT33), .ZN(n788) );
  XOR2_X1 U876 ( .A(G1981), .B(G305), .Z(n999) );
  NAND2_X1 U877 ( .A1(n789), .A2(n523), .ZN(n797) );
  NAND2_X1 U878 ( .A1(n790), .A2(n791), .ZN(n794) );
  NOR2_X1 U879 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n795), .A2(n777), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U884 ( .A1(G1981), .A2(G305), .ZN(n799) );
  XOR2_X1 U885 ( .A(n799), .B(KEYINPUT24), .Z(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n528), .ZN(n832) );
  NAND2_X1 U887 ( .A1(G119), .A2(n916), .ZN(n803) );
  NAND2_X1 U888 ( .A1(G95), .A2(n920), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U890 ( .A1(n917), .A2(G107), .ZN(n804) );
  XOR2_X1 U891 ( .A(KEYINPUT94), .B(n804), .Z(n805) );
  NOR2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U893 ( .A1(n636), .A2(G131), .ZN(n807) );
  NAND2_X1 U894 ( .A1(n808), .A2(n807), .ZN(n905) );
  NAND2_X1 U895 ( .A1(G1991), .A2(n905), .ZN(n818) );
  NAND2_X1 U896 ( .A1(G105), .A2(n920), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT38), .B(n809), .Z(n814) );
  NAND2_X1 U898 ( .A1(G129), .A2(n916), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G117), .A2(n917), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U901 ( .A(KEYINPUT95), .B(n812), .Z(n813) );
  NOR2_X1 U902 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U903 ( .A1(n636), .A2(G141), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n816), .A2(n815), .ZN(n909) );
  NAND2_X1 U905 ( .A1(G1996), .A2(n909), .ZN(n817) );
  NAND2_X1 U906 ( .A1(n818), .A2(n817), .ZN(n937) );
  NOR2_X1 U907 ( .A1(n820), .A2(n819), .ZN(n846) );
  NAND2_X1 U908 ( .A1(n937), .A2(n846), .ZN(n821) );
  XOR2_X1 U909 ( .A(KEYINPUT96), .B(n821), .Z(n837) );
  INV_X1 U910 ( .A(n837), .ZN(n831) );
  NAND2_X1 U911 ( .A1(G128), .A2(n916), .ZN(n823) );
  NAND2_X1 U912 ( .A1(G116), .A2(n917), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U914 ( .A(n824), .B(KEYINPUT35), .ZN(n829) );
  NAND2_X1 U915 ( .A1(G104), .A2(n920), .ZN(n826) );
  NAND2_X1 U916 ( .A1(G140), .A2(n636), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U918 ( .A(KEYINPUT34), .B(n827), .Z(n828) );
  NAND2_X1 U919 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U920 ( .A(n830), .B(KEYINPUT36), .Z(n913) );
  XNOR2_X1 U921 ( .A(G2067), .B(KEYINPUT37), .ZN(n842) );
  NOR2_X1 U922 ( .A1(n913), .A2(n842), .ZN(n938) );
  NAND2_X1 U923 ( .A1(n846), .A2(n938), .ZN(n840) );
  AND2_X1 U924 ( .A1(n832), .A2(n524), .ZN(n834) );
  XNOR2_X1 U925 ( .A(G1986), .B(G290), .ZN(n985) );
  NAND2_X1 U926 ( .A1(n985), .A2(n846), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n849) );
  NOR2_X1 U928 ( .A1(G1996), .A2(n909), .ZN(n940) );
  NOR2_X1 U929 ( .A1(G1986), .A2(G290), .ZN(n835) );
  NOR2_X1 U930 ( .A1(G1991), .A2(n905), .ZN(n947) );
  NOR2_X1 U931 ( .A1(n835), .A2(n947), .ZN(n836) );
  NOR2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U933 ( .A1(n940), .A2(n838), .ZN(n839) );
  XNOR2_X1 U934 ( .A(KEYINPUT39), .B(n839), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n844) );
  AND2_X1 U936 ( .A1(n913), .A2(n842), .ZN(n843) );
  XOR2_X1 U937 ( .A(KEYINPUT106), .B(n843), .Z(n954) );
  NAND2_X1 U938 ( .A1(n844), .A2(n954), .ZN(n845) );
  XOR2_X1 U939 ( .A(KEYINPUT107), .B(n845), .Z(n847) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U941 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U942 ( .A(n850), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U943 ( .A(G223), .ZN(n851) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n851), .ZN(G217) );
  NAND2_X1 U945 ( .A1(G15), .A2(G2), .ZN(n852) );
  XNOR2_X1 U946 ( .A(KEYINPUT109), .B(n852), .ZN(n853) );
  NAND2_X1 U947 ( .A1(n853), .A2(G661), .ZN(n854) );
  XNOR2_X1 U948 ( .A(KEYINPUT110), .B(n854), .ZN(G259) );
  NAND2_X1 U949 ( .A1(G3), .A2(G1), .ZN(n855) );
  NAND2_X1 U950 ( .A1(n856), .A2(n855), .ZN(G188) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  INV_X1 U953 ( .A(n857), .ZN(n859) );
  NOR2_X1 U954 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U955 ( .A(KEYINPUT111), .B(n860), .ZN(G261) );
  INV_X1 U956 ( .A(G261), .ZN(G325) );
  XOR2_X1 U957 ( .A(G2100), .B(G2096), .Z(n862) );
  XNOR2_X1 U958 ( .A(KEYINPUT42), .B(G2678), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U960 ( .A(KEYINPUT43), .B(G2072), .Z(n864) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2090), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U963 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U964 ( .A(G2084), .B(G2078), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(G227) );
  XOR2_X1 U966 ( .A(G1976), .B(G1971), .Z(n870) );
  XNOR2_X1 U967 ( .A(G1986), .B(G1956), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n880) );
  XOR2_X1 U969 ( .A(KEYINPUT112), .B(KEYINPUT41), .Z(n872) );
  XNOR2_X1 U970 ( .A(G1996), .B(KEYINPUT113), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U972 ( .A(G1961), .B(G1966), .Z(n874) );
  XNOR2_X1 U973 ( .A(G1991), .B(G1981), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U975 ( .A(n876), .B(n875), .Z(n878) );
  XNOR2_X1 U976 ( .A(KEYINPUT114), .B(G2474), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(G229) );
  XNOR2_X1 U979 ( .A(n998), .B(G286), .ZN(n883) );
  XNOR2_X1 U980 ( .A(G171), .B(n881), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U983 ( .A1(G37), .A2(n886), .ZN(G397) );
  NAND2_X1 U984 ( .A1(G124), .A2(n916), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(KEYINPUT44), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G136), .A2(n636), .ZN(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT115), .B(n888), .Z(n889) );
  NAND2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n545), .A2(G100), .ZN(n892) );
  NAND2_X1 U990 ( .A1(G112), .A2(n917), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n893) );
  NOR2_X1 U992 ( .A1(n894), .A2(n893), .ZN(G162) );
  XOR2_X1 U993 ( .A(KEYINPUT48), .B(KEYINPUT119), .Z(n903) );
  NAND2_X1 U994 ( .A1(G103), .A2(n920), .ZN(n896) );
  NAND2_X1 U995 ( .A1(G139), .A2(n636), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n901) );
  NAND2_X1 U997 ( .A1(G127), .A2(n916), .ZN(n898) );
  NAND2_X1 U998 ( .A1(G115), .A2(n917), .ZN(n897) );
  NAND2_X1 U999 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n899), .Z(n900) );
  NOR2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n950) );
  XNOR2_X1 U1002 ( .A(n950), .B(KEYINPUT118), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(KEYINPUT46), .B(n904), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n905), .B(KEYINPUT117), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(G164), .B(G160), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1010 ( .A(n912), .B(n943), .Z(n915) );
  XOR2_X1 U1011 ( .A(n913), .B(G162), .Z(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n928) );
  NAND2_X1 U1013 ( .A1(G130), .A2(n916), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(G118), .A2(n917), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n926) );
  NAND2_X1 U1016 ( .A1(n920), .A2(G106), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n921), .B(KEYINPUT116), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(G142), .A2(n636), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1020 ( .A(n924), .B(KEYINPUT45), .Z(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1022 ( .A(n928), .B(n927), .Z(n929) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n929), .ZN(G395) );
  NOR2_X1 U1024 ( .A1(G227), .A2(G229), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT49), .B(n930), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(G401), .A2(n931), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(G397), .A2(n932), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n935), .A2(G395), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(n936), .B(KEYINPUT120), .ZN(G308) );
  INV_X1 U1031 ( .A(G308), .ZN(G225) );
  INV_X1 U1032 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n949) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT51), .B(n941), .Z(n945) );
  XOR2_X1 U1037 ( .A(G2084), .B(G160), .Z(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n957) );
  XOR2_X1 U1042 ( .A(G2072), .B(n950), .Z(n952) );
  XOR2_X1 U1043 ( .A(G164), .B(G2078), .Z(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(KEYINPUT50), .B(n953), .ZN(n955) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1047 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1048 ( .A(KEYINPUT52), .B(n958), .Z(n959) );
  NOR2_X1 U1049 ( .A1(KEYINPUT55), .A2(n959), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(KEYINPUT121), .B(n960), .ZN(n961) );
  NAND2_X1 U1051 ( .A1(n961), .A2(G29), .ZN(n1039) );
  XOR2_X1 U1052 ( .A(G2067), .B(G26), .Z(n962) );
  NAND2_X1 U1053 ( .A1(n962), .A2(G28), .ZN(n967) );
  XNOR2_X1 U1054 ( .A(G32), .B(n963), .ZN(n965) );
  XOR2_X1 U1055 ( .A(G2072), .B(G33), .Z(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n972) );
  XNOR2_X1 U1058 ( .A(G1991), .B(G25), .ZN(n970) );
  XNOR2_X1 U1059 ( .A(G27), .B(n968), .ZN(n969) );
  NOR2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(KEYINPUT53), .B(n973), .ZN(n977) );
  XOR2_X1 U1063 ( .A(G34), .B(KEYINPUT122), .Z(n975) );
  XNOR2_X1 U1064 ( .A(G2084), .B(KEYINPUT54), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n975), .B(n974), .ZN(n976) );
  NAND2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(G35), .B(G2090), .ZN(n978) );
  NOR2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(KEYINPUT55), .B(n980), .ZN(n982) );
  INV_X1 U1070 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n983), .A2(G11), .ZN(n1037) );
  XNOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1074 ( .A(G1956), .B(G299), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n991) );
  AND2_X1 U1076 ( .A1(G303), .A2(G1971), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n996) );
  XNOR2_X1 U1080 ( .A(G171), .B(G1961), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(n992), .B(G1348), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(KEYINPUT124), .B(n997), .ZN(n1006) );
  XNOR2_X1 U1085 ( .A(n998), .B(G1341), .ZN(n1004) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G168), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1001), .B(KEYINPUT57), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT123), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1091 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1092 ( .A1(n1008), .A2(n1007), .ZN(n1035) );
  INV_X1 U1093 ( .A(G16), .ZN(n1033) );
  XOR2_X1 U1094 ( .A(G1981), .B(G6), .Z(n1011) );
  XNOR2_X1 U1095 ( .A(G20), .B(KEYINPUT125), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1009), .B(G1956), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G19), .B(G1341), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(KEYINPUT126), .B(n1014), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1348), .B(KEYINPUT59), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(n1015), .B(G4), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(n1018), .B(KEYINPUT60), .ZN(n1030) );
  XOR2_X1 U1105 ( .A(G1986), .B(G24), .Z(n1022) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(n1024), .B(n1023), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(G1966), .B(G21), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(G5), .B(G1961), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1121 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1040), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

