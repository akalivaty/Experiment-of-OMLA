//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n556, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(G2104), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR3_X1   g040(.A1(new_n465), .A2(KEYINPUT65), .A3(G2105), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(G137), .A3(new_n463), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT66), .ZN(G160));
  NAND2_X1  g054(.A1(new_n476), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT67), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n476), .A2(new_n482), .A3(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n476), .A2(new_n463), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(new_n491), .B2(G136), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n486), .A2(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(new_n463), .A2(G138), .ZN(new_n494));
  INV_X1    g069(.A(new_n472), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(new_n470), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT68), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n476), .A2(new_n498), .A3(new_n494), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(KEYINPUT4), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n496), .A2(KEYINPUT68), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n476), .A2(G126), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n500), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT69), .B1(new_n509), .B2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT6), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(new_n513), .B1(new_n509), .B2(G651), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(new_n512), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n510), .A2(new_n513), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n509), .A2(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n516), .A2(new_n523), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND3_X1  g105(.A1(new_n514), .A2(G51), .A3(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n533), .A2(new_n534), .B1(new_n521), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n531), .B(new_n536), .C1(new_n526), .C2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n519), .B2(new_n520), .ZN(new_n541));
  AND2_X1   g116(.A1(G77), .A2(G543), .ZN(new_n542));
  OAI21_X1  g117(.A(G651), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n524), .A2(G52), .A3(G543), .A4(new_n525), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n524), .A2(new_n521), .A3(G90), .A4(new_n525), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(new_n515), .A2(G43), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n512), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n527), .A2(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g130(.A(KEYINPUT71), .B(KEYINPUT8), .Z(new_n556));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n525), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n514), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n524), .A2(new_n521), .A3(G91), .A4(new_n525), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n564), .B(new_n565), .C1(new_n512), .C2(new_n566), .ZN(G299));
  NAND3_X1  g142(.A1(new_n514), .A2(G49), .A3(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n568), .B(new_n569), .C1(new_n526), .C2(new_n570), .ZN(G288));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n519), .B2(new_n520), .ZN(new_n573));
  AND2_X1   g148(.A1(G73), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n524), .A2(new_n521), .A3(G86), .A4(new_n525), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n524), .A2(G48), .A3(G543), .A4(new_n525), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(new_n515), .A2(G47), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n512), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n527), .A2(G85), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n526), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n514), .A2(KEYINPUT10), .A3(G92), .A4(new_n521), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n519), .B2(new_n520), .ZN(new_n591));
  AND2_X1   g166(.A1(G79), .A2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT72), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n524), .A2(G54), .A3(G543), .A4(new_n525), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n589), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n584), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n584), .B1(new_n599), .B2(G868), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n565), .B1(new_n566), .B2(new_n512), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n561), .B2(new_n563), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n602), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n599), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n599), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n467), .A2(new_n476), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT73), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT13), .Z(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n491), .A2(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n463), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n620), .B1(new_n621), .B2(new_n622), .C1(new_n484), .C2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n618), .A2(new_n619), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT76), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT77), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT77), .ZN(new_n638));
  NAND4_X1  g213(.A1(new_n634), .A2(new_n638), .A3(KEYINPUT14), .A4(new_n635), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n629), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n637), .A2(new_n639), .A3(new_n629), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT75), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n637), .A2(new_n639), .A3(new_n629), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(new_n640), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT78), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n655));
  NAND4_X1  g230(.A1(new_n647), .A2(new_n650), .A3(new_n655), .A4(new_n652), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n647), .A2(new_n650), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(new_n659), .B2(new_n651), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  INV_X1    g237(.A(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n617), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n625), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  INV_X1    g266(.A(new_n689), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n686), .A2(new_n687), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n690), .A2(new_n694), .A3(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(G160), .A2(G29), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT79), .B(G29), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT24), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G34), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n704), .A2(KEYINPUT85), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT85), .B1(new_n704), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(G34), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n702), .A2(G2084), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT86), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G33), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G139), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n490), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n476), .A2(G127), .ZN(new_n720));
  NAND2_X1  g295(.A1(G115), .A2(G2104), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n463), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n714), .B1(new_n723), .B2(new_n713), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT84), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2072), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT27), .B(G1996), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT88), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n713), .A2(G32), .ZN(new_n729));
  INV_X1    g304(.A(G129), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n484), .A2(KEYINPUT87), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(KEYINPUT87), .B1(new_n484), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT26), .Z(new_n735));
  INV_X1    g310(.A(G141), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n490), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G105), .B2(new_n467), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n729), .B1(new_n740), .B2(new_n713), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n712), .B(new_n726), .C1(new_n728), .C2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT89), .Z(new_n743));
  NOR2_X1   g318(.A1(new_n704), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n704), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT29), .Z(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n741), .A2(new_n728), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n704), .A2(G27), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n704), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT91), .B(G2078), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G16), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G19), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n553), .B2(new_n755), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n754), .B1(G1341), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(G1341), .ZN(new_n760));
  AOI21_X1  g335(.A(G2084), .B1(new_n702), .B2(new_n710), .ZN(new_n761));
  INV_X1    g336(.A(G1961), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n755), .A2(G5), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G301), .B2(G16), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n760), .B(new_n761), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n755), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1956), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(G28), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n713), .B1(new_n772), .B2(G28), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n771), .B1(new_n773), .B2(new_n774), .C1(new_n624), .C2(new_n703), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n755), .A2(G21), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G168), .B2(new_n755), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n777), .A2(G1966), .B1(new_n764), .B2(new_n762), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n775), .B(new_n778), .C1(G1966), .C2(new_n777), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n759), .A2(new_n770), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n703), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT28), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n481), .A2(G128), .A3(new_n483), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT81), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT82), .Z(new_n789));
  INV_X1    g364(.A(G116), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n465), .B1(new_n790), .B2(G2105), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n791), .B1(new_n491), .B2(G140), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n784), .B1(new_n794), .B2(new_n713), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT83), .B(G2067), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n599), .A2(new_n755), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G4), .B2(new_n755), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1348), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n743), .A2(new_n782), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n755), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n755), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n755), .A2(G23), .ZN(new_n809));
  INV_X1    g384(.A(G288), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n755), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT33), .B(G1976), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n805), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT34), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n755), .A2(G24), .ZN(new_n816));
  INV_X1    g391(.A(G290), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n755), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT80), .B(G1986), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n485), .A2(G119), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(G107), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G2105), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n491), .B2(G131), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  MUX2_X1   g401(.A(G25), .B(new_n826), .S(new_n704), .Z(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n815), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n801), .B1(new_n831), .B2(new_n832), .ZN(G311));
  XNOR2_X1  g408(.A(new_n830), .B(KEYINPUT36), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n782), .A2(new_n797), .A3(new_n800), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n743), .A3(new_n835), .ZN(G150));
  AOI22_X1  g411(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n512), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n524), .A2(new_n521), .A3(G93), .A4(new_n525), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n524), .A2(G55), .A3(G543), .A4(new_n525), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT92), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n839), .B2(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT93), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(new_n838), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n552), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n844), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n849), .A2(new_n846), .A3(new_n553), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n599), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n844), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XOR2_X1   g435(.A(KEYINPUT95), .B(G37), .Z(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G160), .B(new_n624), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(G162), .Z(new_n864));
  NAND3_X1  g439(.A1(new_n787), .A2(G164), .A3(new_n792), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(G164), .B1(new_n787), .B2(new_n792), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n740), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n739), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n723), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n870), .A3(new_n723), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n826), .B(new_n615), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n491), .A2(G142), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT94), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n485), .A2(G130), .ZN(new_n879));
  OR2_X1    g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n876), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n864), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n873), .A2(new_n874), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n862), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n875), .B1(new_n888), .B2(new_n885), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n873), .A2(KEYINPUT96), .A3(new_n874), .A4(new_n883), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n864), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT40), .B1(new_n887), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G395));
  OAI21_X1  g469(.A(KEYINPUT99), .B1(new_n849), .B2(G868), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n896));
  XNOR2_X1  g471(.A(G303), .B(G288), .ZN(new_n897));
  XNOR2_X1  g472(.A(G290), .B(G305), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n897), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n900), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(KEYINPUT97), .A3(KEYINPUT42), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n906), .A3(new_n902), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT98), .B1(new_n904), .B2(KEYINPUT42), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n903), .A2(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n851), .B(new_n609), .ZN(new_n910));
  NAND2_X1  g485(.A1(G299), .A2(new_n598), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n593), .A2(new_n595), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT72), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n604), .A3(new_n589), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n911), .A2(new_n916), .A3(KEYINPUT41), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n911), .B2(new_n916), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n910), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n909), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G868), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(new_n909), .B2(new_n922), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n895), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT99), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n923), .A2(new_n925), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G295));
  AOI21_X1  g504(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  NAND2_X1  g506(.A1(G301), .A2(KEYINPUT100), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n932), .A2(G286), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G286), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n851), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n848), .A2(new_n937), .A3(new_n850), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n921), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n917), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n848), .A2(new_n937), .A3(new_n850), .ZN(new_n943));
  INV_X1    g518(.A(new_n936), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n932), .A2(G286), .A3(new_n934), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n848), .A2(new_n850), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n942), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n901), .ZN(new_n949));
  INV_X1    g524(.A(G37), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n941), .A2(new_n947), .A3(new_n904), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n949), .A2(KEYINPUT43), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n941), .A2(new_n947), .A3(new_n904), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n904), .B1(new_n941), .B2(new_n947), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(new_n954), .A3(new_n862), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n931), .B(new_n952), .C1(new_n955), .C2(KEYINPUT43), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT101), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n949), .A2(new_n861), .A3(new_n951), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(KEYINPUT101), .A3(new_n931), .A4(new_n952), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n949), .A2(new_n960), .A3(new_n950), .A4(new_n951), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n964), .A2(KEYINPUT102), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(KEYINPUT102), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n931), .B1(new_n959), .B2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(G397));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT45), .B1(new_n507), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT103), .B(G40), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n468), .A2(new_n475), .A3(new_n477), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n828), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n826), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n821), .A2(new_n828), .A3(new_n825), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n497), .A2(KEYINPUT4), .A3(new_n499), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n502), .A2(new_n505), .A3(new_n503), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n970), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(new_n973), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(G1996), .A3(new_n739), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT105), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT104), .B1(new_n975), .B2(G1996), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n740), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n793), .A2(G2067), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n793), .A2(G2067), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n985), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n987), .A2(new_n993), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(G290), .B(G1986), .ZN(new_n999));
  AOI211_X1 g574(.A(new_n979), .B(new_n998), .C1(new_n985), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2078), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n983), .A2(G1384), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n973), .B1(new_n507), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n984), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n1007));
  NOR2_X1   g582(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n973), .B1(new_n507), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n762), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1005), .A2(G2078), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n984), .A2(new_n1003), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1006), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G171), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1004), .A2(new_n1005), .B1(new_n1010), .B2(new_n762), .ZN(new_n1016));
  OR3_X1    g591(.A1(new_n473), .A2(KEYINPUT122), .A3(new_n474), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT122), .B1(new_n473), .B2(new_n474), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(G2105), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n468), .A2(KEYINPUT121), .A3(new_n477), .ZN(new_n1020));
  INV_X1    g595(.A(G40), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n464), .A2(new_n466), .ZN(new_n1022));
  INV_X1    g597(.A(G101), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n477), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT121), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1019), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(new_n984), .A3(KEYINPUT123), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT123), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n971), .B2(new_n1027), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n507), .A2(new_n1002), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .A4(new_n1012), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1016), .A2(new_n1033), .A3(G301), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT54), .B1(new_n1015), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1966), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n974), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(new_n1037), .B2(new_n971), .ZN(new_n1038));
  INV_X1    g613(.A(G2084), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1007), .A2(new_n1039), .A3(new_n1009), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT108), .B(G8), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G286), .A2(new_n1043), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(KEYINPUT51), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1045), .B(KEYINPUT120), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT51), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1045), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT119), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1035), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1007), .A2(new_n747), .A3(new_n1009), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT106), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT106), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1007), .A2(new_n1060), .A3(new_n1009), .A4(new_n747), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n804), .B1(new_n1037), .B2(new_n971), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT107), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(G166), .B2(new_n1049), .ZN(new_n1066));
  NAND3_X1  g641(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT107), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1059), .A2(new_n1069), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1064), .A2(G8), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1062), .A2(new_n1058), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1068), .B1(new_n1072), .B2(new_n1043), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n502), .A2(new_n505), .A3(new_n503), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1384), .B1(new_n1074), .B2(new_n500), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1042), .B1(new_n1075), .B2(new_n974), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n527), .A2(G87), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(new_n568), .A3(new_n569), .A4(G1976), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1043), .B(new_n1079), .C1(new_n982), .C2(new_n973), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT109), .B1(new_n1083), .B2(KEYINPUT52), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n974), .A2(new_n970), .A3(new_n507), .ZN(new_n1085));
  AND4_X1   g660(.A1(new_n1085), .A2(new_n1043), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1981), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT110), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(KEYINPUT111), .A2(G86), .ZN(new_n1092));
  AND2_X1   g667(.A1(KEYINPUT111), .A2(G86), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n526), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n575), .A2(new_n577), .ZN(new_n1095));
  OAI21_X1  g670(.A(G1981), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(KEYINPUT112), .A2(KEYINPUT49), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1091), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1076), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1073), .A2(new_n1087), .A3(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1071), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1016), .A2(new_n1033), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(G171), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1014), .A2(G171), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(KEYINPUT124), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1014), .A2(new_n1109), .A3(G171), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1106), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1057), .A2(new_n1103), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n564), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G299), .B(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT113), .B(G1956), .Z(new_n1117));
  NAND2_X1  g692(.A1(new_n1010), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n984), .A2(new_n1003), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1116), .B1(new_n1120), .B2(new_n1118), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1113), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1116), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT61), .A3(new_n1121), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n984), .A2(new_n989), .A3(new_n1003), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT58), .B(G1341), .Z(new_n1130));
  NAND3_X1  g705(.A1(new_n1085), .A2(KEYINPUT115), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT115), .B1(new_n1085), .B2(new_n1130), .ZN(new_n1133));
  OAI211_X1 g708(.A(KEYINPUT117), .B(new_n553), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT116), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1124), .A2(new_n1128), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n553), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1139), .B(KEYINPUT59), .C1(new_n1135), .C2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1348), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1010), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G2067), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1075), .A2(new_n1144), .A3(new_n974), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(KEYINPUT60), .A3(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(KEYINPUT118), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(KEYINPUT118), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n599), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(KEYINPUT118), .A3(new_n598), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT60), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1138), .B(new_n1141), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n598), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1121), .B1(new_n1123), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1112), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1044), .A2(G286), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1071), .A2(new_n1102), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1064), .A2(G8), .A3(new_n1070), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1068), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1041), .A2(KEYINPUT63), .A3(G168), .A4(new_n1043), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1164), .A2(new_n1087), .A3(new_n1101), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1071), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1007), .A2(new_n1039), .A3(new_n1009), .ZN(new_n1168));
  AOI21_X1  g743(.A(G1966), .B1(new_n984), .B2(new_n1003), .ZN(new_n1169));
  OAI21_X1  g744(.A(G8), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1051), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1171), .A2(KEYINPUT51), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1055), .A2(KEYINPUT119), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT119), .ZN(new_n1174));
  AOI211_X1 g749(.A(new_n1174), .B(new_n1045), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT62), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1015), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1054), .A2(new_n1056), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1103), .A2(new_n1177), .A3(new_n1178), .A4(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1071), .A2(new_n1101), .A3(new_n1087), .ZN(new_n1182));
  OR3_X1    g757(.A1(new_n1101), .A2(G1976), .A3(G288), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1100), .B1(new_n1183), .B2(new_n1091), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1167), .A2(new_n1181), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1000), .B1(new_n1156), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n996), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n998), .B2(new_n978), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n998), .A2(new_n979), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n975), .A2(G1986), .A3(G290), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT48), .Z(new_n1192));
  AOI22_X1  g767(.A1(new_n1189), .A2(new_n985), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT46), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n990), .A2(new_n1194), .A3(new_n991), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1195), .B(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1188), .A2(new_n740), .A3(new_n994), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1198), .A2(new_n985), .B1(new_n992), .B2(KEYINPUT46), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1197), .A2(KEYINPUT126), .A3(new_n1199), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1202), .A2(KEYINPUT47), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1193), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(KEYINPUT47), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1187), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g783(.A1(G227), .A2(new_n460), .ZN(new_n1210));
  XNOR2_X1  g784(.A(new_n1210), .B(KEYINPUT127), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n661), .A2(new_n700), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n887), .B2(new_n891), .ZN(new_n1213));
  AND3_X1   g787(.A1(new_n1213), .A2(new_n961), .A3(new_n952), .ZN(G308));
  NAND3_X1  g788(.A1(new_n1213), .A2(new_n961), .A3(new_n952), .ZN(G225));
endmodule


