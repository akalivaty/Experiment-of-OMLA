//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1188, new_n1189,
    new_n1190, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1240, new_n1241;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G107), .A2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n207), .B(new_n208), .C1(new_n201), .C2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n202), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NOR2_X1   g0023(.A1(G58), .A2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n220), .A2(new_n223), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G264), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n217), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  NOR2_X1   g0038(.A1(new_n201), .A2(new_n202), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(new_n203), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(KEYINPUT64), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT65), .B(G107), .ZN(new_n245));
  INV_X1    g0045(.A(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n244), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n253), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT66), .B(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n259), .A2(new_n213), .B1(new_n217), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n261), .A2(new_n262), .B1(G33), .B2(G97), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n255), .B1(new_n209), .B2(new_n258), .C1(new_n263), .C2(new_n257), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(KEYINPUT13), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(KEYINPUT13), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G190), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n228), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n227), .A2(G33), .ZN(new_n272));
  OAI22_X1  g0072(.A1(new_n272), .A2(new_n202), .B1(new_n227), .B2(G68), .ZN(new_n273));
  XOR2_X1   g0073(.A(new_n273), .B(KEYINPUT70), .Z(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n212), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n271), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(new_n278), .B(KEYINPUT11), .Z(new_n279));
  NAND3_X1  g0079(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n252), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n201), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT12), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(new_n271), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n287), .B(new_n288), .C1(G1), .C2(new_n227), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n201), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n267), .A2(G200), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n269), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n265), .A2(G179), .A3(new_n266), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT71), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT14), .B1(new_n268), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT14), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n267), .A2(new_n299), .A3(G169), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n291), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n294), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n262), .B1(new_n209), .B2(new_n260), .C1(new_n259), .C2(new_n217), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n256), .C1(G107), .C2(new_n262), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n257), .A2(G244), .A3(new_n253), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n255), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(G179), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n297), .B2(new_n307), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G20), .A2(G77), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT8), .B(G58), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n310), .B1(new_n311), .B2(new_n272), .C1(new_n276), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n271), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n284), .A2(new_n202), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n314), .B(new_n315), .C1(new_n202), .C2(new_n289), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n303), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(G20), .B1(new_n225), .B2(G50), .ZN(new_n319));
  INV_X1    g0119(.A(G150), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n216), .A2(KEYINPUT8), .ZN(new_n321));
  MUX2_X1   g0121(.A(new_n312), .B(new_n321), .S(KEYINPUT67), .Z(new_n322));
  OAI221_X1 g0122(.A(new_n319), .B1(new_n320), .B2(new_n276), .C1(new_n322), .C2(new_n272), .ZN(new_n323));
  INV_X1    g0123(.A(new_n289), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n323), .A2(new_n271), .B1(G50), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G50), .B2(new_n287), .ZN(new_n326));
  INV_X1    g0126(.A(G223), .ZN(new_n327));
  INV_X1    g0127(.A(G222), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n262), .B1(new_n327), .B2(new_n260), .C1(new_n259), .C2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(new_n256), .C1(G77), .C2(new_n262), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(new_n255), .C1(new_n213), .C2(new_n258), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n297), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n326), .B(new_n332), .C1(G179), .C2(new_n331), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(G200), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT9), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n335), .B1(new_n336), .B2(new_n331), .C1(new_n326), .C2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n326), .A2(new_n337), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n338), .A2(KEYINPUT10), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT10), .B1(new_n338), .B2(new_n339), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n334), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT3), .ZN(new_n344));
  INV_X1    g0144(.A(G33), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n227), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n346), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n347), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n201), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G159), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n276), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G58), .A2(G68), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n227), .B1(new_n225), .B2(new_n355), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n343), .B1(new_n357), .B2(KEYINPUT16), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n288), .B1(new_n357), .B2(KEYINPUT16), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n227), .ZN(new_n364));
  INV_X1    g0164(.A(new_n351), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n356), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(KEYINPUT72), .B(new_n360), .C1(new_n368), .C2(new_n354), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n358), .A2(new_n359), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n322), .A2(new_n287), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n324), .B2(new_n322), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n257), .A2(G232), .A3(new_n253), .ZN(new_n374));
  INV_X1    g0174(.A(G87), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n345), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G226), .A2(G1698), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n259), .B2(new_n327), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n378), .B2(new_n262), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n255), .B(new_n374), .C1(new_n379), .C2(new_n257), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G169), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n260), .A2(KEYINPUT66), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT66), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G223), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n363), .B1(new_n386), .B2(new_n377), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n256), .B1(new_n387), .B2(new_n376), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n388), .A2(G179), .A3(new_n255), .A4(new_n374), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT73), .B1(new_n381), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n381), .A2(KEYINPUT73), .A3(new_n389), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n373), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n380), .A2(G200), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n380), .A2(new_n336), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n370), .A2(new_n395), .A3(new_n396), .A4(new_n372), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(new_n398), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT74), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n370), .A2(new_n396), .A3(new_n372), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT17), .A3(new_n395), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(new_n398), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT74), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n394), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n307), .A2(new_n336), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n307), .A2(G200), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n409), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  AND4_X1   g0213(.A1(new_n318), .A2(new_n342), .A3(new_n408), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G264), .A2(G1698), .ZN(new_n415));
  INV_X1    g0215(.A(G257), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n262), .B(new_n415), .C1(new_n259), .C2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G303), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n363), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT81), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT81), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(new_n422), .A3(new_n419), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n256), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT5), .B(G41), .ZN(new_n425));
  INV_X1    g0225(.A(G45), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(G1), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(G274), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n425), .A2(new_n430), .A3(G274), .A4(new_n427), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n256), .B1(new_n425), .B2(new_n427), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n429), .A2(new_n431), .B1(new_n432), .B2(G270), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n287), .A2(G116), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT20), .ZN(new_n436));
  INV_X1    g0236(.A(G97), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n227), .B1(new_n437), .B2(G33), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT75), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(G33), .A3(G283), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G283), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT75), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n438), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n270), .A2(new_n228), .B1(G20), .B2(new_n246), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n436), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(new_n440), .ZN(new_n447));
  INV_X1    g0247(.A(new_n438), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n444), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n435), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n252), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n287), .A2(new_n288), .A3(G116), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n297), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT21), .B1(new_n434), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n446), .A2(new_n450), .ZN(new_n456));
  INV_X1    g0256(.A(new_n435), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(new_n453), .ZN(new_n458));
  AND4_X1   g0258(.A1(G179), .A2(new_n458), .A3(new_n424), .A4(new_n433), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n434), .A2(KEYINPUT21), .A3(new_n454), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT82), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n434), .A2(new_n454), .A3(KEYINPUT82), .A4(KEYINPUT21), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n434), .A2(G200), .ZN(new_n465));
  INV_X1    g0265(.A(new_n458), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n424), .A2(new_n433), .A3(G190), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n460), .A2(new_n463), .A3(new_n464), .A4(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  OAI21_X1  g0271(.A(G244), .B1(new_n361), .B2(new_n362), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(new_n259), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n385), .A2(new_n262), .A3(KEYINPUT4), .A4(G244), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n262), .A2(G250), .A3(G1698), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n447), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n256), .ZN(new_n477));
  INV_X1    g0277(.A(G179), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n429), .A2(new_n431), .B1(new_n432), .B2(G257), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT77), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n477), .A2(new_n479), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n297), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n287), .A2(new_n288), .A3(new_n452), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n437), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n284), .A2(new_n437), .ZN(new_n487));
  INV_X1    g0287(.A(G107), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n350), .B2(new_n351), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT6), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n437), .A2(new_n488), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n488), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n227), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n276), .A2(new_n202), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n486), .B(new_n487), .C1(new_n497), .C2(new_n288), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT77), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n477), .A2(new_n499), .A3(new_n478), .A4(new_n479), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n481), .A2(new_n483), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n482), .A2(G200), .ZN(new_n502));
  OAI21_X1  g0302(.A(G107), .B1(new_n364), .B2(new_n365), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n493), .A2(new_n494), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G20), .ZN(new_n505));
  INV_X1    g0305(.A(new_n496), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n485), .B1(new_n507), .B2(new_n271), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n477), .A2(G190), .A3(new_n479), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n502), .A2(new_n487), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n257), .B1(G250), .B2(new_n427), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n426), .A2(G1), .A3(G274), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n209), .B1(new_n382), .B2(new_n384), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT78), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n262), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n472), .A2(new_n260), .B1(new_n345), .B2(new_n246), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n516), .B1(new_n515), .B2(new_n262), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n478), .B(new_n514), .C1(new_n521), .C2(new_n257), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n272), .B2(new_n437), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT79), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n262), .A2(new_n227), .A3(G68), .ZN(new_n526));
  NAND3_X1  g0326(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n227), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n375), .A2(new_n437), .A3(new_n488), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT79), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n523), .C1(new_n272), .C2(new_n437), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n525), .A2(new_n526), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n271), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n284), .A2(new_n311), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n535), .C1(new_n311), .C2(new_n484), .ZN(new_n536));
  INV_X1    g0336(.A(new_n520), .ZN(new_n537));
  INV_X1    g0337(.A(new_n519), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(new_n517), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n513), .B1(new_n539), .B2(new_n256), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n522), .B(new_n536), .C1(G169), .C2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G190), .B(new_n514), .C1(new_n521), .C2(new_n257), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n287), .A2(new_n288), .A3(G87), .A4(new_n452), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n534), .A2(new_n535), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G200), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n542), .B(new_n544), .C1(new_n545), .C2(new_n540), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n501), .A2(new_n510), .A3(new_n541), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n469), .B1(new_n470), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT23), .A2(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(G20), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n227), .A2(KEYINPUT23), .A3(G107), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n552), .A2(KEYINPUT83), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(KEYINPUT83), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n363), .A2(G20), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(G87), .ZN(new_n558));
  NOR4_X1   g0358(.A1(new_n363), .A2(KEYINPUT22), .A3(G20), .A4(new_n375), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n555), .B(KEYINPUT24), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n271), .A3(new_n563), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n484), .A2(new_n488), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n287), .A2(G107), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT25), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n432), .A2(G264), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT84), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT84), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n432), .A2(new_n571), .A3(G264), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n429), .A2(new_n431), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n385), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n575));
  INV_X1    g0375(.A(G294), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n575), .A2(new_n363), .B1(new_n345), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n256), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n545), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n573), .A2(new_n336), .A3(new_n574), .A4(new_n578), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(KEYINPUT85), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n568), .B(new_n582), .C1(KEYINPUT85), .C2(new_n581), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n297), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(G179), .B2(new_n579), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n568), .ZN(new_n586));
  AND4_X1   g0386(.A1(new_n501), .A2(new_n510), .A3(new_n541), .A4(new_n546), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(KEYINPUT80), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n414), .A2(new_n548), .A3(new_n583), .A4(new_n588), .ZN(G372));
  NAND2_X1  g0389(.A1(new_n434), .A2(new_n454), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n458), .A2(new_n424), .A3(G179), .A4(new_n433), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n463), .A2(new_n592), .A3(new_n593), .A4(new_n464), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT86), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n460), .A2(new_n596), .A3(new_n463), .A4(new_n464), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n586), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT87), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n587), .A2(new_n583), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n586), .B1(new_n595), .B2(new_n597), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT87), .B1(new_n605), .B2(new_n602), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT88), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n501), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n508), .A2(new_n487), .B1(new_n482), .B2(new_n297), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n609), .A2(KEYINPUT88), .A3(new_n481), .A4(new_n500), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n541), .A2(new_n546), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(KEYINPUT89), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n612), .A2(new_n501), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT26), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT89), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n612), .B1(new_n608), .B2(new_n610), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(KEYINPUT26), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n616), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n604), .A2(new_n606), .A3(new_n541), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n414), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n381), .A2(new_n389), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n373), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(new_n393), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n401), .B1(new_n399), .B2(new_n400), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n404), .A2(KEYINPUT74), .A3(new_n405), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n293), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n318), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n340), .A2(new_n341), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n334), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n624), .A2(new_n634), .ZN(G369));
  INV_X1    g0435(.A(KEYINPUT91), .ZN(new_n636));
  INV_X1    g0436(.A(G13), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(G20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n252), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n466), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n595), .B2(new_n597), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n469), .A2(new_n647), .ZN(new_n649));
  OR3_X1    g0449(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT90), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT90), .B1(new_n648), .B2(new_n649), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G330), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n636), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n650), .A2(KEYINPUT91), .A3(G330), .A4(new_n651), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n599), .A2(new_n644), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n568), .A2(new_n645), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n583), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n586), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n660), .A2(new_n594), .A3(new_n599), .A4(new_n645), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n658), .A3(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n221), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G1), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n529), .A2(G116), .ZN(new_n670));
  OAI22_X1  g0470(.A1(new_n669), .A2(new_n670), .B1(new_n226), .B2(new_n668), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n672));
  XNOR2_X1  g0472(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n623), .A2(new_n645), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n617), .A2(new_n615), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n541), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(KEYINPUT26), .B2(new_n614), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n603), .B1(new_n594), .B2(new_n586), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n644), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT29), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT31), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n548), .A2(new_n583), .A3(new_n588), .A4(new_n645), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n434), .A2(new_n478), .ZN(new_n686));
  INV_X1    g0486(.A(new_n482), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n573), .A2(new_n578), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n540), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT30), .ZN(new_n690));
  AOI21_X1  g0490(.A(G179), .B1(new_n424), .B2(new_n433), .ZN(new_n691));
  INV_X1    g0491(.A(new_n540), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n482), .A4(new_n579), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n644), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n684), .B1(new_n685), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT31), .B1(new_n694), .B2(new_n644), .ZN(new_n697));
  OAI21_X1  g0497(.A(G330), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n683), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n673), .B1(new_n700), .B2(G1), .ZN(G364));
  AOI21_X1  g0501(.A(new_n228), .B1(G20), .B2(new_n297), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n336), .A2(new_n545), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n227), .A2(G179), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT96), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT96), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n227), .A2(new_n478), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n545), .A2(G190), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n709), .A2(new_n375), .B1(new_n201), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n336), .A2(G200), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n227), .B1(new_n714), .B2(new_n478), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT97), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(KEYINPUT97), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n437), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G190), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n705), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G159), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n713), .B(new_n720), .C1(KEYINPUT32), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n710), .A2(new_n714), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n710), .A2(new_n704), .ZN(new_n727));
  OAI221_X1 g0527(.A(new_n262), .B1(new_n726), .B2(new_n216), .C1(new_n212), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n710), .A2(new_n721), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(G77), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n705), .A2(new_n711), .ZN(new_n733));
  OAI221_X1 g0533(.A(new_n732), .B1(KEYINPUT32), .B2(new_n724), .C1(new_n488), .C2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G283), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n715), .A2(new_n576), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n712), .ZN(new_n737));
  XNOR2_X1  g0537(.A(KEYINPUT33), .B(G317), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n737), .A2(new_n738), .B1(new_n730), .B2(G311), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n723), .A2(G329), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(new_n363), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n727), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n736), .B(new_n741), .C1(G326), .C2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n743), .B1(new_n418), .B2(new_n709), .C1(new_n744), .C2(new_n726), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n703), .B1(new_n734), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n652), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n669), .B1(G45), .B2(new_n638), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n702), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n225), .A2(new_n426), .A3(G50), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n363), .A2(new_n221), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT95), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n754), .B(new_n756), .C1(new_n244), .C2(new_n426), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n666), .A2(new_n363), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n246), .B2(new_n666), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT94), .Z(new_n760));
  NAND2_X1  g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n746), .B(new_n752), .C1(new_n753), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n656), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n652), .A2(KEYINPUT93), .A3(new_n653), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT93), .B1(new_n652), .B2(new_n653), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n764), .A2(new_n765), .A3(new_n751), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n762), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(G396));
  NOR2_X1   g0568(.A1(new_n317), .A2(new_n644), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n316), .A2(new_n644), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n413), .A2(new_n770), .B1(new_n309), .B2(new_n316), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n769), .A2(new_n771), .A3(KEYINPUT100), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT100), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n623), .A2(new_n645), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n699), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n775), .A2(KEYINPUT101), .A3(new_n698), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n774), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(new_n674), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n751), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n674), .A2(new_n780), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n777), .A2(new_n783), .A3(new_n778), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n747), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n702), .A2(new_n747), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT98), .Z(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n202), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n733), .A2(new_n201), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n726), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G143), .A2(new_n792), .B1(new_n737), .B2(G150), .ZN(new_n793));
  INV_X1    g0593(.A(G137), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n794), .B2(new_n727), .C1(new_n353), .C2(new_n729), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n791), .B1(new_n796), .B2(KEYINPUT34), .ZN(new_n797));
  INV_X1    g0597(.A(new_n715), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(G58), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n363), .B1(new_n796), .B2(KEYINPUT34), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(new_n212), .C2(new_n709), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G132), .B2(new_n723), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n709), .A2(new_n488), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n803), .B(new_n720), .C1(G311), .C2(new_n723), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT99), .B(G283), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n363), .B1(new_n733), .B2(new_n375), .C1(new_n806), .C2(new_n712), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G294), .B2(new_n792), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n804), .B(new_n808), .C1(new_n246), .C2(new_n729), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G303), .B2(new_n742), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n702), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n786), .A2(new_n751), .A3(new_n789), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n785), .A2(new_n812), .ZN(G384));
  XNOR2_X1  g0613(.A(new_n769), .B(KEYINPUT103), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n775), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n302), .A2(new_n644), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n303), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n301), .A2(new_n302), .A3(new_n644), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n642), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n359), .B1(KEYINPUT16), .B2(new_n357), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n372), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n407), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n373), .A2(new_n822), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n826), .A2(new_n397), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT104), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n392), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n392), .A2(new_n826), .A3(new_n829), .A4(new_n397), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT104), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n824), .B1(new_n625), .B2(new_n822), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n834), .A2(new_n397), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n833), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n825), .A2(new_n836), .A3(KEYINPUT38), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT38), .B1(new_n825), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n821), .A2(new_n839), .B1(new_n627), .B2(new_n822), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n835), .A2(new_n829), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n830), .B2(new_n832), .ZN(new_n843));
  INV_X1    g0643(.A(new_n824), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n630), .B2(new_n394), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(new_n822), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n827), .A2(new_n626), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n830), .A2(new_n832), .B1(new_n848), .B2(KEYINPUT37), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n399), .A2(new_n400), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n826), .B1(new_n627), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n846), .A2(KEYINPUT38), .B1(new_n852), .B2(KEYINPUT105), .ZN(new_n853));
  AND4_X1   g0653(.A1(KEYINPUT105), .A2(new_n825), .A3(KEYINPUT38), .A4(new_n836), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n841), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n301), .A2(new_n302), .A3(new_n645), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n840), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n414), .A2(new_n676), .A3(new_n682), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n634), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n861), .B(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n820), .B(new_n774), .C1(new_n696), .C2(new_n697), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n866), .B(KEYINPUT40), .C1(new_n853), .C2(new_n854), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT40), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n839), .B2(new_n865), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n869), .A3(G330), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n414), .A2(new_n699), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n696), .A2(new_n697), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n867), .A2(new_n414), .A3(new_n873), .A4(new_n869), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n864), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n252), .B2(new_n638), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n246), .B1(new_n504), .B2(KEYINPUT35), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n228), .A2(new_n227), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n878), .B(new_n879), .C1(KEYINPUT35), .C2(new_n504), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT36), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n355), .A2(G77), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n226), .A2(new_n882), .B1(G50), .B2(new_n201), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(G1), .A3(new_n637), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT102), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n877), .A2(new_n881), .A3(new_n885), .ZN(G367));
  OAI21_X1  g0686(.A(new_n262), .B1(new_n729), .B2(new_n212), .ZN(new_n887));
  INV_X1    g0687(.A(new_n733), .ZN(new_n888));
  AOI22_X1  g0688(.A1(G143), .A2(new_n742), .B1(new_n888), .B2(G77), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n320), .B2(new_n726), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n887), .B(new_n890), .C1(G159), .C2(new_n737), .ZN(new_n891));
  INV_X1    g0691(.A(new_n709), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(G58), .B1(G137), .B2(new_n723), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n719), .A2(new_n201), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT46), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n709), .A2(new_n898), .A3(new_n246), .ZN(new_n899));
  INV_X1    g0699(.A(G311), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n727), .A2(new_n900), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n715), .A2(new_n488), .B1(new_n726), .B2(new_n418), .ZN(new_n902));
  INV_X1    g0702(.A(G317), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n363), .B1(new_n722), .B2(new_n903), .ZN(new_n904));
  NOR4_X1   g0704(.A1(new_n899), .A2(new_n901), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n730), .A2(new_n805), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n888), .A2(G97), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n898), .B1(new_n709), .B2(new_n246), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n905), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n712), .A2(new_n576), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n896), .A2(new_n897), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT47), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n702), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n544), .A2(new_n645), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n613), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n541), .B2(new_n914), .ZN(new_n916));
  INV_X1    g0716(.A(new_n749), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n756), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n753), .B1(new_n221), .B2(new_n311), .C1(new_n233), .C2(new_n919), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n913), .A2(new_n918), .A3(new_n751), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n656), .A2(KEYINPUT106), .ZN(new_n922));
  INV_X1    g0722(.A(new_n594), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n661), .B1(new_n923), .B2(new_n644), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n924), .A2(new_n664), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT106), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n654), .A2(new_n926), .A3(new_n655), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n925), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n656), .A2(KEYINPUT106), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n501), .A2(new_n645), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n498), .A2(new_n644), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n501), .A2(new_n510), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n664), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n938), .B2(new_n657), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(KEYINPUT44), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n664), .A2(new_n658), .A3(new_n936), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT45), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n939), .A2(KEYINPUT44), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n663), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n700), .B1(new_n932), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n667), .B(KEYINPUT41), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(KEYINPUT107), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT107), .ZN(new_n951));
  INV_X1    g0751(.A(new_n700), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n663), .B(new_n945), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n931), .ZN(new_n954));
  INV_X1    g0754(.A(new_n949), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n252), .B1(new_n638), .B2(G45), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n950), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n663), .A2(new_n937), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n664), .A2(new_n935), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT42), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n501), .B2(new_n644), .C1(new_n658), .C2(new_n935), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n961), .B(new_n966), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n958), .A2(new_n967), .A3(KEYINPUT108), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT108), .B1(new_n958), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n921), .B1(new_n968), .B2(new_n969), .ZN(G387));
  NAND2_X1  g0770(.A1(new_n932), .A2(new_n952), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n931), .A2(new_n700), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n667), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n919), .B1(new_n237), .B2(G45), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n670), .B2(new_n758), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n312), .A2(G50), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT50), .Z(new_n977));
  NOR4_X1   g0777(.A1(new_n977), .A2(G45), .A3(new_n239), .A4(new_n670), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n975), .A2(new_n978), .B1(G107), .B2(new_n221), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n782), .B1(new_n979), .B2(new_n753), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G311), .A2(new_n737), .B1(new_n792), .B2(G317), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n418), .B2(new_n729), .C1(new_n744), .C2(new_n727), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT48), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n576), .B2(new_n709), .C1(new_n715), .C2(new_n806), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT49), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n262), .B1(new_n723), .B2(G326), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(new_n246), .C2(new_n733), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n322), .A2(new_n712), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n719), .A2(new_n311), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G159), .C2(new_n742), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n907), .B1(new_n201), .B2(new_n729), .C1(new_n320), .C2(new_n722), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G77), .B2(new_n892), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n792), .A2(G50), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n262), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n980), .B1(new_n662), .B2(new_n917), .C1(new_n995), .C2(new_n703), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n957), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(new_n931), .B2(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n973), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(G393));
  AOI21_X1  g0801(.A(new_n957), .B1(new_n953), .B2(KEYINPUT110), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT110), .B2(new_n953), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n753), .B1(new_n437), .B2(new_n221), .C1(new_n250), .C2(new_n919), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n751), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT111), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n723), .A2(G143), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G150), .A2(new_n742), .B1(new_n792), .B2(G159), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n262), .B(new_n1007), .C1(new_n1008), .C2(KEYINPUT51), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n719), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(G77), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n729), .A2(new_n312), .B1(new_n733), .B2(new_n375), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G50), .B2(new_n737), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(new_n201), .C2(new_n709), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1009), .B(new_n1014), .C1(KEYINPUT51), .C2(new_n1008), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n727), .A2(new_n903), .B1(new_n726), .B2(new_n900), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT52), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n892), .A2(new_n805), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n730), .A2(G294), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G107), .A2(new_n888), .B1(new_n723), .B2(G322), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n262), .B1(new_n798), .B2(G116), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1017), .B(new_n1022), .C1(G303), .C2(new_n737), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n702), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1006), .B(new_n1024), .C1(new_n917), .C2(new_n936), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n668), .B1(new_n972), .B2(new_n947), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n972), .A2(new_n947), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1003), .B(new_n1025), .C1(new_n1027), .C2(new_n1028), .ZN(G390));
  NAND2_X1  g0829(.A1(new_n857), .A2(new_n747), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n788), .A2(new_n322), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1011), .B1(new_n246), .B2(new_n726), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT116), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n791), .B1(new_n576), .B2(new_n722), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n709), .A2(new_n375), .B1(new_n735), .B2(new_n727), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G97), .C2(new_n730), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n363), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G107), .B2(new_n737), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n892), .A2(G150), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT53), .ZN(new_n1040));
  INV_X1    g0840(.A(G128), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n719), .A2(new_n353), .B1(new_n1041), .B2(new_n727), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT54), .B(G143), .Z(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n262), .B1(new_n212), .B2(new_n733), .C1(new_n1045), .C2(new_n729), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G125), .B2(new_n723), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1043), .B(new_n1047), .C1(new_n794), .C2(new_n712), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G132), .B2(new_n792), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n702), .B1(new_n1038), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1030), .A2(new_n751), .A3(new_n1031), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT112), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n821), .A2(new_n1052), .A3(new_n859), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n820), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n775), .B2(new_n815), .ZN(new_n1055));
  OAI21_X1  g0855(.A(KEYINPUT112), .B1(new_n1055), .B2(new_n860), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n857), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n814), .B1(new_n681), .B2(new_n774), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n859), .B1(new_n1058), .B2(new_n1054), .C1(new_n853), .C2(new_n854), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n774), .B(G330), .C1(new_n696), .C2(new_n697), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1061), .A2(new_n1054), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1062), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1057), .A2(new_n1064), .A3(new_n1059), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1051), .B1(new_n1066), .B2(new_n957), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n862), .A2(new_n634), .A3(new_n871), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1061), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT113), .B1(new_n1069), .B2(new_n820), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT113), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1061), .A2(new_n1054), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n816), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n698), .A2(KEYINPUT114), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT114), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(G330), .C1(new_n696), .C2(new_n697), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1075), .A2(new_n774), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n1054), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n1064), .A3(new_n1058), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1068), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT115), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1063), .A2(new_n1065), .A3(new_n1081), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1083), .A2(new_n667), .A3(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1082), .A2(KEYINPUT115), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1067), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G378));
  NAND2_X1  g0888(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT119), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n867), .A2(new_n869), .A3(new_n1090), .A4(G330), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1092));
  XNOR2_X1  g0892(.A(new_n342), .B(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n326), .A2(new_n822), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1089), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n870), .A2(KEYINPUT119), .A3(new_n1095), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1097), .A2(new_n861), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n861), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT120), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1068), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1084), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1102), .B1(new_n1084), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1101), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT57), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1057), .A2(new_n1064), .A3(new_n1059), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1064), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1058), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1111), .B(new_n1062), .C1(new_n1078), .C2(new_n1054), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n816), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1071), .B1(new_n1061), .B2(new_n1054), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1114), .A2(new_n1062), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1113), .B1(new_n1115), .B2(new_n1072), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1103), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n1109), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT120), .B1(new_n1118), .B2(new_n1068), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1084), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1099), .A2(new_n1100), .A3(new_n1107), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n668), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1108), .A2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1099), .A2(new_n1100), .A3(new_n957), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1095), .A2(new_n748), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n212), .B1(new_n361), .B2(G41), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n892), .A2(G77), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n888), .A2(G58), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n262), .B1(new_n723), .B2(G283), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n729), .A2(new_n311), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G97), .B2(new_n737), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n792), .A2(new_n1134), .A3(G107), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n727), .A2(new_n246), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n792), .B2(G107), .ZN(new_n1137));
  NOR4_X1   g0937(.A1(new_n897), .A2(G41), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1133), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1127), .B1(new_n1139), .B2(KEYINPUT58), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT118), .Z(new_n1141));
  INV_X1    g0941(.A(G41), .ZN(new_n1142));
  AOI21_X1  g0942(.A(G33), .B1(new_n723), .B2(G124), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n729), .A2(new_n794), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G125), .A2(new_n742), .B1(new_n737), .B2(G132), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n1041), .B2(new_n726), .C1(new_n709), .C2(new_n1045), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G150), .C2(new_n1010), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT59), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1142), .B(new_n1143), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G159), .B2(new_n888), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1150), .A2(new_n1151), .B1(KEYINPUT58), .B2(new_n1139), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n703), .B1(new_n1141), .B2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n702), .A2(G50), .A3(new_n747), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n1126), .A2(new_n782), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1125), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1124), .A2(new_n1156), .ZN(G375));
  NAND3_X1  g0957(.A1(new_n1074), .A2(new_n1080), .A3(new_n1068), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1117), .A2(new_n949), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n989), .B1(G294), .B2(new_n742), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n437), .B2(new_n709), .C1(new_n418), .C2(new_n722), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n726), .A2(new_n735), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n729), .A2(new_n488), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n363), .B1(new_n733), .B2(new_n202), .C1(new_n246), .C2(new_n712), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n892), .A2(G159), .B1(new_n737), .B2(new_n1044), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n742), .A2(G132), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT121), .Z(new_n1168));
  OAI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(new_n212), .C2(new_n719), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n729), .A2(new_n320), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n726), .A2(new_n794), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1129), .A2(new_n262), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1172), .A2(KEYINPUT122), .B1(G128), .B2(new_n723), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(KEYINPUT122), .B2(new_n1172), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n702), .B1(new_n1165), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n751), .B(new_n1176), .C1(new_n820), .C2(new_n748), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n201), .B2(new_n788), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n998), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1159), .A2(new_n1180), .ZN(G381));
  NOR2_X1   g0981(.A1(G375), .A2(G378), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G381), .A2(G384), .ZN(new_n1183));
  INV_X1    g0983(.A(G390), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n921), .B(new_n1184), .C1(new_n968), .C2(new_n969), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1185), .A2(G396), .A3(G393), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1183), .A3(new_n1186), .ZN(G407));
  NAND2_X1  g0987(.A1(new_n643), .A2(G213), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT123), .Z(new_n1189));
  NAND2_X1  g0989(.A1(new_n1182), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(G407), .A2(G213), .A3(new_n1190), .ZN(G409));
  NAND2_X1  g0991(.A1(G387), .A2(G390), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1000), .B(new_n767), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1185), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n1192), .B2(new_n1185), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT127), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT61), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1189), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1121), .A2(new_n949), .A3(new_n1101), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1087), .A2(new_n1156), .A3(new_n1200), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1125), .A2(new_n1155), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1108), .B2(new_n1123), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1199), .B(new_n1201), .C1(new_n1203), .C2(new_n1087), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1189), .A2(G2897), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT60), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n668), .B1(new_n1158), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1117), .C1(new_n1207), .C2(new_n1158), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(G384), .A3(new_n1180), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G384), .B1(new_n1209), .B2(new_n1180), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1206), .B1(new_n1213), .B2(KEYINPUT124), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1212), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1210), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT124), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n1205), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1214), .A2(new_n1218), .B1(KEYINPUT124), .B2(new_n1213), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT62), .B1(new_n1204), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1204), .A2(new_n1216), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1198), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1204), .A2(KEYINPUT62), .A3(new_n1216), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1197), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT125), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1204), .A2(new_n1225), .A3(new_n1219), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1196), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT63), .B1(new_n1204), .B2(new_n1216), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1189), .B1(G375), .B2(G378), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT63), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1201), .A4(new_n1213), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1227), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1204), .A2(new_n1219), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT61), .B1(new_n1233), .B2(KEYINPUT125), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT126), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1227), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1231), .A2(new_n1228), .ZN(new_n1237));
  AND4_X1   g1037(.A1(KEYINPUT126), .A2(new_n1236), .A3(new_n1234), .A4(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1224), .B1(new_n1235), .B2(new_n1238), .ZN(G405));
  XNOR2_X1  g1039(.A(new_n1203), .B(G378), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(new_n1216), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(new_n1196), .ZN(G402));
endmodule


