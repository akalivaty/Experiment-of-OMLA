//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1196, new_n1197, new_n1198, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G97), .B(G107), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n207), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n248), .A2(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT65), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT66), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n254), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n215), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n261), .ZN(new_n265));
  INV_X1    g0065(.A(G50), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n266), .B1(new_n206), .B2(G20), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n265), .A2(new_n267), .B1(new_n266), .B2(new_n264), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n273), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(G226), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n279), .A2(new_n280), .B1(new_n224), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n283), .A2(new_n285), .A3(G1698), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n281), .B1(G222), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n271), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n277), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(G200), .B2(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n270), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n296), .B(new_n269), .C1(G179), .C2(new_n289), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n295), .A2(KEYINPUT72), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n278), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G226), .ZN(new_n302));
  INV_X1    g0102(.A(G97), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n301), .A2(new_n302), .B1(new_n284), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n282), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G232), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n307), .A2(new_n308), .A3(new_n300), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n271), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n274), .B1(G238), .B2(new_n276), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n310), .B2(new_n312), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n299), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n299), .C1(new_n313), .C2(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n310), .A2(new_n312), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(G179), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n316), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT71), .B1(new_n263), .B2(G68), .ZN(new_n324));
  XOR2_X1   g0124(.A(new_n324), .B(KEYINPUT12), .Z(new_n325));
  NOR2_X1   g0125(.A1(new_n284), .A2(G20), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n266), .B2(new_n252), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT11), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n328), .A2(new_n329), .A3(new_n261), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n328), .B2(new_n261), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n325), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n261), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(KEYINPUT69), .A3(new_n263), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT69), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n264), .B2(new_n261), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n206), .A2(G20), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G68), .A3(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n339), .A2(KEYINPUT70), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(KEYINPUT70), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n332), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n323), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G200), .B1(new_n313), .B2(new_n314), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n320), .A2(G190), .A3(new_n321), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n265), .ZN(new_n350));
  INV_X1    g0150(.A(new_n248), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n338), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n350), .A2(new_n352), .B1(new_n263), .B2(new_n351), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT7), .B1(new_n307), .B2(new_n207), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  AOI211_X1 g0156(.A(new_n356), .B(G20), .C1(new_n305), .C2(new_n306), .ZN(new_n357));
  OAI21_X1  g0157(.A(G68), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(G58), .A2(G68), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(G20), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G159), .ZN(new_n362));
  NOR4_X1   g0162(.A1(new_n362), .A2(KEYINPUT73), .A3(G20), .A4(G33), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n251), .B2(G159), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n361), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT16), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n356), .B1(new_n278), .B2(G20), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT7), .B(new_n207), .C1(new_n283), .C2(new_n285), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n202), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(KEYINPUT16), .B(new_n361), .C1(new_n363), .C2(new_n365), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n261), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT74), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n368), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n372), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n333), .B1(new_n358), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n371), .B2(new_n366), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT74), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n354), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT18), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n278), .A2(G226), .A3(G1698), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n305), .A2(new_n306), .A3(G223), .A4(new_n300), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n271), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n271), .A2(new_n272), .ZN(new_n388));
  AOI22_X1  g0188(.A1(G232), .A2(new_n276), .B1(new_n388), .B2(new_n275), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n295), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n387), .A2(new_n389), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(G179), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n381), .A2(new_n382), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n387), .A2(new_n389), .ZN(new_n395));
  INV_X1    g0195(.A(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n290), .A2(KEYINPUT75), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n290), .A2(KEYINPUT75), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n387), .A2(new_n389), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n354), .B(new_n402), .C1(new_n375), .C2(new_n380), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n374), .B1(new_n368), .B2(new_n373), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n377), .A2(KEYINPUT74), .A3(new_n379), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n353), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT18), .B1(new_n408), .B2(new_n392), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n402), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n394), .A2(new_n405), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT67), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n326), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n418), .A2(KEYINPUT68), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n248), .A2(new_n252), .B1(new_n207), .B2(new_n224), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n418), .B2(KEYINPUT68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n333), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n337), .A2(G77), .A3(new_n338), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G77), .B2(new_n263), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n279), .A2(new_n219), .B1(new_n226), .B2(new_n278), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n307), .A2(new_n308), .A3(G1698), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n271), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n274), .B1(G244), .B2(new_n276), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n295), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G179), .B2(new_n430), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n428), .A2(G190), .A3(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(G200), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n425), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n298), .A2(new_n349), .A3(new_n411), .A4(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n263), .A2(G97), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n350), .B1(new_n206), .B2(G33), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(G97), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT6), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n303), .A2(new_n226), .ZN(new_n445));
  NOR2_X1   g0245(.A1(G97), .A2(G107), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n226), .A2(KEYINPUT6), .A3(G97), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n450));
  OAI21_X1  g0250(.A(G107), .B1(new_n355), .B2(new_n357), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n443), .B1(new_n452), .B2(new_n261), .ZN(new_n453));
  AOI211_X1 g0253(.A(KEYINPUT76), .B(new_n333), .C1(new_n450), .C2(new_n451), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n442), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n300), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT77), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n301), .A2(new_n225), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(KEYINPUT4), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n271), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G179), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n467), .A2(new_n272), .A3(new_n271), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n288), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(G257), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n462), .A2(new_n463), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT77), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n456), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n459), .A2(new_n458), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n286), .A2(G244), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n288), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n471), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n295), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n455), .A2(new_n472), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT78), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT78), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n455), .A2(new_n472), .A3(new_n481), .A4(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n455), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n479), .A2(new_n480), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G190), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n462), .A2(new_n471), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G200), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n483), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n278), .A2(new_n207), .A3(G68), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n249), .A2(new_n303), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT79), .B(G87), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n495), .A2(G97), .A3(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n497), .A2(new_n207), .ZN(new_n498));
  OAI221_X1 g0298(.A(new_n493), .B1(KEYINPUT19), .B2(new_n494), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(new_n261), .B1(new_n264), .B2(new_n416), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n441), .A2(G87), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n278), .A2(G244), .A3(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n278), .A2(G238), .A3(new_n300), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n271), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n271), .A2(new_n221), .A3(new_n466), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n388), .B2(new_n466), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G190), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n502), .B(new_n511), .C1(new_n396), .C2(new_n510), .ZN(new_n512));
  INV_X1    g0312(.A(new_n441), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n500), .B1(new_n416), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n463), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n514), .B(new_n515), .C1(G169), .C2(new_n510), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n468), .B1(new_n470), .B2(G264), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n286), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n305), .A2(new_n306), .A3(G257), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT82), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT82), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n278), .A2(new_n523), .A3(G257), .A4(G1698), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n519), .B(G179), .C1(new_n526), .C2(new_n288), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n288), .B1(new_n520), .B2(new_n525), .ZN(new_n528));
  INV_X1    g0328(.A(new_n467), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n388), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n469), .B2(new_n227), .ZN(new_n531));
  OAI21_X1  g0331(.A(G169), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT83), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n278), .A2(new_n207), .A3(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n278), .A2(new_n537), .A3(new_n207), .A4(G87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n207), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  INV_X1    g0343(.A(new_n505), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n542), .A2(new_n543), .B1(new_n544), .B2(new_n207), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n539), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n540), .B1(new_n539), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n261), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT25), .B1(new_n264), .B2(new_n226), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n441), .A2(G107), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT83), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n527), .A2(new_n554), .A3(new_n532), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n534), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n528), .A2(new_n531), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(G190), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n559), .A2(new_n548), .A3(new_n552), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n458), .B(new_n207), .C1(G33), .C2(new_n303), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT20), .ZN(new_n564));
  INV_X1    g0364(.A(G116), .ZN(new_n565));
  AOI22_X1  g0365(.A1(KEYINPUT81), .A2(new_n564), .B1(new_n565), .B2(G20), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n566), .A3(new_n261), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n564), .A2(KEYINPUT81), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n567), .B(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n334), .B(new_n336), .C1(G1), .C2(new_n284), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G116), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n263), .A2(new_n565), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G303), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n307), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G257), .A2(G1698), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n227), .B2(G1698), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n575), .B(new_n271), .C1(new_n307), .C2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n467), .A2(new_n288), .A3(G270), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n530), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OR3_X1    g0380(.A1(new_n573), .A2(new_n463), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n530), .A2(new_n578), .A3(KEYINPUT80), .A4(new_n579), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n400), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(G200), .A3(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n573), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT21), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n583), .A2(G169), .A3(new_n584), .ZN(new_n591));
  INV_X1    g0391(.A(new_n573), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n583), .A2(G169), .A3(new_n584), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n594), .A2(KEYINPUT21), .A3(new_n573), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n581), .B(new_n589), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n562), .A2(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n439), .A2(new_n492), .A3(new_n518), .A4(new_n597), .ZN(G372));
  INV_X1    g0398(.A(new_n297), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n405), .A2(new_n410), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n344), .B1(new_n434), .B2(new_n347), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(KEYINPUT84), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(KEYINPUT84), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n394), .A2(new_n409), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n599), .B1(new_n606), .B2(new_n294), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n492), .A2(new_n518), .A3(new_n561), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n581), .B1(new_n593), .B2(new_n595), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n553), .B2(new_n533), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n483), .ZN(new_n612));
  INV_X1    g0412(.A(new_n485), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n518), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT26), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT26), .ZN(new_n616));
  INV_X1    g0416(.A(new_n482), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n518), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n516), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n439), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n607), .A2(new_n620), .ZN(G369));
  NAND3_X1  g0421(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n623));
  XOR2_X1   g0423(.A(new_n623), .B(KEYINPUT85), .Z(new_n624));
  OAI21_X1  g0424(.A(G213), .B1(new_n622), .B2(KEYINPUT27), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n562), .B1(new_n553), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n630), .B(KEYINPUT88), .Z(new_n631));
  INV_X1    g0431(.A(new_n629), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n556), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n632), .A2(new_n573), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n596), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n609), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g0439(.A(KEYINPUT86), .B(G330), .Z(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g0442(.A(new_n642), .B(KEYINPUT87), .Z(new_n643));
  NOR2_X1   g0443(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n609), .A2(new_n632), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n631), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n553), .A2(new_n632), .A3(new_n533), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n644), .A2(new_n648), .ZN(G399));
  INV_X1    g0449(.A(new_n210), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G41), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G1), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n496), .A2(new_n565), .ZN(new_n654));
  OAI22_X1  g0454(.A1(new_n653), .A2(new_n654), .B1(new_n213), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  INV_X1    g0456(.A(new_n609), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n608), .B1(new_n657), .B2(new_n556), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n517), .B2(new_n482), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n516), .B(new_n659), .C1(new_n614), .C2(KEYINPUT26), .ZN(new_n660));
  OAI211_X1 g0460(.A(KEYINPUT29), .B(new_n632), .C1(new_n658), .C2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n619), .ZN(new_n662));
  INV_X1    g0462(.A(new_n611), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n629), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n661), .B1(new_n664), .B2(KEYINPUT29), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n585), .A2(G179), .A3(new_n510), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(new_n489), .A3(new_n558), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n528), .A2(new_n531), .A3(new_n463), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n507), .A2(new_n509), .A3(new_n579), .A4(new_n578), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT91), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT90), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n462), .A3(new_n471), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n527), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n487), .A2(KEYINPUT90), .A3(new_n668), .A4(new_n669), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n671), .B1(new_n672), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT91), .A4(new_n677), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n632), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT92), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT31), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n681), .B2(KEYINPUT31), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n492), .A2(new_n597), .A3(new_n518), .A4(new_n632), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n667), .A2(new_n670), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n678), .ZN(new_n687));
  XNOR2_X1  g0487(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(new_n629), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n683), .A2(new_n684), .A3(new_n685), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n641), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n665), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n656), .B1(new_n694), .B2(G1), .ZN(G364));
  AND2_X1   g0495(.A1(new_n207), .A2(G13), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G45), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G1), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n651), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT93), .Z(new_n700));
  NOR2_X1   g0500(.A1(new_n650), .A2(new_n307), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G355), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(G116), .B2(new_n210), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n650), .A2(new_n278), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n465), .B2(new_n214), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n243), .A2(new_n465), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G13), .A2(G33), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G20), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n215), .B1(G20), .B2(new_n295), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n700), .B1(new_n708), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT94), .B1(new_n207), .B2(new_n463), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n207), .A2(new_n463), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT94), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n586), .A2(new_n396), .A3(new_n716), .A4(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G322), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(G200), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G190), .ZN(new_n724));
  XNOR2_X1  g0524(.A(KEYINPUT33), .B(G317), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n207), .A2(G179), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n290), .A3(G200), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n724), .A2(new_n725), .B1(new_n728), .B2(G283), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G190), .A2(G200), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n278), .B1(new_n732), .B2(G329), .ZN(new_n733));
  INV_X1    g0533(.A(G294), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n290), .A2(G179), .A3(G200), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n207), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n729), .B(new_n733), .C1(new_n734), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n719), .A2(new_n730), .A3(new_n716), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n722), .B(new_n737), .C1(G311), .C2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT96), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT96), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G326), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n400), .A2(new_n723), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT95), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n740), .B1(new_n574), .B2(new_n745), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT97), .Z(new_n750));
  OAI22_X1  g0550(.A1(new_n720), .A2(new_n201), .B1(new_n224), .B2(new_n738), .ZN(new_n751));
  INV_X1    g0551(.A(new_n747), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n752), .A2(new_n266), .B1(new_n226), .B2(new_n727), .ZN(new_n753));
  INV_X1    g0553(.A(new_n724), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n754), .A2(new_n202), .B1(new_n736), .B2(new_n303), .ZN(new_n755));
  OR3_X1    g0555(.A1(new_n731), .A2(KEYINPUT32), .A3(new_n362), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n742), .A2(new_n495), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT32), .B1(new_n731), .B2(new_n362), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n756), .A2(new_n757), .A3(new_n278), .A4(new_n758), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n751), .A2(new_n753), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n750), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT98), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n712), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n715), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n711), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n639), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n700), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n643), .B(new_n769), .C1(new_n641), .C2(new_n639), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(G396));
  OAI21_X1  g0572(.A(new_n629), .B1(new_n422), .B2(new_n424), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n437), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n434), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n433), .A2(new_n632), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n664), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n700), .B1(new_n779), .B2(new_n692), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n692), .B2(new_n779), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n307), .B1(new_n732), .B2(G132), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n782), .B1(new_n201), .B2(new_n736), .C1(new_n202), .C2(new_n727), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n747), .A2(G137), .B1(new_n724), .B2(G150), .ZN(new_n784));
  INV_X1    g0584(.A(G143), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n784), .B1(new_n362), .B2(new_n738), .C1(new_n785), .C2(new_n720), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT34), .Z(new_n787));
  INV_X1    g0587(.A(new_n745), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n783), .B(new_n787), .C1(G50), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n278), .B1(new_n732), .B2(G311), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n303), .B2(new_n736), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n752), .A2(new_n574), .B1(new_n220), .B2(new_n727), .ZN(new_n792));
  INV_X1    g0592(.A(new_n720), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n791), .B(new_n792), .C1(G294), .C2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n226), .B2(new_n745), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n739), .A2(G116), .B1(G283), .B2(new_n724), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT100), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n712), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n712), .A2(new_n709), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT99), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n769), .B1(new_n802), .B2(new_n224), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n799), .B(new_n803), .C1(new_n778), .C2(new_n710), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n781), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G384));
  OR2_X1    g0606(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n807), .A2(G116), .A3(new_n216), .A4(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT36), .Z(new_n810));
  OR3_X1    g0610(.A1(new_n213), .A2(new_n224), .A3(new_n359), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n266), .A2(G68), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n206), .B(G13), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n344), .A2(new_n629), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n381), .A2(new_n393), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n381), .A2(new_n626), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT37), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n403), .ZN(new_n819));
  AOI221_X4 g0619(.A(new_n353), .B1(new_n397), .B2(new_n401), .C1(new_n406), .C2(new_n407), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n358), .A2(KEYINPUT102), .A3(new_n367), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT102), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n371), .B2(new_n366), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n821), .A2(new_n823), .A3(new_n378), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n377), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n392), .B1(new_n825), .B2(new_n354), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n627), .B1(new_n825), .B2(new_n354), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n820), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n819), .B1(new_n828), .B2(new_n818), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n604), .B2(new_n600), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT103), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT38), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n831), .A2(KEYINPUT103), .A3(new_n832), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT104), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n836), .A2(KEYINPUT104), .A3(KEYINPUT39), .A4(new_n837), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT39), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT105), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n408), .A2(new_n627), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n411), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n403), .B1(new_n408), .B2(new_n392), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT37), .B1(new_n848), .B2(new_n845), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n849), .A2(new_n819), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n844), .B1(new_n411), .B2(new_n845), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n843), .B(new_n835), .C1(new_n852), .C2(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT106), .ZN(new_n854));
  INV_X1    g0654(.A(new_n851), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n849), .A2(new_n819), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n846), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n832), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT106), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n843), .A4(new_n835), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT107), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n842), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n842), .B2(new_n861), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n815), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n632), .B1(new_n619), .B2(new_n611), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n776), .B1(new_n866), .B2(new_n777), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n342), .A2(new_n632), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n347), .B1(new_n323), .B2(new_n343), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(KEYINPUT101), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n868), .A2(new_n316), .A3(new_n318), .A4(new_n322), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT101), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n836), .A2(new_n837), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n875), .A2(new_n876), .B1(new_n605), .B2(new_n626), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n865), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n439), .B(new_n661), .C1(new_n664), .C2(KEYINPUT29), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(new_n607), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT108), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n879), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n678), .A2(new_n672), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n680), .A3(new_n686), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n886), .B(new_n685), .C1(new_n681), .C2(new_n689), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n777), .A2(new_n870), .A3(new_n873), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT40), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT109), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n858), .A2(new_n890), .A3(new_n835), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n411), .A2(new_n845), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(KEYINPUT105), .B1(new_n819), .B2(new_n849), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n893), .B2(new_n846), .ZN(new_n894));
  INV_X1    g0694(.A(new_n835), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT109), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n887), .A2(new_n888), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n898), .B1(new_n876), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n439), .A2(new_n887), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n640), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n902), .B2(new_n901), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n883), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n206), .B2(new_n696), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n883), .A2(new_n904), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n814), .B1(new_n906), .B2(new_n907), .ZN(G367));
  OAI21_X1  g0708(.A(new_n492), .B1(new_n486), .B2(new_n632), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n617), .A2(new_n629), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n631), .A2(new_n645), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n911), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n483), .B(new_n485), .C1(new_n913), .C2(new_n556), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n912), .A2(KEYINPUT42), .B1(new_n914), .B2(new_n632), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(KEYINPUT42), .B2(new_n912), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n632), .A2(new_n502), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n518), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n917), .A2(new_n516), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n916), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n644), .A2(new_n911), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n921), .B1(new_n916), .B2(new_n922), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n651), .B(KEYINPUT41), .Z(new_n929));
  INV_X1    g0729(.A(new_n644), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n648), .A2(new_n913), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT44), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n646), .A2(new_n647), .A3(new_n911), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT45), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n930), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n932), .A2(new_n644), .A3(new_n935), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n646), .B1(new_n634), .B2(new_n645), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(new_n643), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n693), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n929), .B1(new_n943), .B2(new_n694), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n698), .B(KEYINPUT110), .Z(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n927), .B(new_n928), .C1(new_n944), .C2(new_n946), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n713), .B1(new_n210), .B2(new_n416), .C1(new_n705), .C2(new_n239), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n700), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n736), .A2(new_n202), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G77), .B2(new_n728), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n201), .B2(new_n741), .ZN(new_n952));
  INV_X1    g0752(.A(G137), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n278), .B1(new_n731), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G159), .B2(new_n724), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n266), .B2(new_n738), .C1(new_n250), .C2(new_n720), .ZN(new_n956));
  INV_X1    g0756(.A(new_n748), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n952), .B(new_n956), .C1(G143), .C2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n736), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G107), .A2(new_n959), .B1(new_n724), .B2(G294), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n728), .A2(G97), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n278), .B1(new_n732), .B2(G317), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n788), .A2(KEYINPUT46), .A3(G116), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT46), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n741), .B2(new_n565), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT112), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(KEYINPUT112), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n964), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n963), .B(new_n969), .C1(G283), .C2(new_n739), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n957), .A2(G311), .B1(G303), .B2(new_n793), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT111), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n958), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n949), .B1(new_n920), .B2(new_n767), .C1(new_n974), .C2(new_n764), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n947), .A2(new_n975), .ZN(G387));
  NAND2_X1  g0776(.A1(new_n417), .A2(new_n959), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n202), .B2(new_n738), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n747), .A2(G159), .B1(new_n724), .B2(new_n351), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n278), .A3(new_n961), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT113), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n741), .A2(new_n224), .B1(new_n731), .B2(new_n250), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n981), .B2(new_n982), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n978), .B(new_n984), .C1(G50), .C2(new_n793), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT114), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n793), .A2(G317), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n739), .A2(G303), .B1(G311), .B2(new_n724), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n748), .C2(new_n721), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT48), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n959), .A2(G283), .B1(new_n742), .B2(G294), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT49), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n307), .B1(new_n731), .B2(new_n746), .C1(new_n565), .C2(new_n727), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n764), .B1(new_n986), .B2(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n236), .A2(new_n465), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n1001), .A2(new_n704), .B1(new_n654), .B2(new_n701), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n351), .B2(new_n266), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n465), .B1(new_n202), .B2(new_n224), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n248), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n654), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1002), .A2(new_n1007), .B1(G107), .B2(new_n210), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n769), .B(new_n1000), .C1(new_n713), .C2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT115), .Z(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n635), .B2(new_n711), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n941), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n946), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n694), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n942), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n651), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(G393));
  OAI21_X1  g0817(.A(new_n1015), .B1(new_n937), .B2(new_n938), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n943), .A2(new_n651), .A3(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n793), .A2(G311), .B1(G317), .B2(new_n747), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT52), .Z(new_n1021));
  OAI221_X1 g0821(.A(new_n307), .B1(new_n731), .B2(new_n721), .C1(new_n226), .C2(new_n727), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G116), .A2(new_n959), .B1(new_n724), .B2(G303), .ZN(new_n1023));
  INV_X1    g0823(.A(G283), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n1024), .B2(new_n741), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1022), .B(new_n1025), .C1(G294), .C2(new_n739), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1021), .A2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n720), .A2(new_n362), .B1(new_n752), .B2(new_n250), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT51), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n742), .A2(G68), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G77), .A2(new_n959), .B1(new_n724), .B2(G50), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n278), .B1(new_n731), .B2(new_n785), .C1(new_n220), .C2(new_n727), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n351), .B2(new_n739), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n764), .B1(new_n1027), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n705), .A2(new_n246), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n714), .B(new_n1036), .C1(G97), .C2(new_n650), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1035), .A2(new_n769), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n911), .B2(new_n767), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1019), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n939), .A2(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n939), .A2(KEYINPUT116), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n946), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1040), .A2(new_n1043), .ZN(G390));
  AND2_X1   g0844(.A1(new_n887), .A2(G330), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n439), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n881), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n778), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n874), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT117), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(KEYINPUT117), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n632), .B(new_n775), .C1(new_n658), .C2(new_n660), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1053), .A2(new_n776), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n691), .A2(new_n641), .A3(new_n888), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1049), .B1(new_n692), .B2(new_n777), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1045), .A2(new_n888), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n867), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1047), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n864), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n815), .B1(new_n867), .B2(new_n874), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n842), .A2(new_n861), .A3(new_n862), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1054), .A2(new_n1049), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n815), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n891), .A2(new_n896), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1067), .A2(new_n1055), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1058), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1062), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1058), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n863), .A2(new_n864), .A3(new_n1064), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1071), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1067), .A2(new_n1055), .A3(new_n1071), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n1061), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1074), .A2(new_n651), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n946), .A3(new_n1079), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT119), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n769), .B1(new_n802), .B2(new_n248), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n720), .A2(new_n565), .B1(new_n303), .B2(new_n738), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n278), .B1(new_n959), .B2(G77), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n754), .B2(new_n226), .C1(new_n1024), .C2(new_n752), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(G87), .C2(new_n788), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n727), .A2(new_n202), .B1(new_n731), .B2(new_n734), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT118), .ZN(new_n1090));
  INV_X1    g0890(.A(G128), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n752), .A2(new_n1091), .B1(new_n362), .B2(new_n736), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n307), .B1(new_n732), .B2(G125), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1093), .B1(new_n738), .B2(new_n1094), .C1(new_n754), .C2(new_n953), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1092), .B(new_n1095), .C1(G50), .C2(new_n728), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n742), .A2(G150), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(KEYINPUT53), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1097), .A2(KEYINPUT53), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(G132), .C2(new_n793), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1088), .A2(new_n1090), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1084), .B1(new_n764), .B2(new_n1101), .C1(new_n1102), .C2(new_n710), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1082), .A2(new_n1083), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1083), .B1(new_n1082), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1081), .B1(new_n1104), .B2(new_n1105), .ZN(G378));
  AOI21_X1  g0906(.A(new_n298), .B1(new_n269), .B2(new_n626), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n269), .A2(new_n626), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n294), .B2(new_n297), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n709), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n700), .B1(new_n801), .B2(G50), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n278), .A2(G41), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n266), .B1(G33), .B2(G41), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1024), .B2(new_n731), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n950), .B(new_n1120), .C1(new_n793), .C2(G107), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n724), .A2(G97), .B1(new_n742), .B2(G77), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n747), .A2(G116), .B1(G58), .B2(new_n728), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n417), .A2(new_n739), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT58), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1119), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n720), .A2(new_n1091), .B1(new_n953), .B2(new_n738), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n747), .A2(G125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n959), .A2(G150), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n724), .A2(G132), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n741), .A2(new_n1094), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n728), .A2(G159), .ZN(new_n1138));
  AOI211_X1 g0938(.A(G33), .B(G41), .C1(new_n732), .C2(G124), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1127), .B1(new_n1126), .B2(new_n1125), .C1(new_n1136), .C2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1116), .B1(new_n1141), .B2(new_n712), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1115), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n897), .A2(G330), .A3(new_n900), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1114), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1146), .A2(new_n897), .A3(G330), .A4(new_n900), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n879), .B2(KEYINPUT120), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n879), .A2(KEYINPUT120), .A3(new_n1149), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1143), .B1(new_n1153), .B2(new_n945), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1047), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1080), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT120), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1157), .B(new_n1148), .C1(new_n865), .C2(new_n878), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT57), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n879), .A2(new_n1148), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1149), .A2(new_n865), .A3(new_n878), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1161), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n652), .B1(new_n1156), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1154), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(G375));
  OAI21_X1  g0968(.A(new_n700), .B1(new_n801), .B2(G68), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n307), .B1(new_n731), .B2(new_n574), .C1(new_n224), .C2(new_n727), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n752), .A2(new_n734), .B1(new_n754), .B2(new_n565), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G97), .C2(new_n788), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n739), .A2(G107), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n793), .A2(G283), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1172), .A2(new_n977), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n278), .B1(new_n731), .B2(new_n1091), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G58), .B2(new_n728), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n250), .B2(new_n738), .C1(new_n953), .C2(new_n720), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n747), .A2(G132), .B1(new_n959), .B2(G50), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n754), .B2(new_n1094), .C1(new_n745), .C2(new_n362), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1175), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1169), .B1(new_n1181), .B2(new_n712), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT121), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1049), .B2(new_n709), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1185), .B2(new_n946), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1061), .A2(new_n929), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1185), .A2(new_n1155), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(G381));
  NAND4_X1  g0989(.A1(new_n947), .A2(new_n1040), .A3(new_n975), .A4(new_n1043), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1081), .A2(new_n1082), .A3(new_n1103), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1167), .A3(new_n1193), .A4(new_n1194), .ZN(G407));
  NAND2_X1  g0995(.A1(new_n628), .A2(G213), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1167), .A2(new_n1193), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(G407), .A2(G213), .A3(new_n1198), .ZN(G409));
  XNOR2_X1  g0999(.A(G393), .B(new_n771), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n947), .A2(new_n975), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1201));
  OAI211_X1 g1001(.A(KEYINPUT125), .B(new_n1200), .C1(new_n1191), .C2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(G387), .A2(G390), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1200), .A2(KEYINPUT125), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(KEYINPUT125), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1203), .A2(new_n1190), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1202), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1056), .A2(KEYINPUT60), .A3(new_n1060), .A4(new_n1047), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT123), .Z(new_n1209));
  OAI211_X1 g1009(.A(new_n651), .B(new_n1062), .C1(new_n1188), .C2(KEYINPUT60), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1186), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n805), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G384), .B(new_n1186), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1197), .A2(G2897), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1160), .A2(new_n929), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1143), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(new_n946), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1192), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1219), .B1(new_n1159), .B2(new_n946), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1156), .A2(new_n1165), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n651), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G378), .B(new_n1223), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT122), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT122), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1167), .A2(new_n1229), .A3(G378), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1222), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1217), .B1(new_n1231), .B2(new_n1197), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1207), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1231), .A2(new_n1197), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT63), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1222), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1227), .A2(KEYINPUT122), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1229), .B1(new_n1167), .B2(G378), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1235), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1196), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT63), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1243), .A2(KEYINPUT124), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT124), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1234), .B(new_n1237), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1232), .A2(KEYINPUT126), .A3(new_n1233), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1241), .A2(new_n1196), .A3(new_n1242), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT127), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT62), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1236), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT126), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1248), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1247), .B1(new_n1255), .B2(new_n1207), .ZN(G405));
  NAND2_X1  g1056(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G375), .A2(new_n1193), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(new_n1235), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(new_n1207), .ZN(G402));
endmodule


