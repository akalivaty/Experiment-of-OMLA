//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  INV_X1    g011(.A(G110), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(new_n197), .A3(new_n198), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n194), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(KEYINPUT24), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n198), .A2(KEYINPUT24), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n192), .B1(new_n201), .B2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT74), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT74), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n208), .A3(new_n211), .A4(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n206), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n206), .A2(new_n210), .A3(KEYINPUT75), .A4(new_n212), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n196), .A2(new_n197), .A3(new_n200), .ZN(new_n217));
  INV_X1    g031(.A(new_n202), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n204), .A2(new_n203), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n217), .A2(G110), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(G146), .B1(new_n207), .B2(new_n208), .ZN(new_n221));
  INV_X1    g035(.A(new_n209), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n220), .B(KEYINPUT73), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n221), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n209), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT73), .B1(new_n226), .B2(new_n220), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n215), .B(new_n216), .C1(new_n224), .C2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G137), .ZN(new_n229));
  INV_X1    g043(.A(G953), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(G221), .A3(G234), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n229), .B(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n220), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n223), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n238), .A2(new_n216), .A3(new_n215), .A4(new_n232), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G234), .ZN(new_n241));
  OAI21_X1  g055(.A(G217), .B1(new_n241), .B2(G902), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n234), .A2(new_n239), .A3(new_n243), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT25), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n234), .A2(new_n239), .A3(new_n243), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n242), .B(KEYINPUT72), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n245), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT65), .B(KEYINPUT1), .C1(new_n259), .C2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G128), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT65), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n258), .A3(new_n260), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G137), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G134), .ZN(new_n272));
  OAI21_X1  g086(.A(G131), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT11), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n269), .B2(G137), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(KEYINPUT11), .A3(G134), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT64), .B(G131), .Z(new_n279));
  OAI21_X1  g093(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(G131), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT64), .B(G131), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n283), .A2(new_n275), .A3(new_n276), .A4(new_n277), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT0), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(new_n193), .ZN(new_n287));
  NOR2_X1   g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n261), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(G143), .B(G146), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n286), .B2(new_n193), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n268), .A2(new_n281), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(KEYINPUT2), .A2(G113), .ZN(new_n294));
  AND3_X1   g108(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n199), .A2(G116), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n298), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n298), .B2(new_n300), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n302), .B1(new_n306), .B2(new_n297), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n256), .B1(new_n293), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n280), .B1(new_n267), .B2(new_n265), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n282), .A2(new_n284), .B1(new_n289), .B2(new_n291), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n299), .A2(G119), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n199), .A2(G116), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT67), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n298), .A2(new_n300), .A3(new_n303), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n297), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G116), .B(G119), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n316), .B(new_n294), .C1(new_n296), .C2(new_n295), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NOR4_X1   g132(.A1(new_n309), .A2(new_n310), .A3(new_n318), .A4(KEYINPUT68), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n308), .A2(new_n319), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT30), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n268), .A2(new_n281), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n285), .A2(new_n292), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n318), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G237), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n230), .A3(G210), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT27), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G101), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT69), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT31), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n320), .A2(new_n326), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n332), .A2(KEYINPUT31), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n267), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT1), .B1(new_n259), .B2(G146), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(G128), .A3(new_n262), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n341), .B2(new_n261), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n324), .B(new_n307), .C1(new_n342), .C2(new_n280), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT68), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n293), .A2(new_n256), .A3(new_n307), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT30), .B1(new_n309), .B2(new_n310), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n324), .B(new_n322), .C1(new_n342), .C2(new_n280), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n307), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n335), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n331), .A3(new_n333), .A4(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n318), .B1(new_n309), .B2(new_n310), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n344), .A2(new_n353), .A3(new_n345), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT28), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n343), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n331), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n336), .A2(new_n352), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(G472), .A2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT32), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n359), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n346), .A2(new_n349), .A3(new_n359), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n351), .B1(new_n365), .B2(new_n333), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n334), .A2(new_n335), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(new_n361), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n343), .A2(KEYINPUT70), .A3(new_n356), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT70), .B1(new_n343), .B2(new_n356), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n331), .A2(KEYINPUT29), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n355), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n243), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(KEYINPUT71), .A3(new_n243), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n320), .A2(new_n326), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n381), .B2(new_n359), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n358), .B2(new_n359), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G472), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n255), .B1(new_n371), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT89), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n259), .A2(G128), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n193), .A2(G143), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n269), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n389), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G134), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n299), .A2(G122), .ZN(new_n393));
  INV_X1    g207(.A(G122), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT87), .B1(new_n394), .B2(G116), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n299), .A3(G122), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G107), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n390), .A2(new_n392), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n395), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n393), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n387), .B(new_n400), .C1(new_n406), .C2(new_n399), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n393), .B1(new_n401), .B2(KEYINPUT14), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n399), .B1(new_n408), .B2(new_n404), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n392), .A2(new_n390), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n398), .A2(new_n399), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT89), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n388), .A3(new_n389), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(G134), .C1(new_n388), .C2(new_n414), .ZN(new_n416));
  INV_X1    g230(.A(new_n411), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n398), .A2(new_n399), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n416), .B(new_n390), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n407), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT9), .B(G234), .ZN(new_n421));
  INV_X1    g235(.A(G217), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n421), .A2(new_n422), .A3(G953), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n407), .A2(new_n413), .A3(new_n419), .A4(new_n423), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(KEYINPUT90), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT90), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(new_n428), .A3(new_n424), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n243), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G478), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(KEYINPUT15), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n430), .B(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n327), .A2(new_n230), .A3(G143), .A4(G214), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n327), .A2(new_n230), .A3(G214), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n327), .A2(new_n230), .A3(KEYINPUT82), .A4(G214), .ZN(new_n441));
  AND4_X1   g255(.A1(KEYINPUT83), .A2(new_n440), .A3(new_n259), .A4(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(G143), .B1(new_n438), .B2(new_n439), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT83), .B1(new_n443), .B2(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n437), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(KEYINPUT18), .A3(G131), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT18), .A2(G131), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(new_n437), .C1(new_n442), .C2(new_n444), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n257), .B1(new_n188), .B2(new_n190), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n446), .B(new_n448), .C1(new_n192), .C2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n445), .A2(KEYINPUT17), .A3(new_n279), .ZN(new_n451));
  INV_X1    g265(.A(new_n226), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(KEYINPUT85), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n445), .A2(new_n279), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT17), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n437), .B(new_n283), .C1(new_n442), .C2(new_n444), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT85), .B1(new_n451), .B2(new_n452), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n450), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(G104), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n450), .B(new_n464), .C1(new_n458), .C2(new_n459), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n243), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G475), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n460), .A2(new_n463), .ZN(new_n470));
  INV_X1    g284(.A(new_n463), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n450), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n191), .B(KEYINPUT19), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n210), .B(new_n212), .C1(new_n473), .C2(G146), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n454), .B2(new_n456), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(G475), .A2(G902), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n472), .A2(new_n475), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n460), .B2(new_n463), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(KEYINPUT20), .A3(new_n477), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n434), .A2(new_n469), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT3), .B1(new_n462), .B2(G107), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n399), .A3(G104), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n462), .A2(G107), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G101), .ZN(new_n490));
  INV_X1    g304(.A(G101), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n485), .A2(new_n487), .A3(new_n491), .A4(new_n488), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n494), .A3(G101), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n318), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n462), .A2(G107), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n399), .A2(G104), .ZN(new_n498));
  OAI21_X1  g312(.A(G101), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT5), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n313), .B2(new_n314), .ZN(new_n502));
  OAI21_X1  g316(.A(G113), .B1(new_n298), .B2(KEYINPUT5), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n500), .B(new_n317), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G110), .B(G122), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n496), .A2(new_n504), .A3(new_n506), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(KEYINPUT6), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n292), .A2(G125), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n342), .B2(G125), .ZN(new_n512));
  INV_X1    g326(.A(G224), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(G953), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n512), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n517), .A3(new_n507), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n512), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n492), .A2(new_n499), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(new_n317), .C1(new_n502), .C2(new_n503), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n301), .A2(new_n501), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n317), .B1(new_n524), .B2(new_n503), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n500), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n506), .B(KEYINPUT8), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n509), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(G902), .B1(new_n521), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(G210), .B1(G237), .B2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n519), .A2(new_n530), .A3(new_n532), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT81), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G214), .B1(G237), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT81), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n531), .A2(new_n538), .A3(new_n533), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(KEYINPUT91), .A2(G952), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(KEYINPUT91), .A2(G952), .ZN(new_n543));
  AOI21_X1  g357(.A(G953), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n241), .B2(new_n327), .ZN(new_n545));
  AOI211_X1 g359(.A(new_n243), .B(new_n230), .C1(G234), .C2(G237), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT21), .B(G898), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n484), .A2(new_n540), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n338), .A2(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n261), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n267), .A2(KEYINPUT77), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT77), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n290), .A2(new_n554), .A3(new_n266), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n500), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n282), .A2(new_n284), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n493), .A2(new_n292), .A3(new_n495), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n492), .A2(new_n499), .A3(KEYINPUT10), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n268), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n265), .A2(new_n522), .A3(new_n267), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT12), .B1(new_n566), .B2(new_n285), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n568), .B(new_n560), .C1(new_n557), .C2(new_n565), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n564), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G140), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n230), .A2(G227), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n573), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n564), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n559), .A2(new_n561), .A3(new_n563), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n285), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G469), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT79), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT79), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n570), .A2(new_n573), .B1(new_n576), .B2(new_n578), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(G469), .C1(new_n584), .C2(G902), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n564), .B(new_n575), .C1(new_n567), .C2(new_n569), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n575), .B1(new_n578), .B2(new_n564), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n581), .B(new_n243), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT80), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT80), .ZN(new_n591));
  INV_X1    g405(.A(new_n564), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n557), .A2(new_n558), .B1(new_n268), .B2(new_n562), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n560), .B1(new_n593), .B2(new_n561), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n573), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n595), .B2(new_n586), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n591), .B1(new_n596), .B2(new_n581), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n582), .B(new_n585), .C1(new_n590), .C2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G221), .B1(new_n421), .B2(G902), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n386), .A2(new_n550), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  INV_X1    g416(.A(new_n537), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n534), .B2(new_n535), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n605), .A2(new_n549), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n469), .A2(new_n480), .A3(new_n483), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT93), .B(G478), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n430), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n426), .B(KEYINPUT92), .Z(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(KEYINPUT33), .A3(new_n425), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n427), .A2(new_n613), .A3(new_n429), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n243), .A2(G478), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n608), .A2(new_n617), .A3(KEYINPUT94), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT94), .B1(new_n608), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n607), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n598), .A2(new_n599), .A3(new_n254), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n360), .B2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n368), .A2(new_n361), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT34), .B(G104), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  XOR2_X1   g444(.A(new_n549), .B(KEYINPUT95), .Z(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR4_X1   g446(.A1(new_n608), .A2(new_n605), .A3(new_n434), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n626), .A3(new_n622), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NAND2_X1  g450(.A1(new_n252), .A2(new_n253), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n233), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n228), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n243), .A3(new_n242), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n598), .A2(new_n599), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n550), .A2(new_n626), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT96), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n643), .B(new_n645), .ZN(G12));
  AOI22_X1  g460(.A1(new_n363), .A2(new_n370), .B1(new_n384), .B2(G472), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n598), .A2(new_n599), .A3(new_n641), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n479), .A2(new_n478), .B1(new_n468), .B2(G475), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n430), .A2(new_n432), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n430), .A2(new_n432), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n546), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n545), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n651), .A2(new_n654), .A3(new_n483), .A4(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n650), .B1(new_n659), .B2(new_n605), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n654), .A2(new_n469), .A3(new_n480), .A4(new_n483), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n661), .A2(KEYINPUT97), .A3(new_n604), .A4(new_n658), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n649), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT98), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n649), .A2(new_n660), .A3(new_n662), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n381), .A2(new_n331), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n243), .C1(new_n354), .C2(new_n331), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G472), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n371), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n371), .A2(KEYINPUT99), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n603), .B1(new_n652), .B2(new_n653), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n608), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n536), .A2(new_n539), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(KEYINPUT38), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT38), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n536), .B2(new_n539), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n679), .A2(new_n681), .A3(new_n683), .A4(new_n641), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n657), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n598), .A2(new_n599), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT40), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n669), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n689), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n677), .A3(KEYINPUT101), .A4(new_n684), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT102), .B(G143), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G45));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n608), .A2(new_n617), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n696), .B1(new_n697), .B2(new_n657), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n608), .A2(new_n617), .A3(KEYINPUT103), .A4(new_n658), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n647), .A2(new_n648), .A3(new_n605), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NAND2_X1  g517(.A1(new_n595), .A2(new_n586), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n581), .B1(new_n704), .B2(new_n243), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n589), .A2(KEYINPUT80), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n596), .A2(new_n591), .A3(new_n581), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n599), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n647), .A2(new_n255), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT94), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n697), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n618), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n713), .A3(new_n607), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  INV_X1    g530(.A(new_n599), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n717), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n386), .A2(new_n633), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT104), .B(G116), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G18));
  NAND4_X1  g535(.A1(new_n641), .A2(new_n708), .A3(new_n599), .A4(new_n604), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n647), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n484), .A2(new_n549), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NAND2_X1  g540(.A1(new_n534), .A2(new_n535), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n608), .A2(new_n727), .A3(new_n631), .A4(new_n678), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n355), .A2(new_n374), .ZN(new_n730));
  OAI22_X1  g544(.A1(new_n366), .A2(new_n367), .B1(new_n730), .B2(new_n331), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n361), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n623), .A2(new_n732), .A3(new_n254), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n709), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n734), .A3(KEYINPUT105), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n718), .A2(new_n254), .A3(new_n623), .A4(new_n732), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n736), .B1(new_n737), .B2(new_n728), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  NAND3_X1  g554(.A1(new_n641), .A2(new_n623), .A3(new_n732), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n708), .A2(new_n599), .A3(new_n604), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n698), .A2(new_n699), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n189), .ZN(G27));
  NAND2_X1  g559(.A1(new_n574), .A2(new_n579), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n581), .B1(new_n746), .B2(new_n243), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n706), .B2(new_n707), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT106), .B1(new_n748), .B2(new_n717), .ZN(new_n749));
  OAI21_X1  g563(.A(G469), .B1(new_n584), .B2(G902), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n590), .B2(new_n597), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n599), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n680), .A2(new_n537), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n386), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n700), .A2(new_n757), .A3(KEYINPUT42), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n386), .A2(new_n754), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n698), .A2(new_n699), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  INV_X1    g578(.A(new_n659), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n386), .A2(new_n754), .A3(new_n765), .A4(new_n756), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  INV_X1    g581(.A(new_n608), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n617), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n771), .A3(new_n617), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT107), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n625), .A2(new_n641), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT108), .Z(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(KEYINPUT107), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n774), .A2(new_n776), .A3(KEYINPUT44), .A4(new_n777), .ZN(new_n781));
  NAND2_X1  g595(.A1(G469), .A2(G902), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n584), .A2(KEYINPUT45), .ZN(new_n783));
  OAI21_X1  g597(.A(G469), .B1(new_n584), .B2(KEYINPUT45), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n706), .A2(new_n707), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n783), .A2(new_n784), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n782), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n717), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n792), .A2(new_n687), .A3(new_n756), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n780), .A2(new_n781), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  XOR2_X1   g609(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n796));
  OR2_X1    g610(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n700), .A2(new_n647), .A3(new_n255), .A4(new_n756), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n187), .ZN(G42));
  NOR2_X1   g617(.A1(new_n773), .A2(new_n545), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n755), .A2(new_n709), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n386), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT48), .ZN(new_n807));
  INV_X1    g621(.A(new_n545), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n770), .A2(new_n808), .A3(new_n734), .A4(new_n772), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n605), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT117), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n755), .A2(new_n709), .A3(new_n545), .A4(new_n255), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n713), .A3(new_n675), .A4(new_n676), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n544), .A2(new_n807), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  INV_X1    g629(.A(new_n733), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n804), .A2(new_n816), .A3(new_n756), .ZN(new_n817));
  INV_X1    g631(.A(new_n800), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n708), .A2(new_n717), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n820), .B1(new_n800), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n817), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n603), .B1(new_n681), .B2(new_n683), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n809), .A2(KEYINPUT114), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n826), .B2(KEYINPUT115), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n608), .A2(new_n617), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n812), .A2(new_n675), .A3(new_n676), .A4(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT116), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n809), .A2(new_n825), .B1(KEYINPUT114), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n741), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n804), .A2(new_n833), .A3(new_n805), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n827), .A2(new_n830), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n815), .B1(new_n823), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n818), .A2(new_n820), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT51), .B1(new_n837), .B2(new_n817), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n814), .B(new_n836), .C1(new_n835), .C2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n710), .A2(new_n633), .B1(new_n723), .B2(new_n724), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n843), .A2(new_n714), .A3(new_n739), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n763), .A3(KEYINPUT53), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n651), .A2(new_n654), .A3(new_n483), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n697), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n540), .A2(new_n632), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n622), .A3(new_n626), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n766), .A2(new_n849), .A3(new_n601), .A4(new_n643), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n623), .A2(new_n732), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n749), .B2(new_n753), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n698), .A3(new_n699), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n371), .A2(new_n385), .ZN(new_n855));
  INV_X1    g669(.A(new_n484), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n600), .A3(new_n856), .A4(new_n658), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n756), .A2(new_n641), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT111), .B1(new_n851), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n854), .B2(new_n857), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n850), .A3(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n845), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n744), .B1(new_n664), .B2(new_n666), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(KEYINPUT110), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT110), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n869), .B(new_n744), .C1(new_n664), .C2(new_n666), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n608), .A2(new_n727), .A3(new_n678), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n637), .A2(new_n640), .A3(new_n658), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n871), .A2(new_n717), .A3(new_n748), .A4(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n700), .A2(new_n701), .B1(new_n677), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT52), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n868), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT52), .B1(new_n867), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n866), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n863), .A2(new_n850), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n879), .A2(new_n844), .A3(new_n763), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n867), .A2(KEYINPUT52), .A3(new_n874), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n880), .B1(new_n881), .B2(new_n877), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n842), .B1(new_n885), .B2(KEYINPUT54), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n878), .A2(new_n884), .A3(KEYINPUT112), .A4(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n883), .B(new_n880), .C1(new_n876), .C2(new_n877), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n882), .A2(KEYINPUT53), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n841), .A2(new_n892), .B1(G952), .B2(G953), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n708), .B(KEYINPUT49), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n537), .A3(new_n599), .A4(new_n254), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n681), .A2(new_n683), .ZN(new_n896));
  OR4_X1    g710(.A1(new_n677), .A2(new_n895), .A3(new_n896), .A4(new_n769), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n230), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n243), .B1(new_n878), .B2(new_n884), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT56), .B1(new_n901), .B2(G210), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n510), .A2(new_n518), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT119), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT120), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(new_n516), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n900), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  AOI211_X1 g723(.A(KEYINPUT56), .B(new_n907), .C1(new_n901), .C2(G210), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n885), .A2(G210), .A3(G902), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n907), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n902), .A2(new_n908), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .A4(new_n900), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n911), .A2(new_n918), .ZN(G51));
  XNOR2_X1  g733(.A(new_n885), .B(new_n887), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n782), .B(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n704), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n901), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n923), .A2(new_n790), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n899), .B1(new_n922), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  INV_X1    g740(.A(new_n482), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n899), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n612), .A2(new_n614), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n900), .B1(new_n920), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n892), .A2(new_n933), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n615), .ZN(G63));
  XOR2_X1   g751(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND3_X1  g754(.A1(new_n885), .A2(new_n639), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n843), .A2(new_n739), .A3(new_n714), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n762), .B2(new_n758), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n864), .B1(new_n863), .B2(new_n850), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n851), .A2(new_n861), .A3(KEYINPUT111), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n943), .A2(KEYINPUT53), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n744), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n667), .A2(new_n947), .A3(new_n874), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT52), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n667), .A2(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n869), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n867), .A2(KEYINPUT110), .ZN(new_n953));
  INV_X1    g767(.A(new_n875), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n946), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n867), .A2(KEYINPUT52), .A3(new_n874), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n950), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT53), .B1(new_n958), .B2(new_n880), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n940), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n899), .B1(new_n960), .B2(new_n240), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n941), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g777(.A(KEYINPUT123), .B(new_n899), .C1(new_n960), .C2(new_n240), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n938), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n961), .A2(KEYINPUT61), .A3(new_n941), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(G66));
  NAND4_X1  g781(.A1(new_n844), .A2(new_n601), .A3(new_n643), .A4(new_n849), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n230), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n547), .B2(new_n513), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT124), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n904), .B1(G898), .B2(new_n230), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n975), .B(new_n976), .Z(G69));
  NAND2_X1  g791(.A1(new_n347), .A2(new_n348), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n473), .B(KEYINPUT126), .Z(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(G953), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n952), .A2(new_n693), .A3(new_n702), .A4(new_n953), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n868), .A2(new_n870), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(KEYINPUT62), .A3(new_n693), .A4(new_n702), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n802), .ZN(new_n988));
  INV_X1    g802(.A(new_n688), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n386), .A2(new_n847), .A3(new_n989), .A4(new_n756), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n794), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n987), .A2(KEYINPUT127), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT127), .B1(new_n987), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n981), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(G227), .ZN(new_n995));
  OAI21_X1  g809(.A(G953), .B1(new_n995), .B2(new_n655), .ZN(new_n996));
  NAND2_X1  g810(.A1(G900), .A2(G953), .ZN(new_n997));
  INV_X1    g811(.A(new_n871), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n792), .A2(new_n386), .A3(new_n687), .A4(new_n998), .ZN(new_n999));
  AND4_X1   g813(.A1(new_n763), .A2(new_n988), .A3(new_n766), .A4(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n1000), .A2(new_n702), .A3(new_n794), .A4(new_n985), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n997), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n980), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n994), .A2(new_n996), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n996), .B1(new_n994), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n1001), .B2(new_n968), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1009), .A2(new_n359), .A3(new_n350), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n350), .B(new_n331), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n889), .A2(new_n890), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1010), .A2(new_n900), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n993), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n987), .A2(KEYINPUT127), .A3(new_n991), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1008), .B1(new_n1016), .B2(new_n968), .ZN(new_n1017));
  INV_X1    g831(.A(new_n670), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(G57));
endmodule


