//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT66), .Z(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT67), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n215), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT64), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n221), .A2(G1), .A3(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NAND4_X1  g0032(.A1(new_n217), .A2(new_n218), .A3(new_n229), .A4(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT68), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT69), .B(G50), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT70), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n220), .A2(new_n222), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT73), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT73), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n220), .A2(new_n222), .A3(new_n257), .A4(new_n254), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G58), .A2(G68), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n225), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G150), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n225), .A2(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n259), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G20), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n268), .B1(G50), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n256), .A2(new_n258), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n271), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n225), .A2(G1), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n274), .A2(new_n261), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g0077(.A(new_n277), .B(KEYINPUT9), .Z(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n284), .A2(G223), .B1(G77), .B2(new_n282), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n282), .A2(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G222), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n285), .A2(KEYINPUT71), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT71), .B1(new_n285), .B2(new_n287), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n223), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT72), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT72), .B1(new_n223), .B2(new_n290), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OR3_X1    g0095(.A1(new_n288), .A2(new_n289), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G274), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  AOI21_X1  g0100(.A(G1), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n297), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n305), .B2(G226), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G190), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(G200), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n278), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n305), .A2(KEYINPUT76), .ZN(new_n315));
  INV_X1    g0115(.A(G238), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT76), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n316), .B1(new_n304), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n303), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n284), .A2(KEYINPUT75), .A3(G232), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT3), .ZN(new_n322));
  INV_X1    g0122(.A(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n279), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n321), .B1(new_n326), .B2(new_n236), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n286), .A2(G226), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  AND4_X1   g0129(.A1(new_n320), .A2(new_n327), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n319), .B1(new_n330), .B2(new_n295), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT13), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n331), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G190), .ZN(new_n336));
  INV_X1    g0136(.A(G68), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G77), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n266), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n259), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(KEYINPUT77), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT11), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(KEYINPUT77), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n346));
  INV_X1    g0146(.A(new_n271), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n337), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT12), .ZN(new_n349));
  OAI21_X1  g0149(.A(G68), .B1(new_n225), .B2(G1), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n274), .B2(new_n350), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n345), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n333), .A2(new_n336), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n352), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT14), .B1(new_n335), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n335), .A2(G179), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n332), .A2(new_n359), .A3(G169), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n354), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n307), .A2(G179), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n277), .B(new_n363), .C1(new_n356), .C2(new_n307), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n303), .ZN(new_n366));
  INV_X1    g0166(.A(G244), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n304), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT74), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n286), .A2(G232), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n284), .A2(G238), .B1(G107), .B2(new_n282), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n295), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G190), .ZN(new_n374));
  INV_X1    g0174(.A(new_n265), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n266), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n259), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G77), .B2(new_n271), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n274), .A2(new_n339), .A3(new_n275), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n374), .B(new_n382), .C1(new_n383), .C2(new_n373), .ZN(new_n384));
  INV_X1    g0184(.A(G179), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n373), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n382), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n356), .B1(new_n369), .B2(new_n372), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n314), .A2(new_n362), .A3(new_n365), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n323), .A2(KEYINPUT78), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT78), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G33), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n322), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(G223), .B(new_n283), .C1(new_n395), .C2(new_n281), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT80), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT78), .B(G33), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n324), .B1(new_n398), .B2(new_n322), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT80), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(G223), .A4(new_n283), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(G226), .A3(G1698), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n397), .A2(new_n401), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n291), .B(new_n292), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n366), .B1(new_n236), .B2(new_n304), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(G200), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AOI211_X1 g0209(.A(G190), .B(new_n407), .C1(new_n404), .C2(new_n405), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n274), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n265), .A2(new_n275), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n412), .A2(new_n413), .B1(new_n347), .B2(new_n265), .ZN(new_n414));
  INV_X1    g0214(.A(G58), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n337), .ZN(new_n416));
  OAI21_X1  g0216(.A(G20), .B1(new_n416), .B2(new_n260), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n263), .A2(G159), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(G20), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n399), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT79), .B1(new_n395), .B2(new_n281), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT79), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n324), .C1(new_n398), .C2(new_n322), .ZN(new_n430));
  AOI21_X1  g0230(.A(G20), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n427), .B1(new_n431), .B2(KEYINPUT7), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n422), .B1(new_n432), .B2(G68), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n392), .A2(new_n394), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n424), .B(new_n279), .C1(new_n434), .C2(KEYINPUT3), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n423), .B1(new_n325), .B2(G20), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n419), .B1(new_n437), .B2(G68), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n259), .B1(new_n438), .B2(KEYINPUT16), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n414), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n411), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n414), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n432), .A2(G68), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n421), .ZN(new_n448));
  INV_X1    g0248(.A(new_n439), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G190), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n406), .A2(new_n451), .A3(new_n408), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n407), .B1(new_n404), .B2(new_n405), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(G200), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n445), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT82), .B1(new_n443), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n406), .A2(G179), .A3(new_n408), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n356), .B2(new_n453), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n458), .A2(new_n459), .A3(new_n440), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(new_n458), .B2(new_n440), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n444), .B1(new_n411), .B2(new_n440), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n450), .A2(new_n454), .A3(new_n441), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n456), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n399), .A2(G257), .A3(new_n283), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n399), .A2(G264), .A3(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n282), .A2(G303), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n405), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n300), .A2(G1), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(G274), .A3(new_n297), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n297), .ZN(new_n477));
  INV_X1    g0277(.A(G270), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n225), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT83), .B(G97), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(new_n323), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n255), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n482), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n225), .B(new_n483), .C1(new_n485), .C2(G33), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(KEYINPUT20), .A3(new_n255), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G1), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G33), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n273), .A2(G116), .A3(new_n271), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n270), .A2(G20), .A3(new_n488), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n481), .A2(new_n499), .A3(KEYINPUT21), .A4(G169), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n479), .B1(new_n471), .B2(new_n405), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n501), .A3(G179), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n501), .A2(new_n356), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT21), .B1(new_n505), .B2(new_n499), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n499), .B1(new_n481), .B2(G200), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n451), .B2(new_n481), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n399), .A2(new_n225), .A3(G68), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n225), .B1(new_n329), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n485), .A2(new_n203), .ZN(new_n514));
  XNOR2_X1  g0314(.A(KEYINPUT86), .B(G87), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n512), .B1(new_n485), .B2(new_n266), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n511), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(new_n259), .B1(new_n347), .B2(new_n377), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n273), .A2(G87), .A3(new_n271), .A4(new_n496), .ZN(new_n520));
  INV_X1    g0320(.A(new_n474), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n521), .A2(G250), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n297), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n298), .B2(new_n521), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n399), .A2(G244), .A3(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n399), .A2(G238), .A3(new_n283), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n398), .A2(new_n488), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n524), .B1(new_n529), .B2(new_n405), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n519), .B(new_n520), .C1(new_n531), .C2(new_n451), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n530), .A2(new_n383), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n518), .A2(new_n259), .ZN(new_n534));
  INV_X1    g0334(.A(new_n377), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n273), .A2(new_n271), .A3(new_n535), .A4(new_n496), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n347), .A2(new_n377), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n531), .B2(G179), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n530), .A2(G169), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n532), .A2(new_n533), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n510), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n476), .A2(G264), .A3(new_n297), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n399), .A2(G257), .A3(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n399), .A2(G250), .A3(new_n283), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n434), .A2(G294), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(new_n405), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n475), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n383), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n405), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT87), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT87), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(new_n553), .A3(new_n405), .ZN(new_n554));
  INV_X1    g0354(.A(new_n475), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n543), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n552), .A2(new_n451), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n412), .A2(G107), .A3(new_n496), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n271), .A2(G107), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n560), .B(KEYINPUT25), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n399), .A2(KEYINPUT22), .A3(new_n225), .A4(G87), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n225), .B2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n527), .A2(new_n225), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n225), .A2(G87), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n282), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n563), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT24), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n562), .B1(new_n572), .B2(new_n259), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n558), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n259), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n559), .A2(new_n561), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n556), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n551), .B2(KEYINPUT87), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n356), .B1(new_n581), .B2(new_n554), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n549), .A2(new_n385), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n263), .A2(G77), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n203), .A2(KEYINPUT6), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n485), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G97), .A2(G107), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT6), .B1(new_n204), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n586), .B1(new_n591), .B2(new_n225), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n203), .B1(new_n435), .B2(new_n436), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n259), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n273), .A2(G97), .A3(new_n271), .A4(new_n496), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n347), .A2(new_n202), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n477), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n555), .B1(new_n598), .B2(G257), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT4), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n600), .A2(new_n367), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(new_n283), .C1(new_n280), .C2(new_n281), .ZN(new_n602));
  OAI211_X1 g0402(.A(G250), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n483), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G244), .B(new_n283), .C1(new_n395), .C2(new_n281), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n599), .B1(new_n606), .B2(new_n295), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n599), .B(KEYINPUT84), .C1(new_n606), .C2(new_n295), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n597), .B1(new_n611), .B2(new_n356), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n599), .B(new_n385), .C1(new_n606), .C2(new_n295), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(G200), .B2(new_n607), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n609), .A2(G190), .A3(new_n610), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n612), .A2(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n542), .A2(new_n585), .A3(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n391), .A2(new_n467), .A3(new_n620), .ZN(G372));
  NOR2_X1   g0421(.A1(new_n391), .A2(new_n467), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n503), .A2(new_n506), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n584), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n385), .A2(new_n530), .B1(new_n519), .B2(new_n536), .ZN(new_n625));
  INV_X1    g0425(.A(new_n524), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT88), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n529), .A2(new_n405), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n529), .B2(new_n405), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n356), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(G200), .ZN(new_n632));
  AOI211_X1 g0432(.A(new_n451), .B(new_n524), .C1(new_n529), .C2(new_n405), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n519), .A2(new_n520), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n625), .A2(new_n631), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n624), .A2(new_n619), .A3(new_n574), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n629), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n529), .A2(new_n405), .A3(new_n627), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n524), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n625), .B1(new_n640), .B2(G169), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT89), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n612), .A2(new_n615), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT26), .B1(new_n643), .B2(new_n636), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n612), .A2(new_n615), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n645), .A2(new_n541), .A3(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n637), .B(new_n642), .C1(new_n644), .C2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n622), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n462), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n361), .A2(new_n355), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n354), .B1(new_n651), .B2(new_n389), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n456), .A2(new_n466), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n314), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n365), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n649), .A2(new_n656), .ZN(G369));
  NAND2_X1  g0457(.A1(new_n270), .A2(new_n225), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT90), .Z(new_n660));
  OAI21_X1  g0460(.A(G213), .B1(new_n658), .B2(KEYINPUT27), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n499), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT91), .Z(new_n666));
  INV_X1    g0466(.A(new_n623), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n510), .B2(new_n666), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n664), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n585), .B1(new_n573), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n584), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n585), .A2(new_n667), .A3(new_n671), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n584), .A2(new_n664), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n230), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G1), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n514), .A2(new_n515), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n488), .ZN(new_n685));
  OAI22_X1  g0485(.A1(new_n683), .A2(new_n685), .B1(new_n227), .B2(new_n682), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n542), .A2(new_n585), .A3(new_n619), .A4(new_n671), .ZN(new_n689));
  AND4_X1   g0489(.A1(new_n385), .A2(new_n549), .A3(new_n481), .A4(new_n607), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n501), .A2(new_n548), .A3(new_n530), .A4(G179), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n611), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n630), .A2(new_n690), .B1(new_n692), .B2(KEYINPUT30), .ZN(new_n693));
  AND4_X1   g0493(.A1(G179), .A2(new_n501), .A3(new_n548), .A4(new_n530), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(KEYINPUT92), .A3(new_n609), .A4(new_n610), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n611), .B2(new_n691), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n671), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n689), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n690), .A2(new_n630), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n548), .A2(new_n530), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n501), .A2(G179), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n609), .A4(new_n610), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n705), .B1(new_n708), .B2(new_n696), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n699), .A2(KEYINPUT93), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT93), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n695), .A2(new_n711), .A3(new_n698), .A4(new_n696), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n709), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n701), .B1(new_n713), .B2(new_n671), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT94), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n704), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT30), .B1(new_n708), .B2(new_n697), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n711), .B1(new_n717), .B2(new_n695), .ZN(new_n718));
  INV_X1    g0518(.A(new_n712), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n693), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n720), .B2(new_n664), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT94), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n688), .B1(new_n716), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT29), .B1(new_n648), .B2(new_n671), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n632), .A2(new_n635), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n641), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT26), .B1(new_n726), .B2(new_n645), .ZN(new_n727));
  INV_X1    g0527(.A(new_n541), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n643), .A2(new_n728), .A3(new_n646), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n727), .A2(new_n729), .A3(new_n642), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT95), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n617), .A2(new_n618), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n643), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n636), .A2(new_n574), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n619), .A2(KEYINPUT95), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n733), .A2(new_n734), .A3(new_n624), .A4(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n664), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n724), .B1(KEYINPUT29), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n723), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n687), .B1(new_n739), .B2(G1), .ZN(G364));
  NOR2_X1   g0540(.A1(new_n269), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n495), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n681), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n670), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G330), .B2(new_n669), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n224), .B1(G20), .B2(new_n356), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n225), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n385), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n339), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n225), .B1(new_n756), .B2(G190), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT98), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G97), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n225), .A2(new_n451), .A3(new_n383), .A4(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n760), .A2(new_n515), .B1(G68), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n761), .A2(new_n451), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n759), .B(new_n763), .C1(new_n261), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n750), .A2(G20), .A3(G190), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n225), .A2(new_n383), .A3(G179), .A4(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n325), .B1(new_n415), .B2(new_n767), .C1(new_n769), .C2(new_n203), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n749), .A2(new_n756), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n773), .B(new_n774), .ZN(new_n775));
  OR4_X1    g0575(.A1(new_n755), .A2(new_n766), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n767), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n282), .B1(new_n751), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n771), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n778), .B(new_n780), .C1(G329), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n764), .A2(G326), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n760), .A2(G303), .B1(new_n762), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n757), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G294), .B1(new_n768), .B2(G283), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n782), .A2(new_n783), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n748), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n747), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n228), .A2(new_n300), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n428), .A2(new_n430), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n680), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n795), .B(new_n798), .C1(new_n248), .C2(new_n300), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n680), .A2(new_n282), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G355), .B1(new_n488), .B2(new_n680), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n794), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n744), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n789), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n792), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n669), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n746), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NOR2_X1   g0608(.A1(new_n747), .A2(new_n790), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n803), .B1(new_n809), .B2(new_n339), .ZN(new_n810));
  INV_X1    g0610(.A(new_n754), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G116), .ZN(new_n812));
  INV_X1    g0612(.A(new_n760), .ZN(new_n813));
  INV_X1    g0613(.A(G303), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n203), .B1(new_n814), .B2(new_n765), .ZN(new_n815));
  INV_X1    g0615(.A(G87), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  INV_X1    g0617(.A(new_n762), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n769), .A2(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n282), .B1(new_n771), .B2(new_n779), .ZN(new_n821));
  INV_X1    g0621(.A(new_n767), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(G294), .B2(new_n822), .ZN(new_n823));
  AND4_X1   g0623(.A1(new_n759), .A2(new_n812), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n822), .A2(G143), .B1(G137), .B2(new_n764), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n826), .B2(new_n818), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G159), .B2(new_n811), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n769), .A2(new_n337), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G50), .B2(new_n760), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G132), .A2(new_n781), .B1(new_n786), .B2(G58), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n831), .A2(new_n797), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n828), .B2(KEYINPUT34), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n824), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n389), .A2(new_n664), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n384), .B1(new_n382), .B2(new_n671), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n389), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n810), .B1(new_n748), .B2(new_n835), .C1(new_n838), .C2(new_n791), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n648), .A2(new_n671), .A3(new_n838), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT99), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n648), .A2(KEYINPUT99), .A3(new_n671), .A4(new_n838), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n648), .A2(new_n671), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n838), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n716), .A2(new_n722), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(G330), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n803), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n846), .A2(new_n848), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n839), .B1(new_n850), .B2(new_n851), .ZN(G384));
  INV_X1    g0652(.A(new_n591), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n226), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OAI211_X1 g0657(.A(new_n228), .B(G77), .C1(new_n415), .C2(new_n337), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n261), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n495), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n741), .A2(new_n495), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n450), .A2(new_n454), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n447), .A2(new_n417), .A3(new_n418), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n420), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n433), .A2(new_n273), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n446), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n458), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n662), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n662), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n440), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n863), .B(new_n873), .C1(new_n868), .C2(new_n450), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n871), .B1(KEYINPUT37), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT100), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n467), .A2(new_n876), .A3(new_n870), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n467), .B2(new_n870), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT38), .B(new_n875), .C1(new_n877), .C2(new_n878), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n874), .B(KEYINPUT37), .Z(new_n884));
  NOR2_X1   g0684(.A1(new_n443), .A2(new_n455), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n873), .B1(new_n885), .B2(new_n462), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n880), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n361), .A2(new_n355), .A3(new_n671), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n355), .A2(new_n664), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n651), .A2(new_n353), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n355), .B(new_n664), .C1(new_n354), .C2(new_n361), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n836), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n844), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT101), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n881), .A2(new_n901), .A3(new_n882), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n881), .B2(new_n882), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n898), .B(new_n900), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n650), .A2(new_n662), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n894), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n656), .B1(new_n738), .B2(new_n622), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n906), .B(new_n907), .Z(new_n908));
  NAND2_X1  g0708(.A1(new_n898), .A2(new_n838), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT102), .ZN(new_n910));
  INV_X1    g0710(.A(new_n702), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n689), .B1(new_n713), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(new_n721), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n720), .A2(new_n702), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n714), .A2(new_n914), .A3(KEYINPUT102), .A4(new_n689), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n909), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(KEYINPUT40), .A3(new_n888), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n916), .B1(new_n902), .B2(new_n903), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n913), .A2(new_n915), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n622), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(G330), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n921), .B1(new_n622), .B2(new_n922), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n862), .B1(new_n908), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n927), .A2(new_n928), .B1(new_n908), .B2(new_n926), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n861), .B1(new_n929), .B2(new_n930), .ZN(G367));
  NAND2_X1  g0731(.A1(new_n664), .A2(new_n634), .ZN(new_n932));
  MUX2_X1   g0732(.A(new_n642), .B(new_n726), .S(new_n932), .Z(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n792), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n822), .A2(G303), .B1(new_n781), .B2(G317), .ZN(new_n935));
  INV_X1    g0735(.A(G294), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n936), .B2(new_n818), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G283), .B2(new_n811), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n769), .A2(new_n485), .B1(new_n779), .B2(new_n765), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G107), .B2(new_n786), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT46), .B1(new_n813), .B2(new_n488), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n813), .A2(KEYINPUT46), .A3(new_n488), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n797), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT110), .ZN(new_n945));
  INV_X1    g0745(.A(new_n758), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(new_n337), .ZN(new_n947));
  INV_X1    g0747(.A(G143), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n818), .A2(new_n772), .B1(new_n765), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n769), .A2(new_n339), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(G58), .C2(new_n760), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n767), .A2(new_n826), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n282), .B(new_n952), .C1(G137), .C2(new_n781), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(new_n261), .C2(new_n754), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n945), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT47), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n747), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n798), .A2(new_n242), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n958), .B(new_n793), .C1(new_n230), .C2(new_n377), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n934), .A2(new_n957), .A3(new_n744), .A4(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n933), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n664), .A2(new_n616), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n733), .A2(new_n735), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n643), .A2(new_n664), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n675), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT105), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(KEYINPUT105), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT42), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n967), .A2(KEYINPUT105), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT42), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n968), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n645), .B1(new_n964), .B2(new_n584), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n671), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT104), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n933), .A2(new_n961), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n977), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n962), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n977), .A2(new_n979), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT104), .ZN(new_n984));
  INV_X1    g0784(.A(new_n962), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n674), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n966), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n982), .A2(new_n987), .B1(KEYINPUT106), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n681), .B(KEYINPUT41), .Z(new_n992));
  INV_X1    g0792(.A(new_n675), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n667), .A2(new_n671), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n993), .B1(new_n673), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n670), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT109), .B1(new_n739), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n739), .A2(KEYINPUT109), .A3(new_n997), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n966), .A2(new_n678), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1001), .B1(new_n966), .B2(new_n678), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n966), .A2(new_n678), .ZN(new_n1006));
  XOR2_X1   g0806(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1008), .A3(new_n674), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n988), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n999), .A2(new_n1000), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n992), .B1(new_n1012), .B2(new_n739), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n990), .A2(new_n991), .B1(new_n743), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n982), .A2(new_n987), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n991), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n960), .B1(new_n1014), .B2(new_n1019), .ZN(G387));
  AND3_X1   g0820(.A1(new_n739), .A2(KEYINPUT109), .A3(new_n997), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n998), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1022), .A2(KEYINPUT115), .A3(new_n682), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT115), .B1(new_n1022), .B2(new_n682), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n739), .C2(new_n997), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n997), .A2(new_n743), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT111), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n673), .A2(new_n805), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n798), .B1(new_n239), .B2(new_n300), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n685), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n800), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1033));
  OR3_X1    g0833(.A1(new_n265), .A2(new_n1033), .A3(G50), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n265), .B2(G50), .ZN(new_n1035));
  AOI21_X1  g0835(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1030), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1032), .A2(new_n1037), .B1(new_n203), .B2(new_n680), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n744), .B1(new_n1038), .B2(new_n794), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n751), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1040), .A2(G68), .B1(new_n781), .B2(G150), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n261), .B2(new_n767), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n813), .A2(new_n339), .B1(new_n772), .B2(new_n765), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n769), .A2(new_n202), .B1(new_n265), .B2(new_n818), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n758), .A2(new_n535), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n797), .A3(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n813), .A2(new_n936), .B1(new_n817), .B2(new_n757), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n822), .A2(G317), .B1(G311), .B2(new_n762), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n777), .B2(new_n765), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G303), .B2(new_n811), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1048), .B1(new_n1051), .B2(KEYINPUT48), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT113), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(KEYINPUT48), .B2(new_n1051), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n781), .A2(G326), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n796), .B(new_n1057), .C1(new_n488), .C2(new_n769), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT114), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1047), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1039), .B1(new_n1061), .B2(new_n747), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1027), .B1(new_n1028), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1025), .A2(new_n1063), .ZN(G393));
  INV_X1    g0864(.A(KEYINPUT117), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1011), .A2(new_n743), .A3(new_n1009), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n822), .A2(G311), .B1(G317), .B2(new_n764), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n282), .B1(new_n771), .B2(new_n777), .C1(new_n936), .C2(new_n751), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n769), .A2(new_n203), .B1(new_n814), .B2(new_n818), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n813), .A2(new_n817), .B1(new_n488), .B2(new_n757), .ZN(new_n1071));
  OR4_X1    g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n769), .A2(new_n816), .B1(new_n948), .B2(new_n771), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n813), .A2(new_n337), .B1(new_n261), .B2(new_n818), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n811), .C2(new_n375), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n758), .A2(G77), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n765), .A2(new_n826), .B1(new_n767), .B2(new_n772), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n797), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n748), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n793), .B1(new_n230), .B2(new_n485), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n252), .B2(new_n798), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1080), .A2(new_n803), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n966), .B2(new_n805), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1066), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT116), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1066), .B2(new_n1084), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1011), .A2(new_n1009), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1021), .B2(new_n998), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1012), .A2(new_n1091), .A3(new_n681), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1065), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(KEYINPUT117), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(G390));
  AOI211_X1 g0896(.A(new_n688), .B(new_n909), .C1(new_n913), .C2(new_n915), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n900), .A2(new_n898), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1098), .A2(new_n892), .B1(new_n883), .B2(new_n890), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n837), .A2(new_n389), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n737), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n899), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n893), .B1(new_n1102), .B2(new_n898), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n888), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1097), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n922), .A2(G330), .A3(new_n622), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n907), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n898), .B1(new_n723), .B2(new_n838), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n900), .B1(new_n1109), .B2(new_n1097), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1102), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n847), .A2(G330), .A3(new_n838), .A4(new_n898), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n838), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n688), .B(new_n1113), .C1(new_n913), .C2(new_n915), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1111), .B(new_n1112), .C1(new_n1114), .C2(new_n898), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1108), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n893), .B1(new_n900), .B2(new_n898), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1104), .B(new_n1112), .C1(new_n891), .C2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1106), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT118), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT118), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1106), .A2(new_n1116), .A3(new_n1121), .A4(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1106), .A2(new_n1118), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1116), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n682), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n803), .B1(new_n809), .B2(new_n265), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT119), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n813), .A2(new_n816), .B1(new_n203), .B2(new_n818), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n830), .B(new_n1130), .C1(G283), .C2(new_n764), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n811), .A2(new_n486), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n282), .B1(new_n771), .B2(new_n936), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G116), .B2(new_n822), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1131), .A2(new_n1076), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n811), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G132), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n325), .B1(new_n767), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G125), .B2(new_n781), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n813), .A2(KEYINPUT53), .A3(new_n826), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT53), .B1(new_n813), .B2(new_n826), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1138), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n762), .A2(G137), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n768), .A2(G50), .B1(G128), .B2(new_n764), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n946), .C2(new_n772), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1135), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1129), .B1(new_n1148), .B2(new_n747), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n891), .B2(new_n791), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1124), .B2(new_n742), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1127), .A2(new_n1151), .ZN(G378));
  AOI21_X1  g0952(.A(new_n803), .B1(new_n809), .B2(new_n261), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n760), .A2(new_n1137), .B1(G125), .B2(new_n764), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n822), .A2(G128), .B1(new_n1040), .B2(G137), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n1139), .C2(new_n818), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G150), .B2(new_n758), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n768), .A2(G159), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G33), .B(G41), .C1(new_n781), .C2(G124), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(G41), .B1(new_n781), .B2(G283), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n203), .B2(new_n767), .C1(new_n377), .C2(new_n751), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n760), .A2(G77), .B1(G116), .B2(new_n764), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n768), .A2(G58), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n202), .C2(new_n818), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n947), .A2(new_n1165), .A3(new_n1168), .A4(new_n797), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT58), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT58), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n299), .B1(new_n796), .B2(new_n323), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n261), .ZN(new_n1173));
  AND4_X1   g0973(.A1(new_n1163), .A2(new_n1170), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n314), .A2(new_n365), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n277), .A2(new_n662), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1153), .B1(new_n748), .B2(new_n1174), .C1(new_n1180), .C2(new_n791), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n906), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1180), .B1(new_n921), .B2(G330), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n916), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n467), .A2(new_n870), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT100), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n467), .A2(new_n876), .A3(new_n870), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT38), .B1(new_n1189), .B2(new_n875), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n882), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT101), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n881), .A2(new_n901), .A3(new_n882), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1185), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(G330), .B(new_n917), .C1(new_n1194), .C2(KEYINPUT40), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(new_n1179), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1183), .B1(new_n1184), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1179), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n919), .A2(new_n920), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1199), .A2(G330), .A3(new_n917), .A4(new_n1180), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1200), .A3(new_n906), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1197), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1182), .B1(new_n1202), .B2(new_n743), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1108), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1198), .A2(new_n906), .A3(new_n1200), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n906), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT120), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT120), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1201), .A2(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1204), .B(new_n1205), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1108), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1123), .A2(new_n1212), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n681), .B1(new_n1213), .B2(KEYINPUT57), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1203), .B1(new_n1211), .B2(new_n1214), .ZN(G375));
  AND2_X1   g1015(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1108), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1218), .A2(new_n992), .A3(new_n1116), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n813), .A2(new_n202), .B1(new_n936), .B2(new_n765), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n950), .B(new_n1220), .C1(G116), .C2(new_n762), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n811), .A2(G107), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n282), .B1(new_n771), .B2(new_n814), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G283), .B2(new_n822), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1221), .A2(new_n1046), .A3(new_n1222), .A4(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n758), .A2(G50), .B1(G150), .B2(new_n1040), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT121), .Z(new_n1227));
  OAI22_X1  g1027(.A1(new_n1139), .A2(new_n765), .B1(new_n818), .B2(new_n1136), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G159), .B2(new_n760), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n822), .A2(G137), .B1(new_n781), .B2(G128), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n797), .A3(new_n1167), .A4(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1225), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n747), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n803), .B1(new_n809), .B2(new_n337), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n898), .C2(new_n791), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1216), .B2(new_n742), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1219), .A2(new_n1236), .ZN(G381));
  NAND3_X1  g1037(.A1(new_n1025), .A2(new_n807), .A3(new_n1063), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1238), .ZN(new_n1239));
  OR4_X1    g1039(.A1(G387), .A2(new_n1239), .A3(G375), .A4(G378), .ZN(G407));
  NOR2_X1   g1040(.A1(new_n1127), .A2(new_n1151), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n663), .A2(G213), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G407), .B(G213), .C1(G375), .C2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT122), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1245), .B(new_n1246), .ZN(G409));
  OAI211_X1 g1047(.A(G378), .B(new_n1203), .C1(new_n1211), .C2(new_n1214), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1123), .A2(new_n1212), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1202), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1181), .B1(new_n1250), .B2(new_n992), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n742), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1241), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1243), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1217), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n681), .B1(new_n1255), .B2(new_n1217), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(new_n1236), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  XOR2_X1   g1062(.A(G384), .B(KEYINPUT124), .Z(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1259), .B2(new_n1236), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1254), .A2(KEYINPUT63), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G393), .A2(G396), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1238), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G387), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n990), .A2(new_n991), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1013), .A2(new_n743), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G390), .B1(new_n1276), .B2(new_n960), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1270), .B1(new_n1272), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(new_n1271), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1276), .A2(G390), .A3(new_n960), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1238), .A3(new_n1269), .A4(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1268), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT123), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1248), .A2(new_n1253), .A3(KEYINPUT123), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1290), .A2(new_n1242), .A3(new_n1267), .A4(new_n1291), .ZN(new_n1292));
  XOR2_X1   g1092(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1290), .A2(new_n1242), .A3(new_n1291), .ZN(new_n1295));
  INV_X1    g1095(.A(G2897), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1267), .B1(new_n1296), .B2(new_n1242), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1266), .A2(G2897), .A3(new_n1243), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1295), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1287), .A2(new_n1294), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1279), .B1(new_n1301), .B2(new_n1254), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1292), .A2(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1266), .A2(new_n1303), .ZN(new_n1305));
  AND4_X1   g1105(.A1(KEYINPUT127), .A2(new_n1288), .A3(new_n1242), .A4(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT127), .B1(new_n1254), .B2(new_n1305), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1302), .B1(new_n1304), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1300), .B1(new_n1309), .B2(new_n1311), .ZN(G405));
  XNOR2_X1  g1112(.A(G375), .B(G378), .ZN(new_n1313));
  OR2_X1    g1113(.A1(new_n1313), .A2(new_n1266), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1266), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1310), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1314), .A2(new_n1311), .A3(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


