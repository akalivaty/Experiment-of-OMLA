//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1295, new_n1296,
    new_n1297, new_n1299, new_n1300, new_n1301, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374, new_n1375;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n210), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT8), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT8), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n211), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(new_n256), .B1(G150), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n203), .A2(G20), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n249), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n249), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G50), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n263), .A2(new_n265), .B1(G50), .B2(new_n262), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT65), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(KEYINPUT65), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G77), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n271), .A2(new_n276), .A3(G222), .A4(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n271), .A2(new_n276), .A3(G223), .A4(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n278), .A2(new_n284), .A3(new_n280), .A4(new_n281), .ZN(new_n285));
  AND2_X1   g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n210), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n283), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT64), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n286), .B2(new_n210), .ZN(new_n290));
  AND2_X1   g0090(.A1(G1), .A2(G13), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(KEYINPUT64), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n290), .A2(new_n293), .A3(G274), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n290), .A2(new_n293), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n295), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(G226), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n267), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  INV_X1    g0104(.A(new_n300), .ZN(new_n305));
  INV_X1    g0105(.A(new_n287), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n282), .B2(KEYINPUT66), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n307), .B2(new_n285), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n303), .A2(KEYINPUT67), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(KEYINPUT67), .B2(new_n303), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n217), .A2(G20), .ZN(new_n311));
  INV_X1    g0111(.A(new_n257), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n255), .B2(new_n223), .C1(new_n312), .C2(new_n202), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n248), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT11), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n262), .A2(KEYINPUT70), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n317), .A2(new_n261), .A3(G13), .A4(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT12), .B1(new_n319), .B2(G68), .ZN(new_n320));
  INV_X1    g0120(.A(G13), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G1), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(KEYINPUT12), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n320), .B1(new_n311), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n248), .B1(new_n316), .B2(new_n318), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G68), .A3(new_n264), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n315), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G226), .A2(G1698), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n232), .B2(G1698), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n271), .A2(new_n330), .A3(new_n276), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G97), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n287), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n290), .A2(new_n293), .A3(G238), .A4(new_n294), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n296), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n306), .B1(new_n331), .B2(new_n332), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n296), .A2(new_n336), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT13), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(G169), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(G179), .A3(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n342), .B2(G169), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n328), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n328), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n342), .A2(G200), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n349), .B(new_n350), .C1(new_n351), .C2(new_n342), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n254), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT69), .B1(new_n354), .B2(new_n255), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n354), .A2(KEYINPUT69), .A3(new_n255), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n248), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n319), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n223), .B1(new_n261), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n359), .A2(new_n223), .B1(new_n326), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n297), .B1(G244), .B2(new_n299), .ZN(new_n363));
  NOR2_X1   g0163(.A1(G232), .A2(G1698), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n218), .B2(G1698), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n277), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n277), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT68), .B(G107), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n287), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n363), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n362), .B1(new_n302), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(G179), .B2(new_n370), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(G200), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n362), .C1(new_n351), .C2(new_n370), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n352), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n310), .A2(new_n348), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n288), .A2(G190), .A3(new_n300), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n267), .A2(KEYINPUT9), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n260), .B2(new_n266), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n377), .B(new_n382), .C1(new_n308), .C2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n377), .A2(new_n382), .A3(KEYINPUT71), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT10), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n381), .B1(new_n308), .B2(G190), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n301), .A2(G200), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n388), .B(new_n389), .C1(KEYINPUT71), .C2(KEYINPUT10), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G41), .A2(G45), .ZN(new_n393));
  OAI21_X1  g0193(.A(G232), .B1(new_n393), .B2(G1), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n261), .B(G274), .C1(G41), .C2(G45), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT74), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n396), .A2(new_n298), .A3(new_n397), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n286), .A2(new_n289), .A3(new_n210), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT64), .B1(new_n291), .B2(new_n292), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n394), .A2(new_n395), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT74), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  OR2_X1    g0205(.A1(G223), .A2(G1698), .ZN(new_n406));
  INV_X1    g0206(.A(G226), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n269), .A2(new_n270), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(G179), .B1(new_n411), .B2(new_n287), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n392), .B1(new_n404), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n397), .B1(new_n396), .B2(new_n298), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n401), .A2(KEYINPUT74), .A3(new_n402), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n412), .A2(new_n414), .A3(new_n392), .A4(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n396), .A2(new_n298), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n274), .A2(new_n275), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n406), .A3(new_n408), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n306), .B1(new_n419), .B2(new_n405), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n302), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT76), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT75), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT76), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n421), .A4(new_n416), .ZN(new_n427));
  INV_X1    g0227(.A(new_n263), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n254), .A2(new_n264), .ZN(new_n429));
  INV_X1    g0229(.A(new_n254), .ZN(new_n430));
  INV_X1    g0230(.A(new_n262), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n428), .A2(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT7), .B1(new_n277), .B2(new_n211), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n275), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT73), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT73), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n410), .A2(new_n437), .A3(KEYINPUT7), .A4(new_n211), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n250), .A2(new_n217), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n441), .A2(new_n201), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(G20), .B1(G159), .B2(new_n257), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n433), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT7), .B1(new_n410), .B2(new_n211), .ZN(new_n445));
  INV_X1    g0245(.A(new_n435), .ZN(new_n446));
  OAI21_X1  g0246(.A(G68), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(KEYINPUT16), .A3(new_n443), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n248), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n432), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n423), .A2(new_n427), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT18), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n423), .A2(new_n450), .A3(new_n453), .A4(new_n427), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n411), .A2(new_n287), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n414), .A2(new_n415), .A3(new_n455), .A4(new_n351), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n383), .B1(new_n417), .B2(new_n420), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n432), .C1(new_n444), .C2(new_n449), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT17), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT17), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n452), .A2(new_n454), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n376), .A2(new_n391), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(new_n290), .A3(G270), .A4(new_n293), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n261), .A2(G45), .A3(G274), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n290), .A2(new_n293), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT78), .A2(G303), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT78), .A2(G303), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n271), .B2(new_n276), .ZN(new_n480));
  INV_X1    g0280(.A(G257), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n279), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n226), .A2(G1698), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(new_n483), .C1(new_n269), .C2(new_n270), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n287), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n302), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n261), .A2(G33), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n319), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G116), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n326), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n247), .A2(new_n210), .B1(G20), .B2(new_n491), .ZN(new_n493));
  AOI21_X1  g0293(.A(G20), .B1(G33), .B2(G283), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(G33), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT79), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n492), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n492), .B2(new_n501), .ZN(new_n504));
  OAI211_X1 g0304(.A(KEYINPUT21), .B(new_n487), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n476), .A2(new_n486), .A3(G179), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n503), .B2(new_n504), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n319), .A2(new_n249), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(G116), .B1(new_n319), .B2(new_n489), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT20), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT20), .B1(new_n493), .B2(new_n496), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT79), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n492), .A2(new_n501), .A3(new_n502), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT21), .B1(new_n516), .B2(new_n487), .ZN(new_n517));
  INV_X1    g0317(.A(new_n479), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n277), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n306), .B1(new_n519), .B2(new_n484), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n471), .A2(new_n475), .ZN(new_n521));
  OAI21_X1  g0321(.A(G200), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n476), .A2(new_n486), .A3(G190), .ZN(new_n523));
  AND4_X1   g0323(.A1(new_n515), .A2(new_n522), .A3(new_n514), .A4(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n508), .A2(new_n517), .A3(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n470), .A2(new_n290), .A3(G257), .A4(new_n293), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n475), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(new_n279), .C1(new_n269), .C2(new_n270), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n529), .B1(G33), .B2(G283), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n224), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n271), .A2(new_n276), .A3(new_n279), .A4(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n271), .A2(new_n276), .A3(G250), .A4(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI211_X1 g0334(.A(G179), .B(new_n527), .C1(new_n534), .C2(new_n287), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n368), .B1(new_n434), .B2(new_n439), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n537), .A2(new_n495), .A3(G107), .ZN(new_n538));
  XNOR2_X1  g0338(.A(G97), .B(G107), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n540), .A2(new_n211), .B1(new_n223), .B2(new_n312), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n248), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n431), .A2(new_n495), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n262), .A2(new_n488), .A3(new_n210), .A4(new_n247), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n495), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n535), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n527), .B1(new_n534), .B2(new_n287), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n302), .ZN(new_n552));
  AOI21_X1  g0352(.A(G20), .B1(new_n271), .B2(new_n276), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n436), .B(new_n438), .C1(new_n553), .C2(KEYINPUT7), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n541), .B1(new_n554), .B2(new_n368), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n548), .B1(new_n555), .B2(new_n249), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(new_n351), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G200), .B2(new_n550), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n549), .A2(new_n552), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n470), .A2(new_n290), .A3(G264), .A4(new_n293), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G250), .A2(G1698), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n481), .B2(G1698), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n418), .B1(G33), .B2(G294), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n475), .B(new_n561), .C1(new_n564), .C2(new_n306), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G169), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT80), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n470), .A2(new_n290), .A3(new_n293), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n481), .A2(G1698), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G250), .B2(G1698), .ZN(new_n570));
  INV_X1    g0370(.A(G294), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n570), .A2(new_n410), .B1(new_n273), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n568), .A2(G264), .B1(new_n572), .B2(new_n287), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(G179), .A3(new_n475), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n573), .A2(KEYINPUT80), .A3(G179), .A4(new_n475), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n219), .A2(KEYINPUT22), .A3(G20), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n271), .A2(new_n276), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n211), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT22), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n225), .A2(G20), .ZN(new_n582));
  OAI22_X1  g0382(.A1(KEYINPUT23), .A2(new_n582), .B1(new_n255), .B2(new_n491), .ZN(new_n583));
  OR2_X1    g0383(.A1(KEYINPUT68), .A2(G107), .ZN(new_n584));
  NAND2_X1  g0384(.A1(KEYINPUT68), .A2(G107), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(G20), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n583), .B1(KEYINPUT23), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT24), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n581), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n581), .B2(new_n587), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n248), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n323), .A2(new_n582), .ZN(new_n592));
  XOR2_X1   g0392(.A(new_n592), .B(KEYINPUT25), .Z(new_n593));
  NOR2_X1   g0393(.A1(new_n546), .A2(new_n225), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n575), .A2(new_n576), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n473), .B1(new_n467), .B2(new_n220), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n290), .A3(new_n293), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT77), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n224), .A2(G1698), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G238), .B2(G1698), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n603), .B2(new_n410), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n287), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n597), .A2(KEYINPUT77), .A3(new_n290), .A4(new_n293), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n302), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n599), .A2(new_n598), .B1(new_n604), .B2(new_n287), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n304), .A3(new_n606), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT19), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n211), .B1(new_n332), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n219), .A2(new_n495), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n368), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n418), .A2(new_n211), .A3(G68), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n255), .B2(new_n495), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n248), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n316), .A2(new_n318), .A3(new_n354), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n546), .A2(new_n354), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n608), .A2(new_n610), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n607), .A2(G200), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n546), .A2(new_n219), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n619), .B(new_n625), .C1(new_n617), .C2(new_n248), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n607), .A2(new_n351), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n565), .A2(new_n383), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n572), .A2(new_n287), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n351), .A3(new_n475), .A4(new_n561), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n591), .A2(new_n595), .A3(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n596), .A2(new_n629), .A3(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n465), .A2(new_n525), .A3(new_n560), .A4(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n535), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n552), .A2(new_n556), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(new_n629), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT83), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n549), .A2(new_n641), .A3(new_n552), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(KEYINPUT83), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n383), .B1(new_n609), .B2(new_n606), .ZN(new_n645));
  INV_X1    g0445(.A(new_n625), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n618), .A2(new_n620), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT81), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n628), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT81), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n624), .A2(new_n626), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n623), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT82), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(KEYINPUT82), .A3(new_n623), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n644), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n640), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n652), .A2(KEYINPUT82), .A3(new_n623), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT82), .B1(new_n652), .B2(new_n623), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n591), .A2(new_n595), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT80), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n565), .B2(G169), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n565), .A2(new_n304), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n576), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n487), .B1(new_n503), .B2(new_n504), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT21), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n667), .A2(new_n670), .A3(new_n507), .A4(new_n505), .ZN(new_n671));
  INV_X1    g0471(.A(new_n634), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n560), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n623), .B1(new_n661), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n658), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n465), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT84), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n391), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n387), .A2(new_n390), .A3(KEYINPUT84), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n459), .B(KEYINPUT17), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n372), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n352), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n685), .B2(new_n348), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n425), .A2(new_n421), .A3(new_n416), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n688), .A2(new_n453), .A3(new_n450), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n453), .B1(new_n688), .B2(new_n450), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n681), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n677), .A2(new_n310), .A3(new_n693), .ZN(G369));
  OR3_X1    g0494(.A1(new_n323), .A2(KEYINPUT27), .A3(G20), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT27), .B1(new_n323), .B2(G20), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n516), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT85), .Z(new_n701));
  NAND3_X1  g0501(.A1(new_n670), .A2(new_n507), .A3(new_n505), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT86), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(KEYINPUT86), .A3(new_n702), .ZN(new_n706));
  INV_X1    g0506(.A(new_n525), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n705), .B(new_n706), .C1(new_n707), .C2(new_n701), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n672), .A2(new_n667), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n662), .ZN(new_n711));
  INV_X1    g0511(.A(new_n699), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n596), .A2(new_n699), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n708), .A2(G330), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n702), .A2(new_n712), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n717), .A2(new_n709), .B1(new_n667), .B2(new_n699), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(G399));
  NOR3_X1   g0520(.A1(new_n368), .A2(G116), .A3(new_n613), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT87), .Z(new_n722));
  INV_X1    g0522(.A(new_n207), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G1), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n722), .A2(new_n726), .B1(new_n215), .B2(new_n725), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n676), .A2(new_n729), .A3(new_n712), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n519), .A2(new_n484), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n521), .B1(new_n731), .B2(new_n287), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n550), .A2(new_n732), .A3(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n573), .A2(new_n609), .A3(KEYINPUT88), .A4(new_n606), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT88), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n631), .A2(new_n561), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n607), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n733), .A2(KEYINPUT30), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(new_n734), .A3(new_n506), .A4(new_n550), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n476), .A2(new_n486), .ZN(new_n742));
  AND4_X1   g0542(.A1(new_n304), .A2(new_n742), .A3(new_n607), .A4(new_n565), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n551), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n738), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n699), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT31), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n635), .A2(new_n525), .A3(new_n560), .A4(new_n712), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT26), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n639), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n623), .B(new_n754), .C1(new_n661), .C2(new_n673), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n655), .A2(new_n656), .ZN(new_n756));
  INV_X1    g0556(.A(new_n644), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n712), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n730), .A2(new_n752), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n728), .B1(new_n762), .B2(G1), .ZN(G364));
  NAND2_X1  g0563(.A1(new_n708), .A2(G330), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n321), .A2(G20), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G45), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT89), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT89), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n768), .A2(G1), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n724), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n708), .ZN(new_n773));
  INV_X1    g0573(.A(new_n771), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n210), .B1(G20), .B2(new_n302), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n211), .A2(G179), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n351), .A3(G200), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT95), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT95), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G107), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n304), .A2(new_n383), .A3(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G97), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n777), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n791));
  NAND3_X1  g0591(.A1(new_n790), .A2(G159), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(new_n790), .B2(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n211), .A2(new_n304), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n795), .A2(new_n351), .A3(new_n383), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n793), .B1(G50), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n783), .A2(new_n787), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n794), .A2(new_n788), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT93), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G77), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n794), .A2(G190), .A3(new_n383), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n277), .B1(G58), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n794), .A2(new_n351), .A3(G200), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n211), .A2(new_n351), .A3(new_n383), .A4(G179), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n810), .A2(G68), .B1(new_n811), .B2(G87), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n805), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n798), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(KEYINPUT33), .A2(G317), .ZN(new_n815));
  AND2_X1   g0615(.A1(KEYINPUT33), .A2(G317), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n810), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n796), .ZN(new_n818));
  INV_X1    g0618(.A(G326), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G303), .B2(new_n811), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n782), .A2(G283), .ZN(new_n822));
  INV_X1    g0622(.A(G322), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n806), .A2(new_n823), .B1(new_n799), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G329), .B2(new_n790), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n367), .B1(G294), .B2(new_n785), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n821), .A2(new_n822), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n776), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G13), .A2(G33), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT92), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(G20), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n277), .A2(new_n723), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(G355), .B1(new_n491), .B2(new_n723), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n245), .A2(G45), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT90), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n723), .A2(new_n418), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(G45), .B2(new_n215), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n834), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT91), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n832), .B(new_n775), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n774), .B(new_n829), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n832), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n708), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n773), .A2(new_n845), .ZN(G396));
  NAND2_X1  g0646(.A1(new_n676), .A2(new_n712), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n374), .B1(new_n362), .B2(new_n712), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n372), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n684), .A2(new_n712), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(new_n640), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n643), .B(new_n642), .C1(new_n659), .C2(new_n660), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n753), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n712), .B(new_n853), .C1(new_n856), .C2(new_n674), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n771), .B1(new_n858), .B2(new_n752), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n752), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n775), .A2(new_n830), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n774), .B1(new_n223), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n782), .A2(G68), .ZN(new_n863));
  INV_X1    g0663(.A(G132), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n418), .B1(new_n789), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G58), .B2(new_n785), .ZN(new_n866));
  INV_X1    g0666(.A(new_n811), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n863), .B(new_n866), .C1(new_n202), .C2(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n796), .A2(G137), .B1(new_n807), .B2(G143), .ZN(new_n869));
  INV_X1    g0669(.A(G150), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n869), .B1(new_n870), .B2(new_n809), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G159), .B2(new_n804), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n868), .B1(new_n872), .B2(KEYINPUT34), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n872), .A2(KEYINPUT34), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n277), .B1(new_n824), .B2(new_n789), .C1(new_n571), .C2(new_n806), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n796), .A2(G303), .B1(new_n810), .B2(G283), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n225), .B2(new_n867), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n875), .B(new_n877), .C1(G116), .C2(new_n804), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n782), .A2(G87), .B1(G97), .B2(new_n786), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n873), .A2(new_n874), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n862), .B1(new_n776), .B2(new_n880), .C1(new_n853), .C2(new_n831), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n860), .A2(new_n881), .ZN(G384));
  INV_X1    g0682(.A(new_n540), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n491), .B(new_n213), .C1(new_n883), .C2(KEYINPUT35), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(KEYINPUT35), .B2(new_n883), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT36), .Z(new_n886));
  OR3_X1    g0686(.A1(new_n215), .A2(new_n223), .A3(new_n441), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n202), .A2(G68), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n261), .B(G13), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  INV_X1    g0691(.A(new_n697), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n450), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n451), .A2(new_n891), .A3(new_n459), .A4(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n447), .A2(new_n443), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n448), .B(new_n248), .C1(new_n895), .C2(new_n433), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n687), .A2(new_n697), .B1(new_n896), .B2(new_n432), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT37), .B1(new_n897), .B2(new_n462), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT98), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n697), .B1(new_n896), .B2(new_n432), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n464), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n894), .A2(KEYINPUT98), .A3(new_n898), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT38), .A4(new_n904), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT40), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT100), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n751), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n739), .A2(new_n740), .B1(new_n743), .B2(new_n551), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n747), .B(new_n712), .C1(new_n912), .C2(new_n738), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT31), .B1(new_n745), .B2(new_n699), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(KEYINPUT100), .A3(new_n749), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT97), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n348), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT97), .B(new_n328), .C1(new_n346), .C2(new_n347), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n328), .A2(new_n699), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n918), .A2(new_n352), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n346), .A2(new_n347), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n352), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n328), .A3(new_n699), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n851), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n911), .A2(new_n916), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n909), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n893), .B1(new_n691), .B2(new_n682), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n893), .A2(new_n891), .A3(new_n459), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n688), .A2(new_n450), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n893), .A3(new_n459), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n930), .A2(new_n451), .B1(new_n932), .B2(KEYINPUT37), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n906), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n908), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT40), .B1(new_n935), .B2(new_n926), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n465), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n911), .A2(new_n916), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n937), .A2(new_n940), .ZN(new_n942));
  INV_X1    g0742(.A(G330), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n908), .A2(new_n934), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT99), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n918), .A2(new_n919), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n712), .ZN(new_n951));
  AOI211_X1 g0751(.A(KEYINPUT99), .B(new_n699), .C1(new_n918), .C2(new_n919), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n945), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n857), .A2(new_n850), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n907), .A2(new_n908), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n921), .A2(new_n924), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n692), .A2(new_n697), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n955), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n938), .B1(new_n730), .B2(new_n760), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n693), .A2(new_n310), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n961), .B(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n944), .A2(new_n965), .B1(new_n261), .B2(new_n766), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n944), .A2(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n890), .B1(new_n966), .B2(new_n967), .ZN(G367));
  INV_X1    g0768(.A(KEYINPUT105), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n560), .B1(new_n557), .B2(new_n712), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n549), .A2(new_n552), .A3(new_n699), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n719), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  INV_X1    g0774(.A(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n718), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n975), .B2(new_n718), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT104), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n973), .A2(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n979), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n718), .A3(new_n978), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(KEYINPUT104), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n716), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n984), .A3(new_n716), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n717), .A2(new_n709), .ZN(new_n989));
  INV_X1    g0789(.A(new_n715), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n989), .B1(new_n990), .B2(new_n717), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n764), .B(new_n991), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n762), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n724), .B(KEYINPUT41), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n770), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n972), .A2(new_n989), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT42), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n638), .B1(new_n970), .B2(new_n667), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n712), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n647), .A2(new_n699), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n756), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n623), .A2(new_n1003), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT43), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT102), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n708), .A2(G330), .A3(new_n715), .A4(new_n972), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1002), .A2(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n999), .A2(new_n1001), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1006), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT101), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT101), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1002), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1010), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1009), .A2(new_n1008), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1019), .B(new_n1010), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n969), .B1(new_n996), .B2(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n770), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n987), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1027), .A2(new_n985), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n992), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n761), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1026), .B1(new_n1030), .B2(new_n994), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1025), .A2(new_n1031), .A3(KEYINPUT105), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1024), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n832), .A2(new_n775), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n837), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1034), .B1(new_n207), .B2(new_n354), .C1(new_n238), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT106), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n774), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n1037), .B2(new_n1036), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n811), .A2(G116), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT46), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n807), .A2(new_n518), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n418), .B1(new_n790), .B2(G317), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n796), .A2(G311), .B1(new_n810), .B2(G294), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n804), .A2(G283), .B1(new_n368), .B2(new_n785), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT107), .Z(new_n1047));
  AOI211_X1 g0847(.A(new_n1045), .B(new_n1047), .C1(G97), .C2(new_n782), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT108), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT109), .B(G137), .Z(new_n1050));
  OAI221_X1 g0850(.A(new_n367), .B1(new_n870), .B2(new_n806), .C1(new_n789), .C2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G50), .B2(new_n804), .ZN(new_n1052));
  INV_X1    g0852(.A(G159), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n867), .A2(new_n250), .B1(new_n1053), .B2(new_n809), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G143), .B2(new_n796), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n786), .A2(G68), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n782), .A2(G77), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1052), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1049), .A2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT47), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1039), .B1(new_n1060), .B2(new_n775), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n844), .B2(new_n1012), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1033), .A2(new_n1062), .ZN(G387));
  NAND2_X1  g0863(.A1(new_n1029), .A2(new_n762), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n992), .A2(new_n761), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n724), .A3(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n235), .A2(new_n466), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1067), .A2(new_n837), .B1(new_n722), .B2(new_n833), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n430), .A2(G50), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT50), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n466), .B1(new_n217), .B2(new_n223), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1071), .B(new_n722), .C1(new_n1070), .C2(new_n1069), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1068), .A2(new_n1072), .B1(G107), .B2(new_n207), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n774), .B1(new_n1073), .B2(new_n1034), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n799), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n807), .A2(G50), .B1(new_n1075), .B2(G68), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n810), .A2(new_n254), .B1(new_n811), .B2(G77), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n410), .B1(new_n790), .B2(G150), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n796), .A2(G159), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n786), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(new_n354), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(G97), .C2(new_n782), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n811), .A2(G294), .B1(new_n785), .B2(G283), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT110), .Z(new_n1085));
  AOI22_X1  g0885(.A1(G311), .A2(new_n810), .B1(new_n807), .B2(G317), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n823), .B2(new_n818), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n518), .B2(new_n804), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1088), .B2(KEYINPUT48), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT111), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(KEYINPUT48), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1092), .A2(KEYINPUT49), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n410), .B1(new_n819), .B2(new_n789), .C1(new_n781), .C2(new_n491), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1092), .B2(KEYINPUT49), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1083), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1074), .B1(new_n1096), .B2(new_n776), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n990), .B2(new_n832), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1029), .B2(new_n770), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1066), .A2(new_n1099), .ZN(G393));
  OR3_X1    g0900(.A1(new_n1027), .A2(new_n985), .A3(KEYINPUT112), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1027), .B1(new_n985), .B2(KEYINPUT112), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1026), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n975), .A2(new_n832), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1034), .B1(new_n495), .B2(new_n207), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n242), .A2(new_n837), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n771), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n810), .A2(new_n518), .B1(G116), .B2(new_n785), .ZN(new_n1108));
  INV_X1    g0908(.A(G283), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n867), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n799), .A2(new_n571), .B1(new_n789), .B2(new_n823), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1110), .A2(new_n367), .A3(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n796), .A2(G317), .B1(new_n807), .B2(G311), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1113), .A2(KEYINPUT52), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(KEYINPUT52), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1112), .A2(new_n783), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n804), .A2(new_n254), .B1(G50), .B2(new_n810), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(KEYINPUT113), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n410), .B1(new_n790), .B2(G143), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n217), .B2(new_n867), .C1(new_n781), .C2(new_n219), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(KEYINPUT113), .B2(new_n1118), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n818), .A2(new_n870), .B1(new_n1053), .B2(new_n806), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT51), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n786), .A2(G77), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1116), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1107), .B1(new_n1130), .B2(new_n775), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1103), .B1(new_n1104), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1101), .A2(new_n1064), .A3(new_n1102), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1133), .B(new_n724), .C1(new_n1064), .C2(new_n988), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(G390));
  OAI211_X1 g0935(.A(new_n712), .B(new_n849), .C1(new_n755), .C2(new_n758), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n850), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n958), .A2(KEYINPUT114), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT114), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n921), .A2(new_n1139), .A3(new_n924), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n946), .A2(new_n953), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n958), .A2(G330), .A3(new_n751), .A4(new_n853), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n945), .A2(new_n948), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n954), .B1(new_n956), .B2(new_n958), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1144), .B(new_n1145), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n911), .A2(new_n916), .A3(new_n925), .A4(G330), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n938), .A2(new_n939), .A3(new_n943), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n962), .A2(new_n1153), .A3(new_n963), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1141), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n911), .A2(new_n916), .A3(G330), .A4(new_n853), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1145), .A2(new_n1136), .A3(new_n850), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n921), .B(new_n924), .C1(new_n752), .C2(new_n851), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1150), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1157), .A2(new_n1158), .B1(new_n1160), .B2(new_n956), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1154), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1148), .B(new_n1152), .C1(new_n1162), .C2(KEYINPUT115), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1152), .A2(new_n1148), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1160), .A2(new_n956), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n962), .A2(new_n1153), .A3(new_n963), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT115), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1163), .A2(new_n1170), .A3(new_n724), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1152), .A2(new_n770), .A3(new_n1148), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n774), .B1(new_n430), .B2(new_n861), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n818), .A2(new_n1109), .B1(new_n867), .B2(new_n219), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n368), .B2(new_n810), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n277), .B1(new_n571), .B2(new_n789), .C1(new_n491), .C2(new_n806), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n804), .B2(G97), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1175), .A2(new_n863), .A3(new_n1127), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n811), .A2(G150), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT53), .Z(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n202), .B2(new_n781), .C1(new_n1053), .C2(new_n1081), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT54), .B(G143), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n804), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1050), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n796), .A2(G128), .B1(new_n810), .B2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n807), .A2(G132), .B1(new_n790), .B2(G125), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n367), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1178), .B1(new_n1181), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT116), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n775), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1173), .B1(new_n1191), .B2(new_n1193), .C1(new_n1146), .C2(new_n831), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1172), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1171), .A2(new_n1195), .ZN(G378));
  AOI21_X1  g0996(.A(KEYINPUT100), .B1(new_n915), .B2(new_n749), .ZN(new_n1197));
  AND4_X1   g0997(.A1(KEYINPUT100), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n946), .A3(new_n925), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(KEYINPUT40), .A2(new_n1200), .B1(new_n909), .B2(new_n927), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n681), .A2(new_n310), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n267), .A2(new_n697), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1205));
  INV_X1    g1005(.A(new_n1203), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n387), .A2(new_n390), .A3(KEYINPUT84), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT84), .B1(new_n387), .B2(new_n390), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n310), .B(new_n1206), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1204), .A2(new_n1205), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1205), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1206), .B1(new_n681), .B2(new_n310), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1209), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1201), .A2(new_n1215), .A3(new_n943), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n937), .B2(G330), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n961), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1215), .B1(new_n1201), .B2(new_n943), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n961), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n937), .A2(G330), .A3(new_n1217), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n770), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n861), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n771), .B1(G50), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n789), .A2(new_n1109), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n418), .A2(G41), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(G107), .C2(new_n807), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n796), .A2(G116), .B1(G77), .B2(new_n811), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1229), .A2(new_n1056), .A3(new_n1230), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n809), .A2(new_n495), .B1(new_n799), .B2(new_n354), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT117), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n782), .A2(G58), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1231), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  XOR2_X1   g1037(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1238));
  XNOR2_X1  g1038(.A(new_n1237), .B(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1228), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n786), .A2(G150), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n810), .A2(G132), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n807), .A2(G128), .B1(new_n1075), .B2(G137), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n796), .A2(G125), .B1(new_n811), .B2(new_n1183), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1247));
  AOI211_X1 g1047(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n1053), .C2(new_n781), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1239), .B(new_n1240), .C1(new_n1246), .C2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1226), .B1(new_n1250), .B2(new_n775), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1215), .B2(new_n831), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1224), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1219), .A2(KEYINPUT57), .A3(new_n1223), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1136), .A2(new_n850), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n946), .A2(new_n953), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n956), .A2(new_n958), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n953), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n945), .A2(new_n948), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1148), .B(new_n1167), .C1(new_n1262), .C2(new_n1150), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1263), .A2(new_n1168), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n724), .B1(new_n1255), .B2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1221), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1263), .A2(new_n1168), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT57), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1254), .B1(new_n1265), .B2(new_n1270), .ZN(G375));
  NOR2_X1   g1071(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1162), .A2(new_n1272), .A3(new_n994), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1273), .A2(KEYINPUT119), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1235), .A2(new_n418), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT120), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n790), .A2(G128), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1277), .B1(new_n870), .B2(new_n799), .C1(new_n806), .C2(new_n1050), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n810), .A2(new_n1183), .B1(new_n811), .B2(G159), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n864), .B2(new_n818), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n1278), .B(new_n1280), .C1(G50), .C2(new_n786), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n790), .A2(G303), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1282), .B(new_n277), .C1(new_n1109), .C2(new_n806), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n796), .A2(G294), .B1(new_n810), .B2(G116), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n495), .B2(new_n867), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1283), .B(new_n1285), .C1(new_n368), .C2(new_n804), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1082), .B1(G77), .B2(new_n782), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1276), .A2(new_n1281), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  OAI221_X1 g1088(.A(new_n771), .B1(G68), .B2(new_n1225), .C1(new_n1288), .C2(new_n776), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1155), .B2(new_n830), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1167), .B2(new_n770), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(KEYINPUT121), .Z(new_n1292));
  NAND2_X1  g1092(.A1(new_n1273), .A2(KEYINPUT119), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1274), .A2(new_n1292), .A3(new_n1293), .ZN(G381));
  NAND4_X1  g1094(.A1(new_n1066), .A2(new_n773), .A3(new_n845), .A4(new_n1099), .ZN(new_n1295));
  OR3_X1    g1095(.A1(G390), .A2(G384), .A3(new_n1295), .ZN(new_n1296));
  NOR4_X1   g1096(.A1(new_n1296), .A2(G387), .A3(G381), .A4(G378), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1297), .B(new_n1254), .C1(new_n1270), .C2(new_n1265), .ZN(G407));
  INV_X1    g1098(.A(G378), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n698), .A2(G213), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G407), .B(G213), .C1(G375), .C2(new_n1302), .ZN(G409));
  NAND3_X1  g1103(.A1(new_n1033), .A2(new_n1062), .A3(G390), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G390), .B1(new_n1033), .B2(new_n1062), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G393), .A2(G396), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1295), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1307), .B2(new_n1295), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1305), .A2(new_n1306), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(G390), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G387), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1310), .B1(new_n1314), .B2(new_n1304), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT122), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1219), .A2(new_n995), .A3(new_n1223), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1318), .B1(new_n1319), .B2(new_n1264), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1268), .A2(KEYINPUT122), .A3(new_n995), .A4(new_n1269), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT123), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1253), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1224), .A2(KEYINPUT123), .A3(new_n1252), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G378), .B1(new_n1322), .B2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G378), .B(new_n1254), .C1(new_n1265), .C2(new_n1270), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1317), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1154), .A2(new_n1161), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT60), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1331), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1162), .A2(new_n725), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1272), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1292), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(G384), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1292), .A2(new_n1338), .A3(G384), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1224), .A2(KEYINPUT123), .A3(new_n1252), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT123), .B1(new_n1224), .B2(new_n1252), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1299), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1349), .A2(KEYINPUT124), .A3(new_n1328), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1330), .A2(new_n1300), .A3(new_n1344), .A4(new_n1350), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1351), .A2(KEYINPUT62), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1300), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1301), .A2(G2897), .ZN(new_n1354));
  XOR2_X1   g1154(.A(new_n1354), .B(KEYINPUT126), .Z(new_n1355));
  INV_X1    g1155(.A(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1343), .A2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1341), .A2(new_n1342), .A3(new_n1355), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(KEYINPUT61), .B1(new_n1353), .B2(new_n1359), .ZN(new_n1360));
  OAI211_X1 g1160(.A(new_n1300), .B(new_n1344), .C1(new_n1327), .C2(new_n1329), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(KEYINPUT62), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1360), .A2(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1316), .B1(new_n1352), .B2(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT63), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1351), .A2(new_n1365), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1330), .A2(new_n1300), .A3(new_n1350), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(new_n1359), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1316), .A2(KEYINPUT61), .ZN(new_n1369));
  OR2_X1    g1169(.A1(new_n1361), .A2(new_n1365), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1366), .A2(new_n1368), .A3(new_n1369), .A4(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1364), .A2(new_n1371), .ZN(G405));
  AND2_X1   g1172(.A1(G375), .A2(new_n1299), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1373), .A2(new_n1329), .ZN(new_n1374));
  XNOR2_X1  g1174(.A(new_n1374), .B(new_n1343), .ZN(new_n1375));
  XNOR2_X1  g1175(.A(new_n1375), .B(new_n1316), .ZN(G402));
endmodule


