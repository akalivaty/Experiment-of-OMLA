//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(KEYINPUT64), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(KEYINPUT64), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n216), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n209), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G222), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  OR2_X1    g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n257), .A2(G223), .B1(new_n251), .B2(G77), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n264), .A2(G274), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(KEYINPUT66), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(G274), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(new_n267), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n267), .A2(KEYINPUT67), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n267), .A2(KEYINPUT67), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n274), .A2(new_n275), .A3(new_n260), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n261), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n278), .A2(G179), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT71), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n266), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n213), .B1(new_n206), .B2(new_n262), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n266), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G50), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G50), .B2(new_n285), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n212), .A2(G33), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n287), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n298), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n278), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n302), .A2(KEYINPUT70), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT70), .B1(new_n302), .B2(new_n304), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n280), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n300), .A2(KEYINPUT9), .A3(new_n301), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT74), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n278), .A2(G200), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n278), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n302), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT10), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n310), .A2(new_n318), .A3(new_n315), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n307), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n288), .A2(G77), .A3(new_n289), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(G77), .B2(new_n285), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  INV_X1    g0123(.A(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n262), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n212), .A2(new_n323), .B1(new_n295), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT64), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(KEYINPUT64), .A2(G20), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n262), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT15), .B(G87), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n326), .A2(KEYINPUT72), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(KEYINPUT72), .B2(new_n326), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n322), .B1(new_n287), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n276), .A2(G244), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n273), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n252), .A2(G232), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n257), .A2(G238), .B1(new_n251), .B2(G107), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n264), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(G200), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n336), .A2(KEYINPUT73), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n338), .A2(new_n341), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G190), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT73), .B1(new_n336), .B2(new_n342), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n344), .A2(G169), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n338), .A2(G179), .A3(new_n341), .ZN(new_n350));
  OR3_X1    g0150(.A1(new_n336), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n294), .B2(new_n323), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n354), .A2(KEYINPUT76), .A3(new_n287), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT76), .B1(new_n354), .B2(new_n287), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT11), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT11), .B1(new_n355), .B2(new_n356), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT12), .B1(new_n285), .B2(G68), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n216), .B1(new_n266), .B2(G20), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n359), .A2(new_n360), .B1(new_n288), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n357), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n276), .A2(G238), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G97), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n237), .A2(G1698), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G226), .B2(G1698), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n251), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n260), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n273), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n273), .A2(new_n364), .A3(KEYINPUT13), .A4(new_n369), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(KEYINPUT75), .ZN(new_n376));
  OAI21_X1  g0176(.A(G179), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(G169), .A3(new_n375), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT14), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n378), .A2(KEYINPUT14), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n363), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(G190), .B1(new_n374), .B2(new_n376), .ZN(new_n383));
  INV_X1    g0183(.A(new_n363), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n372), .A2(G200), .A3(new_n375), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n320), .A2(new_n352), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT78), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n324), .B1(new_n217), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G159), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n325), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n392), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n201), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n292), .A2(G159), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(KEYINPUT78), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n212), .A2(new_n251), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n255), .A2(new_n324), .A3(new_n256), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT7), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n405), .A3(G68), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n287), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n255), .A2(new_n256), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(new_n330), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n251), .A2(new_n402), .A3(new_n324), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G68), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n393), .A2(new_n395), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT16), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT79), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n413), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT79), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(new_n287), .A4(new_n407), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n295), .B1(new_n266), .B2(G20), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n288), .A2(new_n422), .B1(new_n286), .B2(new_n295), .ZN(new_n423));
  INV_X1    g0223(.A(G223), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n254), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G226), .B2(new_n254), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n426), .A2(new_n251), .B1(new_n262), .B2(new_n223), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n269), .A2(new_n272), .B1(new_n260), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n276), .A2(G232), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n312), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n428), .A2(new_n429), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(G200), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n421), .A2(new_n423), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT80), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n423), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n415), .B2(new_n420), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT80), .B1(new_n437), .B2(new_n432), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT17), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n421), .A2(new_n423), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n303), .B1(new_n428), .B2(new_n429), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(G179), .B2(new_n431), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT18), .B1(new_n437), .B2(new_n443), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n433), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n439), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n390), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n264), .A2(new_n266), .A3(G45), .A4(G274), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n224), .B1(new_n266), .B2(G45), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n264), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n409), .A2(G238), .A3(new_n254), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n262), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(G244), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n455), .B1(new_n461), .B2(new_n260), .ZN(new_n462));
  INV_X1    g0262(.A(G200), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT19), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n294), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n223), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n365), .A2(new_n465), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n330), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n409), .A2(new_n212), .A3(G68), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(new_n287), .B1(new_n286), .B2(new_n332), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n266), .A2(G33), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT83), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n288), .A2(G87), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n462), .A2(G190), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n462), .A2(G169), .ZN(new_n480));
  INV_X1    g0280(.A(G179), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n462), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n288), .A2(new_n476), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n474), .B1(new_n332), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n464), .A2(new_n479), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n285), .A2(G97), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n483), .B2(new_n466), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n492), .A2(new_n466), .A3(G107), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n212), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n292), .A2(G77), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT81), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n410), .A2(G107), .A3(new_n411), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n490), .B1(new_n501), .B2(new_n287), .ZN(new_n502));
  INV_X1    g0302(.A(new_n287), .ZN(new_n503));
  AOI211_X1 g0303(.A(KEYINPUT82), .B(new_n503), .C1(new_n499), .C2(new_n500), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n489), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n254), .C1(new_n249), .C2(new_n250), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n506), .A2(new_n507), .B1(G33), .B2(G283), .ZN(new_n509));
  NOR4_X1   g0309(.A1(new_n251), .A2(KEYINPUT84), .A3(new_n224), .A4(new_n254), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT84), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n257), .B2(G250), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT85), .B1(new_n514), .B2(G41), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT85), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n263), .A3(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n266), .B(G45), .C1(new_n263), .C2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n260), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n513), .A2(new_n260), .B1(G257), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n519), .B1(new_n515), .B2(new_n517), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n265), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n303), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(new_n481), .A3(new_n524), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n505), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n513), .A2(new_n260), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(G257), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n529), .A2(G190), .A3(new_n524), .A4(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n500), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n497), .B(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n494), .B1(new_n492), .B2(new_n491), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n212), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n287), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT82), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n501), .A2(new_n490), .A3(new_n287), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n488), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n525), .A2(G200), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n485), .B(new_n528), .C1(new_n533), .C2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n288), .A2(new_n476), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT25), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n285), .B2(G107), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n468), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n546), .A2(G107), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n328), .B(new_n329), .C1(new_n249), .C2(new_n250), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT87), .B1(new_n552), .B2(new_n223), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT87), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n409), .A2(new_n212), .A3(new_n554), .A4(G87), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(KEYINPUT22), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n409), .A2(new_n212), .A3(new_n557), .A4(G87), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT88), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n553), .A2(KEYINPUT88), .A3(KEYINPUT22), .A4(new_n555), .ZN(new_n562));
  NOR2_X1   g0362(.A1(KEYINPUT23), .A2(G107), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n330), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n324), .B1(new_n458), .B2(KEYINPUT23), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n468), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n561), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(KEYINPUT24), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n567), .B1(new_n556), .B2(new_n560), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(new_n562), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n287), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT89), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(KEYINPUT24), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(new_n571), .A3(new_n562), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(KEYINPUT89), .A3(new_n287), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n551), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n409), .A2(G257), .A3(G1698), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n409), .A2(G250), .A3(new_n254), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G294), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n260), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n521), .A2(G264), .B1(new_n265), .B2(new_n523), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(new_n312), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(G200), .B2(new_n588), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n545), .B1(new_n581), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n546), .A2(G116), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G283), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n466), .B2(G33), .ZN(new_n594));
  OAI221_X1 g0394(.A(new_n287), .B1(new_n324), .B2(G116), .C1(new_n330), .C2(new_n594), .ZN(new_n595));
  XOR2_X1   g0395(.A(new_n595), .B(KEYINPUT20), .Z(new_n596));
  NAND2_X1  g0396(.A1(new_n286), .A2(new_n457), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n409), .A2(G264), .A3(G1698), .ZN(new_n599));
  OAI211_X1 g0399(.A(G257), .B(new_n254), .C1(new_n249), .C2(new_n250), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n251), .A2(G303), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n260), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n521), .A2(G270), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n524), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n598), .B(new_n606), .C1(new_n312), .C2(new_n605), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(G169), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n598), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n611));
  AND4_X1   g0411(.A1(G179), .A2(new_n603), .A3(new_n524), .A4(new_n604), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n611), .A2(KEYINPUT21), .A3(G169), .A4(new_n605), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n607), .A2(new_n610), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT89), .B1(new_n579), .B2(new_n287), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n575), .B(new_n503), .C1(new_n577), .C2(new_n578), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n550), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n588), .A2(new_n303), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(G179), .B2(new_n588), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n615), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n451), .A2(new_n591), .A3(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n386), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n382), .B1(new_n624), .B2(new_n351), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n439), .A3(new_n449), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n447), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n317), .A2(new_n319), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n307), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n451), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n482), .A2(new_n484), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n528), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(KEYINPUT26), .A3(new_n485), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n479), .A2(new_n464), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n631), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n635), .B1(new_n637), .B2(new_n528), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n632), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT90), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n581), .A2(new_n643), .A3(new_n620), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT90), .B1(new_n618), .B2(new_n621), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n640), .B1(new_n646), .B2(new_n591), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n629), .B1(new_n630), .B2(new_n647), .ZN(G369));
  NAND3_X1  g0448(.A1(new_n212), .A2(new_n266), .A3(G13), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n598), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n641), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n615), .B2(new_n656), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT91), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n581), .A2(new_n590), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n618), .A2(new_n621), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n618), .A2(new_n654), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n618), .A2(new_n621), .A3(new_n654), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n643), .B1(new_n581), .B2(new_n620), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n618), .A2(KEYINPUT90), .A3(new_n621), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n655), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n642), .A2(new_n654), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n669), .A2(new_n672), .A3(new_n674), .ZN(G399));
  INV_X1    g0475(.A(new_n207), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n266), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n469), .A2(G116), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n678), .A2(new_n679), .B1(new_n219), .B2(new_n677), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT28), .Z(new_n681));
  AOI21_X1  g0481(.A(new_n641), .B1(new_n670), .B2(new_n671), .ZN(new_n682));
  INV_X1    g0482(.A(new_n591), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n639), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT94), .B1(new_n684), .B2(new_n655), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT94), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n684), .B2(new_n655), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n642), .B1(new_n581), .B2(new_n620), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n640), .B1(new_n591), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT29), .B1(new_n689), .B2(new_n654), .ZN(new_n690));
  OAI22_X1  g0490(.A1(KEYINPUT29), .A2(new_n685), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n655), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n462), .A2(new_n587), .A3(new_n586), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n612), .A3(new_n522), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n461), .A2(new_n260), .ZN(new_n699));
  INV_X1    g0499(.A(new_n455), .ZN(new_n700));
  AOI21_X1  g0500(.A(G179), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n701), .A2(new_n588), .A3(new_n605), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n696), .A2(new_n697), .B1(new_n702), .B2(new_n525), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT92), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n698), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n696), .A2(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n525), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n706), .A2(new_n707), .A3(new_n704), .ZN(new_n708));
  OAI211_X1 g0508(.A(KEYINPUT93), .B(new_n694), .C1(new_n705), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n698), .A2(new_n703), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n654), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n693), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n706), .A2(new_n707), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT92), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n703), .A2(new_n704), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n716), .A3(new_n698), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT93), .B1(new_n717), .B2(new_n694), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n591), .A2(new_n622), .A3(new_n655), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n692), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n691), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n681), .B1(new_n722), .B2(G1), .ZN(G364));
  AND2_X1   g0523(.A1(new_n212), .A2(G13), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G45), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n678), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n662), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n660), .A2(G330), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n658), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n409), .A2(new_n207), .ZN(new_n737));
  INV_X1    g0537(.A(G355), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n737), .A2(new_n738), .B1(G116), .B2(new_n207), .ZN(new_n739));
  INV_X1    g0539(.A(G45), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n244), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n676), .A2(new_n409), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n740), .B2(new_n219), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n739), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n213), .B1(G20), .B2(new_n303), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n734), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT96), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n728), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT97), .Z(new_n750));
  NOR4_X1   g0550(.A1(new_n324), .A2(new_n312), .A3(new_n463), .A4(G179), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT98), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT98), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n212), .A2(new_n481), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n312), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n756), .A2(G303), .B1(G322), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n212), .B1(new_n481), .B2(new_n758), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n764), .A2(G311), .B1(new_n766), .B2(G294), .ZN(new_n767));
  NOR3_X1   g0567(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n330), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G329), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n212), .A2(G179), .A3(G190), .A4(new_n463), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n251), .B(new_n771), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n757), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n776), .A2(new_n312), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G326), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n761), .A2(new_n767), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n765), .A2(new_n466), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n756), .B2(G87), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT32), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n769), .A2(new_n394), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n786), .B1(new_n763), .B2(new_n323), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n409), .B1(new_n773), .B2(new_n468), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G58), .B2(new_n760), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G50), .A2(new_n780), .B1(new_n777), .B2(G68), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n784), .A2(new_n788), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n782), .A2(new_n792), .A3(KEYINPUT99), .ZN(new_n793));
  AOI21_X1  g0593(.A(KEYINPUT99), .B1(new_n782), .B2(new_n792), .ZN(new_n794));
  INV_X1    g0594(.A(new_n746), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n750), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n729), .A2(new_n731), .B1(new_n736), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  OAI22_X1  g0599(.A1(new_n346), .A2(new_n347), .B1(new_n336), .B2(new_n655), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n351), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n351), .A2(new_n654), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n647), .B2(new_n654), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n352), .A2(new_n655), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n647), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n721), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n728), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n808), .B2(new_n807), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n755), .A2(new_n468), .B1(new_n811), .B2(new_n759), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n783), .B(new_n812), .C1(G116), .C2(new_n764), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n251), .B1(new_n814), .B2(new_n769), .C1(new_n773), .C2(new_n223), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G303), .B2(new_n780), .ZN(new_n816));
  INV_X1    g0616(.A(new_n777), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n813), .B(new_n816), .C1(new_n774), .C2(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G159), .A2(new_n764), .B1(new_n760), .B2(G143), .ZN(new_n819));
  INV_X1    g0619(.A(new_n780), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n819), .B1(new_n820), .B2(new_n821), .C1(new_n822), .C2(new_n817), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n773), .A2(new_n216), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G58), .B2(new_n766), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n202), .B2(new_n755), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n409), .B1(new_n769), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT101), .ZN(new_n831));
  OR3_X1    g0631(.A1(new_n825), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n823), .A2(new_n824), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n818), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n795), .B1(new_n834), .B2(KEYINPUT102), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(KEYINPUT102), .B2(new_n834), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n746), .A2(new_n732), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT100), .Z(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n727), .B1(new_n323), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n804), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n836), .B(new_n840), .C1(new_n733), .C2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n810), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G384));
  NAND2_X1  g0644(.A1(new_n363), .A2(new_n654), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT103), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n387), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n387), .A2(new_n846), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n804), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n711), .B(KEYINPUT31), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n720), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT105), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n433), .A2(new_n434), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n437), .A2(KEYINPUT80), .A3(new_n432), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n448), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n445), .A2(new_n446), .ZN(new_n858));
  INV_X1    g0658(.A(new_n449), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT16), .B1(new_n401), .B2(new_n406), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n423), .B1(new_n408), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n652), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n854), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n864), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n450), .A2(KEYINPUT105), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n440), .A2(KEYINPUT106), .A3(new_n444), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n440), .A2(new_n863), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT106), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n437), .B2(new_n443), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n869), .A2(new_n870), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n435), .A2(new_n438), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n862), .B1(new_n444), .B2(new_n863), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n855), .A2(new_n877), .A3(new_n856), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n875), .A2(new_n876), .B1(KEYINPUT37), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n868), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n882), .B(new_n879), .C1(new_n865), .C2(new_n867), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n853), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n888), .A2(new_n876), .A3(KEYINPUT107), .A4(new_n869), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT107), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n855), .A2(new_n856), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n890), .B1(new_n874), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n870), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n433), .B1(new_n437), .B2(new_n443), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n450), .A2(new_n893), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n879), .B1(new_n865), .B2(new_n867), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n849), .A2(KEYINPUT40), .A3(new_n851), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n887), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT110), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n451), .A2(new_n851), .ZN(new_n905));
  OAI21_X1  g0705(.A(G330), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n691), .A2(new_n451), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n629), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT108), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n450), .A2(KEYINPUT105), .A3(new_n866), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT105), .B1(new_n450), .B2(new_n866), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n880), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n882), .ZN(new_n914));
  OAI211_X1 g0714(.A(KEYINPUT38), .B(new_n880), .C1(new_n911), .C2(new_n912), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n896), .A2(new_n897), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n882), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n382), .A2(new_n654), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n916), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT104), .ZN(new_n924));
  INV_X1    g0724(.A(new_n806), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n802), .B1(new_n684), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n847), .A2(new_n848), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n924), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n803), .B1(new_n647), .B2(new_n806), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(KEYINPUT104), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n914), .A2(new_n915), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n858), .A2(new_n652), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n923), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n910), .B(new_n935), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n907), .A2(new_n936), .B1(new_n266), .B2(new_n724), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n907), .ZN(new_n938));
  INV_X1    g0738(.A(new_n537), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(KEYINPUT35), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(KEYINPUT35), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n940), .A2(G116), .A3(new_n214), .A4(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT36), .Z(new_n943));
  NAND3_X1  g0743(.A1(new_n219), .A2(G77), .A3(new_n392), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n202), .A2(G68), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n266), .B(G13), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n938), .A2(new_n943), .A3(new_n946), .ZN(G367));
  NAND2_X1  g0747(.A1(new_n234), .A2(new_n742), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n746), .B(new_n734), .C1(new_n676), .C2(new_n333), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n727), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n474), .A2(new_n477), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n654), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT111), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n632), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT112), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(KEYINPUT112), .C1(new_n637), .C2(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n765), .A2(new_n216), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n755), .A2(new_n215), .B1(new_n202), .B2(new_n763), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(G150), .C2(new_n760), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT115), .B(G137), .Z(new_n962));
  OAI221_X1 g0762(.A(new_n409), .B1(new_n769), .B2(new_n962), .C1(new_n773), .C2(new_n323), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G143), .B2(new_n780), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n961), .B(new_n964), .C1(new_n394), .C2(new_n817), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n755), .A2(new_n457), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n966), .A2(KEYINPUT46), .B1(G294), .B2(new_n777), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n814), .B2(new_n820), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n763), .A2(new_n774), .B1(new_n765), .B2(new_n468), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G303), .B2(new_n760), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n409), .B1(new_n772), .B2(G97), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n770), .A2(G317), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n970), .B(new_n973), .C1(new_n966), .C2(KEYINPUT46), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n965), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n950), .B1(new_n958), .B2(new_n735), .C1(new_n976), .C2(new_n795), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n726), .A2(G1), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n674), .A2(new_n672), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n528), .B1(new_n542), .B2(new_n655), .C1(new_n533), .C2(new_n544), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n633), .A2(new_n654), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT44), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n674), .A2(new_n672), .A3(new_n982), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n669), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(KEYINPUT114), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT114), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n986), .B(new_n989), .C1(new_n993), .C2(new_n669), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n674), .B1(new_n668), .B2(new_n673), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n661), .B(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n722), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT113), .B(KEYINPUT41), .Z(new_n999));
  XNOR2_X1  g0799(.A(new_n677), .B(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n978), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n664), .A2(new_n980), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n654), .B1(new_n1003), .B2(new_n528), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n674), .A2(new_n983), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1004), .B1(new_n1005), .B2(KEYINPUT42), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT42), .B2(new_n1005), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n1007), .A2(KEYINPUT43), .A3(new_n958), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n957), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n669), .A2(new_n983), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1013), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n977), .B1(new_n1002), .B2(new_n1016), .ZN(G387));
  INV_X1    g0817(.A(new_n722), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(new_n997), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n997), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n1020), .A3(new_n677), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n978), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n997), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n666), .A2(new_n667), .A3(new_n734), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n737), .A2(new_n679), .B1(G107), .B2(new_n207), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n240), .A2(G45), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n679), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1027), .C1(G68), .C2(G77), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n295), .A2(G50), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n743), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1025), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n728), .B1(new_n1032), .B2(new_n748), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n409), .B1(new_n822), .B2(new_n769), .C1(new_n773), .C2(new_n466), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G159), .B2(new_n780), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n756), .A2(G77), .B1(G50), .B2(new_n760), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n764), .A2(G68), .B1(new_n766), .B2(new_n333), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n295), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n777), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n409), .B1(new_n770), .B2(G326), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n755), .A2(new_n811), .B1(new_n774), .B2(new_n765), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G303), .A2(new_n764), .B1(new_n760), .B2(G317), .ZN(new_n1043));
  INV_X1    g0843(.A(G322), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n820), .B2(new_n1044), .C1(new_n814), .C2(new_n817), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1041), .B1(new_n457), .B2(new_n773), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1040), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1033), .B1(new_n1052), .B2(new_n746), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1023), .B1(new_n1024), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1021), .A2(new_n1054), .ZN(G393));
  NAND2_X1  g0855(.A1(new_n990), .A2(new_n991), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n986), .A2(new_n989), .A3(new_n669), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n978), .A3(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n747), .B1(new_n466), .B2(new_n207), .C1(new_n247), .C2(new_n743), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n728), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n770), .A2(G143), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n409), .B(new_n1061), .C1(new_n773), .C2(new_n223), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n756), .A2(G68), .B1(G77), .B2(new_n766), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n295), .B2(new_n763), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1062), .B(new_n1064), .C1(G50), .C2(new_n777), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n780), .A2(G150), .B1(new_n760), .B2(G159), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT116), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n780), .A2(G317), .B1(new_n760), .B2(G311), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n251), .B1(new_n1044), .B2(new_n769), .C1(new_n773), .C2(new_n468), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G303), .B2(new_n777), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n764), .A2(G294), .B1(new_n766), .B2(G116), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n774), .C2(new_n755), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1070), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1060), .B1(new_n1077), .B2(new_n746), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n982), .B2(new_n735), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n677), .B1(new_n1019), .B2(new_n995), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1018), .A2(new_n997), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1058), .B(new_n1079), .C1(new_n1080), .C2(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(new_n677), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n719), .A2(new_n720), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1086), .A2(G330), .A3(new_n841), .A4(new_n927), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n591), .A2(new_n688), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n654), .B1(new_n1088), .B2(new_n639), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n802), .B1(new_n1089), .B2(new_n801), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(new_n928), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n922), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(new_n919), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n916), .A2(new_n921), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n922), .B1(new_n930), .B2(new_n927), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1087), .B(new_n1093), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n692), .B1(new_n720), .B2(new_n850), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1097), .A2(new_n849), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n921), .B2(new_n916), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1091), .A2(new_n1092), .A3(new_n919), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n451), .A2(new_n1097), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n908), .A2(new_n629), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n927), .B1(new_n1097), .B2(new_n841), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT117), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n591), .A2(new_n622), .A3(new_n655), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n694), .B1(new_n705), .B2(new_n708), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT93), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n709), .A3(new_n712), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n841), .C1(new_n1109), .C2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1114), .A2(new_n928), .B1(new_n849), .B2(new_n1097), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1108), .B1(new_n1115), .B2(new_n926), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n927), .B1(new_n721), .B2(new_n841), .ZN(new_n1117));
  OAI211_X1 g0917(.A(KEYINPUT117), .B(new_n930), .C1(new_n1117), .C2(new_n1098), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1107), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1104), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1085), .B1(new_n1102), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1104), .A2(new_n1119), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n1096), .A3(new_n1101), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1096), .A2(new_n1101), .A3(new_n978), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n728), .B1(new_n1038), .B2(new_n838), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n409), .B(new_n826), .C1(G294), .C2(new_n770), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n468), .B2(new_n817), .C1(new_n774), .C2(new_n820), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G97), .A2(new_n764), .B1(new_n760), .B2(G116), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n323), .B2(new_n765), .C1(new_n223), .C2(new_n755), .ZN(new_n1130));
  OR3_X1    g0930(.A1(new_n755), .A2(KEYINPUT53), .A3(new_n822), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n780), .A2(G128), .ZN(new_n1132));
  OAI21_X1  g0932(.A(KEYINPUT53), .B1(new_n755), .B2(new_n822), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n759), .A2(new_n829), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n817), .A2(new_n962), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n770), .A2(G125), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n409), .B(new_n1137), .C1(new_n773), .C2(new_n202), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n763), .A2(new_n1139), .B1(new_n765), .B2(new_n394), .ZN(new_n1140));
  OR4_X1    g0940(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1128), .A2(new_n1130), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1126), .B1(new_n1142), .B2(new_n746), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1094), .B2(new_n733), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1125), .A2(KEYINPUT118), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT118), .B1(new_n1125), .B2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1124), .B1(new_n1146), .B2(new_n1147), .ZN(G378));
  OAI21_X1  g0948(.A(new_n728), .B1(G50), .B2(new_n838), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n302), .A2(new_n863), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT55), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n320), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n320), .A2(new_n1153), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1151), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1156), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n1150), .A3(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(new_n733), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n409), .A2(G41), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G50), .B(new_n1162), .C1(new_n262), .C2(new_n263), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1162), .B1(new_n774), .B2(new_n769), .C1(new_n773), .C2(new_n215), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G77), .B2(new_n756), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT119), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n959), .B1(new_n333), .B2(new_n764), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n468), .B2(new_n759), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n466), .A2(new_n817), .B1(new_n820), .B2(new_n457), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1163), .B1(new_n1170), .B2(KEYINPUT58), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n755), .A2(new_n1139), .B1(new_n821), .B2(new_n763), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G128), .B2(new_n760), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n780), .A2(G125), .B1(G150), .B2(new_n766), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT120), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1173), .B1(new_n829), .B2(new_n817), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n262), .B(new_n263), .C1(new_n773), .C2(new_n394), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G124), .B2(new_n770), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1171), .B1(KEYINPUT58), .B2(new_n1170), .C1(new_n1179), .C2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1149), .B(new_n1161), .C1(new_n746), .C2(new_n1184), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n923), .A2(new_n933), .A3(new_n934), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n885), .B1(new_n932), .B2(new_n853), .ZN(new_n1187));
  OAI21_X1  g0987(.A(G330), .B1(new_n900), .B2(new_n901), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n1160), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1160), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n901), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n692), .B1(new_n919), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1190), .B1(new_n887), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1186), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT123), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT123), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT122), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n935), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1160), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n887), .A2(new_n1192), .A3(new_n1190), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT123), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n935), .A2(new_n1198), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1195), .A2(new_n1200), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1185), .B1(new_n1206), .B2(new_n978), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1104), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1123), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1123), .A2(new_n1208), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1201), .A2(new_n935), .A3(new_n1202), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n935), .B1(new_n1202), .B2(new_n1201), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n677), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1207), .B1(new_n1210), .B2(new_n1215), .ZN(G375));
  OR3_X1    g1016(.A1(new_n1119), .A2(KEYINPUT124), .A3(new_n1022), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n838), .A2(G68), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n760), .A2(G283), .B1(new_n766), .B2(new_n333), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n468), .B2(new_n763), .C1(new_n755), .C2(new_n466), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n251), .B1(new_n773), .B2(new_n323), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G303), .B2(new_n770), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n457), .B2(new_n817), .C1(new_n811), .C2(new_n820), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n409), .B1(new_n773), .B2(new_n215), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G128), .B2(new_n770), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n829), .B2(new_n820), .C1(new_n817), .C2(new_n1139), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n764), .A2(G150), .B1(new_n766), .B2(G50), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n759), .B2(new_n962), .C1(new_n755), .C2(new_n394), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1220), .A2(new_n1223), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n727), .B(new_n1218), .C1(new_n1229), .C2(new_n746), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n927), .B2(new_n733), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT124), .B1(new_n1119), .B2(new_n1022), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1217), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1104), .A2(new_n1119), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1122), .A2(new_n1000), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(G381));
  INV_X1    g1037(.A(G390), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n843), .A3(new_n1239), .ZN(new_n1240));
  OR3_X1    g1040(.A1(new_n1240), .A2(G387), .A3(G381), .ZN(new_n1241));
  OR3_X1    g1041(.A1(new_n1241), .A2(G378), .A3(G375), .ZN(G407));
  NAND2_X1  g1042(.A1(new_n653), .A2(G213), .ZN(new_n1243));
  OR3_X1    g1043(.A1(G375), .A2(G378), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G407), .A2(G213), .A3(new_n1244), .ZN(G409));
  OAI211_X1 g1045(.A(G378), .B(new_n1207), .C1(new_n1210), .C2(new_n1215), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1213), .A2(new_n1196), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1001), .B(new_n1209), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1201), .A2(new_n935), .A3(new_n1202), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1194), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1185), .B1(new_n1251), .B2(new_n978), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1147), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1254), .A2(new_n1145), .B1(new_n1123), .B2(new_n1121), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1246), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1104), .A2(new_n1119), .A3(KEYINPUT60), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT125), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT60), .B1(new_n1104), .B2(new_n1119), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1260), .A2(new_n1122), .A3(new_n1085), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1233), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G384), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n843), .B(new_n1233), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1257), .A2(new_n1243), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1246), .A2(new_n1256), .B1(G213), .B2(new_n653), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(KEYINPUT126), .A3(new_n1266), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1269), .A2(KEYINPUT127), .A3(new_n1272), .A4(new_n1270), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(new_n1238), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G393), .B(new_n798), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G390), .B(new_n977), .C1(new_n1002), .C2(new_n1016), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1278), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n653), .A2(G213), .A3(G2897), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1266), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1284), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1282), .B(new_n1283), .C1(new_n1288), .C2(new_n1271), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1275), .A2(new_n1276), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1282), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT62), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1267), .A2(KEYINPUT62), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1257), .A2(new_n1243), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1297), .A3(new_n1283), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1293), .B1(new_n1294), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1292), .A2(new_n1299), .ZN(G405));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1255), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1246), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1266), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(new_n1293), .ZN(G402));
endmodule


