//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT29), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G211gat), .B(G218gat), .Z(new_n212));
  OAI21_X1  g011(.A(new_n204), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n203), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n217));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT2), .ZN(new_n219));
  INV_X1    g018(.A(G155gat), .ZN(new_n220));
  INV_X1    g019(.A(G162gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n217), .A2(new_n219), .B1(new_n222), .B2(new_n218), .ZN(new_n223));
  INV_X1    g022(.A(G141gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G148gat), .ZN(new_n225));
  INV_X1    g024(.A(G148gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G141gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n219), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n218), .ZN(new_n231));
  NOR2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n219), .B(new_n228), .C1(new_n233), .C2(new_n217), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT73), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n214), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n210), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n239), .A2(new_n210), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(new_n230), .B2(new_n234), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(KEYINPUT29), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n237), .A2(new_n245), .B1(G228gat), .B2(G233gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n204), .B1(new_n241), .B2(new_n242), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT82), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n203), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n212), .A2(KEYINPUT73), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n211), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT29), .B1(new_n251), .B2(new_n240), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(KEYINPUT82), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n236), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n245), .A2(G228gat), .A3(G233gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n246), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT83), .B(G22gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n202), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n258), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT3), .B1(new_n252), .B2(KEYINPUT82), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n247), .A2(new_n248), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n235), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n245), .A2(G228gat), .A3(G233gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g064(.A(KEYINPUT84), .B(new_n257), .C1(new_n265), .C2(new_n246), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n259), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G78gat), .B(G106gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT31), .B(G50gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(KEYINPUT81), .Z(new_n271));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT85), .B1(new_n265), .B2(new_n246), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n270), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n256), .B2(new_n258), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n267), .A2(new_n271), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n243), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT66), .ZN(new_n287));
  NOR2_X1   g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n283), .A2(KEYINPUT65), .A3(new_n285), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n287), .A2(new_n289), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  AND4_X1   g098(.A1(KEYINPUT25), .A2(new_n296), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  INV_X1    g101(.A(new_n290), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n303), .A2(new_n304), .A3(new_n288), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT67), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n310), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n284), .A2(KEYINPUT28), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n324), .A2(new_n299), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n295), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n317), .A2(new_n318), .ZN(new_n328));
  NOR2_X1   g127(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n325), .A2(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n309), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n313), .B1(new_n311), .B2(new_n312), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT67), .A3(new_n318), .ZN(new_n333));
  AOI21_X1  g132(.A(G190gat), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n309), .C1(new_n334), .C2(new_n321), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n308), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n323), .A2(new_n330), .B1(new_n301), .B2(new_n307), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n341), .B(new_n338), .C1(new_n342), .C2(KEYINPUT29), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n330), .B1(new_n334), .B2(new_n321), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n308), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT75), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  AND4_X1   g145(.A1(new_n282), .A2(new_n340), .A3(new_n343), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n308), .A2(new_n344), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT74), .B1(new_n348), .B2(new_n339), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n350));
  AOI211_X1 g149(.A(new_n350), .B(new_n338), .C1(new_n308), .C2(new_n344), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n353), .A2(new_n335), .B1(new_n307), .B2(new_n301), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n338), .B1(new_n354), .B2(KEYINPUT29), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n282), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n281), .B1(new_n347), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n339), .B1(new_n337), .B2(new_n204), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n350), .B1(new_n342), .B2(new_n338), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n339), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n243), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n340), .A2(new_n282), .A3(new_n346), .A4(new_n343), .ZN(new_n363));
  INV_X1    g162(.A(new_n281), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n357), .A2(KEYINPUT30), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n347), .A2(new_n356), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT30), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n368), .A3(new_n364), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT40), .ZN(new_n371));
  OR2_X1    g170(.A1(G127gat), .A2(G134gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G113gat), .B(G120gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(KEYINPUT1), .ZN(new_n374));
  OR2_X1    g173(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(G127gat), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT70), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  INV_X1    g179(.A(G113gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(G120gat), .ZN(new_n382));
  INV_X1    g181(.A(G120gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(G113gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n380), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT70), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n372), .A4(new_n377), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(G127gat), .B(G134gat), .Z(new_n389));
  NOR2_X1   g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n393));
  INV_X1    g192(.A(new_n244), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n235), .A3(new_n391), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n390), .B1(new_n379), .B2(new_n387), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n235), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n402), .B(KEYINPUT77), .Z(new_n403));
  XOR2_X1   g202(.A(KEYINPUT86), .B(KEYINPUT39), .Z(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT80), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n407), .B(G57gat), .Z(new_n408));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409));
  INV_X1    g208(.A(G85gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n408), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n392), .A2(new_n236), .ZN(new_n414));
  INV_X1    g213(.A(new_n403), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n396), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT39), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n403), .B2(new_n401), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n371), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n417), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n403), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n422), .A2(KEYINPUT40), .A3(new_n412), .A4(new_n405), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n415), .B(new_n395), .C1(new_n397), .C2(new_n400), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT78), .ZN(new_n425));
  AOI221_X4 g224(.A(new_n390), .B1(new_n230), .B2(new_n234), .C1(new_n379), .C2(new_n387), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n235), .B1(new_n388), .B2(new_n391), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n403), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT5), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT78), .ZN(new_n432));
  INV_X1    g231(.A(new_n412), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n419), .A2(new_n423), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n278), .B1(new_n370), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n362), .A2(new_n438), .A3(new_n363), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n281), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n362), .B2(new_n363), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT38), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT88), .B(KEYINPUT38), .C1(new_n440), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n282), .B1(new_n358), .B2(new_n361), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n340), .A2(new_n243), .A3(new_n346), .A4(new_n343), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT37), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n447), .A2(KEYINPUT87), .A3(KEYINPUT37), .A4(new_n448), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n364), .A2(KEYINPUT38), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n439), .A4(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT78), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n429), .B1(KEYINPUT78), .B2(new_n424), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n412), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n434), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n431), .A2(KEYINPUT6), .A3(new_n432), .A4(new_n433), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n454), .A2(new_n459), .A3(new_n460), .A4(new_n365), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n436), .B(new_n437), .C1(new_n446), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n459), .A2(new_n460), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n452), .A2(new_n439), .A3(new_n453), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n465), .A2(new_n451), .B1(new_n367), .B2(new_n364), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n464), .A2(new_n466), .A3(new_n444), .A4(new_n445), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n437), .B1(new_n467), .B2(new_n436), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n278), .B1(new_n464), .B2(new_n370), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  INV_X1    g270(.A(G227gat), .ZN(new_n472));
  INV_X1    g271(.A(G233gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT64), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n337), .A2(new_n392), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n354), .A2(new_n399), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT32), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G43gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(G71gat), .B(G99gat), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n337), .A2(new_n392), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n354), .A2(new_n399), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n475), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n489), .B2(KEYINPUT33), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT32), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n487), .A2(new_n488), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n476), .A2(KEYINPUT34), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n487), .B(new_n488), .C1(new_n472), .C2(new_n473), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n495), .A2(new_n496), .B1(new_n497), .B2(KEYINPUT34), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n486), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n486), .B2(new_n493), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n471), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n495), .A2(new_n496), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(KEYINPUT34), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n492), .ZN(new_n506));
  AOI221_X4 g305(.A(new_n491), .B1(KEYINPUT33), .B2(new_n485), .C1(new_n494), .C2(new_n476), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(KEYINPUT71), .A3(new_n499), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n471), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n502), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI211_X1 g313(.A(KEYINPUT72), .B(new_n471), .C1(new_n509), .C2(new_n511), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n470), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n464), .A2(new_n370), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n278), .B1(new_n509), .B2(new_n511), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n278), .A2(new_n500), .A3(new_n501), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OAI22_X1  g322(.A1(new_n469), .A2(new_n516), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(KEYINPUT90), .ZN(new_n526));
  INV_X1    g325(.A(G1gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(KEYINPUT90), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n526), .A2(new_n528), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(G1gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G8gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n529), .B2(KEYINPUT91), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n535), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  OR3_X1    g338(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n540), .A2(new_n541), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n538), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n536), .A2(new_n537), .ZN(new_n550));
  INV_X1    g349(.A(new_n548), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT94), .B1(new_n550), .B2(new_n551), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT92), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT13), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(KEYINPUT17), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n548), .A2(KEYINPUT17), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n556), .B1(KEYINPUT93), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n552), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n562), .A2(KEYINPUT93), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n561), .A2(new_n565), .A3(new_n552), .A4(new_n563), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n558), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  INV_X1    g369(.A(G197gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT11), .B(G169gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n558), .A2(new_n567), .A3(new_n568), .A4(new_n575), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(KEYINPUT95), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n566), .A2(new_n564), .B1(new_n554), .B2(new_n557), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n575), .B1(new_n581), .B2(new_n568), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT98), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT7), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT8), .ZN(new_n592));
  AND2_X1   g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  OAI221_X1 g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .C1(G85gat), .C2(G92gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n594), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G57gat), .B(G64gat), .Z(new_n599));
  INV_X1    g398(.A(KEYINPUT9), .ZN(new_n600));
  INV_X1    g399(.A(G71gat), .ZN(new_n601));
  INV_X1    g400(.A(G78gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G71gat), .B(G78gat), .Z(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n598), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n594), .B(new_n596), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n608), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n608), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n598), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n610), .B2(new_n612), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n589), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n614), .A2(new_n617), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT97), .ZN(new_n625));
  INV_X1    g424(.A(new_n619), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n618), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n622), .A2(new_n588), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n623), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n585), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n616), .A2(KEYINPUT21), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n609), .A2(KEYINPUT21), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n538), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n550), .B1(KEYINPUT21), .B2(new_n609), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n316), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G211gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n638), .B(new_n641), .Z(new_n642));
  XOR2_X1   g441(.A(G127gat), .B(G155gat), .Z(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n638), .B(new_n641), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AND3_X1   g449(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n598), .A2(KEYINPUT17), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n548), .ZN(new_n655));
  MUX2_X1   g454(.A(new_n653), .B(new_n652), .S(new_n655), .Z(new_n656));
  XOR2_X1   g455(.A(G134gat), .B(G162gat), .Z(new_n657));
  XNOR2_X1  g456(.A(G190gat), .B(G218gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n656), .B(new_n659), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n650), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n633), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n524), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n464), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT99), .B(G1gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1324gat));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n370), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT42), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT101), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n663), .A2(KEYINPUT42), .A3(new_n370), .A4(new_n671), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n673), .B(new_n674), .C1(new_n534), .C2(new_n669), .ZN(G1325gat));
  NOR2_X1   g474(.A1(new_n500), .A2(new_n501), .ZN(new_n676));
  AOI21_X1  g475(.A(G15gat), .B1(new_n663), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n514), .A2(new_n515), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n663), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n278), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  XNOR2_X1  g482(.A(new_n656), .B(new_n659), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n524), .A2(KEYINPUT44), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n580), .A2(new_n582), .ZN(new_n687));
  AOI211_X1 g486(.A(KEYINPUT95), .B(new_n575), .C1(new_n581), .C2(new_n568), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n579), .A2(new_n583), .A3(KEYINPUT103), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n690), .A2(new_n692), .A3(new_n631), .A4(new_n650), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n469), .B2(new_n516), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n436), .B1(new_n446), .B2(new_n461), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT89), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n462), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n509), .A2(new_n511), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT72), .B1(new_n699), .B2(new_n471), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n512), .A2(new_n513), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n701), .A3(new_n502), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n698), .A2(new_n702), .A3(KEYINPUT104), .A4(new_n470), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n695), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n520), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(KEYINPUT105), .A3(new_n522), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n523), .B2(new_n520), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n660), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n685), .B(new_n693), .C1(new_n711), .C2(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT106), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n709), .B1(new_n695), .B2(new_n703), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n660), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n685), .A4(new_n693), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n464), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n524), .A2(new_n684), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n633), .A2(new_n650), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n726), .A2(G29gat), .A3(new_n721), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n722), .A2(new_n729), .ZN(G1328gat));
  INV_X1    g529(.A(new_n370), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n720), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n726), .A2(G36gat), .A3(new_n731), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1329gat));
  OAI21_X1  g534(.A(G43gat), .B1(new_n712), .B2(new_n702), .ZN(new_n736));
  INV_X1    g535(.A(G43gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n725), .A2(new_n737), .A3(new_n676), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(KEYINPUT47), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n738), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n719), .A2(new_n678), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(G43gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g542(.A(G50gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n725), .A2(new_n744), .A3(new_n278), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n278), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n713), .B2(new_n718), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(new_n744), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  OAI21_X1  g550(.A(G50gat), .B1(new_n712), .B2(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n745), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT48), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n750), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n751), .B1(new_n750), .B2(new_n754), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(G1331gat));
  NAND2_X1  g556(.A1(new_n704), .A2(new_n710), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n690), .A2(new_n692), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n759), .A2(new_n632), .A3(new_n661), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n464), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g563(.A(new_n761), .B(KEYINPUT108), .Z(new_n765));
  XOR2_X1   g564(.A(new_n370), .B(KEYINPUT109), .Z(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n767), .B2(new_n768), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n765), .B2(new_n702), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n762), .A2(new_n601), .A3(new_n676), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1334gat));
  NOR2_X1   g575(.A1(new_n765), .A2(new_n748), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n602), .ZN(G1335gat));
  NOR3_X1   g577(.A1(new_n759), .A2(new_n632), .A3(new_n650), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n716), .A2(new_n685), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780), .B2(new_n721), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n759), .A2(new_n650), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n711), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT51), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n711), .A2(new_n785), .A3(new_n782), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n631), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n464), .A2(new_n410), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n781), .B1(new_n787), .B2(new_n788), .ZN(G1336gat));
  OR3_X1    g588(.A1(new_n787), .A2(G92gat), .A3(new_n766), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  OAI21_X1  g590(.A(G92gat), .B1(new_n780), .B2(new_n766), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G92gat), .B1(new_n780), .B2(new_n731), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(new_n791), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n780), .B2(new_n702), .ZN(new_n797));
  INV_X1    g596(.A(G99gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n676), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n787), .B2(new_n799), .ZN(G1338gat));
  NOR2_X1   g599(.A1(new_n748), .A2(G106gat), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n784), .A2(new_n631), .A3(new_n786), .A4(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n716), .A2(new_n278), .A3(new_n685), .A4(new_n779), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n808), .A3(G106gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n809), .A3(new_n802), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT53), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n810), .B2(KEYINPUT53), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(G1339gat));
  INV_X1    g613(.A(new_n521), .ZN(new_n815));
  INV_X1    g614(.A(new_n650), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n588), .B1(new_n620), .B2(KEYINPUT54), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n618), .B2(new_n619), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n818), .B(KEYINPUT55), .C1(new_n629), .C2(new_n819), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n629), .A2(new_n630), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n819), .B1(new_n625), .B2(new_n628), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n817), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n689), .A2(new_n691), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n554), .A2(new_n557), .ZN(new_n827));
  INV_X1    g626(.A(new_n556), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n561), .B2(new_n552), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n574), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n631), .A2(new_n578), .A3(new_n830), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT113), .Z(new_n832));
  AOI21_X1  g631(.A(new_n684), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n825), .A2(new_n578), .A3(new_n684), .A4(new_n830), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n816), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n661), .A2(new_n631), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n690), .B2(new_n692), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n815), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n766), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n721), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n584), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n721), .B1(new_n836), .B2(new_n838), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n519), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n766), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n759), .A2(new_n381), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(G1340gat));
  NOR3_X1   g647(.A1(new_n846), .A2(G120gat), .A3(new_n632), .ZN(new_n849));
  INV_X1    g648(.A(new_n842), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n383), .B1(new_n850), .B2(new_n631), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT114), .ZN(G1341gat));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT115), .B1(new_n846), .B2(new_n816), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n845), .A2(new_n856), .A3(new_n650), .A4(new_n766), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(G127gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n850), .B2(new_n650), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n854), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT116), .B(new_n861), .C1(new_n858), .C2(new_n859), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(G1342gat));
  XNOR2_X1  g664(.A(KEYINPUT69), .B(G134gat), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n845), .A2(new_n866), .A3(new_n731), .A4(new_n684), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n842), .B2(new_n660), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G1343gat));
  NOR2_X1   g670(.A1(new_n678), .A2(new_n748), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n844), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n840), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n584), .A2(G141gat), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT58), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n748), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n825), .A2(new_n583), .A3(new_n579), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n831), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n660), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n834), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT117), .B1(new_n882), .B2(new_n816), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n684), .B1(new_n879), .B2(new_n831), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT117), .B(new_n816), .C1(new_n884), .C2(new_n835), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n838), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n878), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n748), .B1(new_n836), .B2(new_n838), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n841), .A2(new_n702), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(KEYINPUT119), .A3(new_n585), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G141gat), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT119), .B1(new_n892), .B2(new_n585), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n876), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n889), .A2(KEYINPUT118), .A3(new_n891), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT118), .B1(new_n889), .B2(new_n891), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n759), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n899), .A2(G141gat), .B1(new_n874), .B2(new_n875), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(G1344gat));
  NAND3_X1  g701(.A1(new_n874), .A2(new_n226), .A3(new_n631), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G148gat), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n897), .A2(new_n898), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n631), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n837), .A2(new_n584), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT120), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n882), .A2(new_n816), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(KEYINPUT121), .A3(new_n910), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n748), .A2(KEYINPUT57), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n888), .A2(new_n877), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n916), .A2(new_n631), .A3(new_n891), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n904), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n903), .B1(new_n907), .B2(new_n919), .ZN(G1345gat));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n650), .B1(new_n897), .B2(new_n898), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G155gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n874), .A2(new_n220), .A3(new_n650), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n924), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT122), .B(new_n926), .C1(new_n922), .C2(G155gat), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n925), .A2(new_n927), .ZN(G1346gat));
  AND2_X1   g727(.A1(new_n906), .A2(new_n684), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n684), .A2(new_n221), .A3(new_n731), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n929), .A2(new_n221), .B1(new_n873), .B2(new_n930), .ZN(G1347gat));
  AOI21_X1  g730(.A(new_n464), .B1(new_n836), .B2(new_n838), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n766), .A2(new_n699), .A3(new_n278), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(G169gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n936), .A3(new_n759), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n731), .A2(new_n464), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n839), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(new_n585), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n940), .B2(new_n936), .ZN(G1348gat));
  AOI21_X1  g740(.A(G176gat), .B1(new_n935), .B2(new_n631), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n631), .A2(G176gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n939), .B2(new_n943), .ZN(G1349gat));
  OAI211_X1 g743(.A(new_n935), .B(new_n650), .C1(new_n319), .C2(new_n314), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n939), .A2(new_n946), .A3(new_n650), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G183gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n939), .B2(new_n650), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g750(.A(new_n310), .B1(new_n939), .B2(new_n684), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT61), .Z(new_n953));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n310), .A3(new_n684), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1351gat));
  NAND2_X1  g754(.A1(new_n916), .A2(new_n917), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n702), .A2(new_n938), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(G197gat), .B1(new_n959), .B2(new_n584), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n872), .A2(new_n840), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n963), .A2(new_n932), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n571), .A3(new_n759), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n960), .A2(new_n966), .ZN(G1352gat));
  OAI21_X1  g766(.A(G204gat), .B1(new_n959), .B2(new_n632), .ZN(new_n968));
  INV_X1    g767(.A(G204gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n965), .A2(new_n969), .A3(new_n631), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n973));
  OAI221_X1 g772(.A(new_n968), .B1(KEYINPUT62), .B2(new_n970), .C1(new_n972), .C2(new_n973), .ZN(G1353gat));
  NAND3_X1  g773(.A1(new_n965), .A2(new_n207), .A3(new_n650), .ZN(new_n975));
  INV_X1    g774(.A(new_n957), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n916), .A2(new_n650), .A3(new_n917), .A4(new_n976), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n207), .B1(new_n977), .B2(KEYINPUT127), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n978), .A2(KEYINPUT63), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  NOR3_X1   g781(.A1(new_n959), .A2(new_n208), .A3(new_n660), .ZN(new_n983));
  AOI21_X1  g782(.A(G218gat), .B1(new_n965), .B2(new_n684), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


