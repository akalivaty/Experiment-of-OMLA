//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(new_n203), .A2(G50), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(new_n207), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G77), .A2(G244), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G97), .A2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G87), .A2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G50), .A2(G226), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G68), .A2(G238), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n216), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n209), .B(new_n230), .C1(KEYINPUT1), .C2(new_n227), .ZN(G361));
  XOR2_X1   g0031(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G226), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT18), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT16), .ZN(new_n249));
  INV_X1    g0049(.A(G68), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n251), .A2(new_n252), .A3(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  OAI211_X1 g0055(.A(KEYINPUT7), .B(new_n207), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(KEYINPUT7), .B1(new_n260), .B2(new_n207), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n250), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(G58), .A2(G68), .ZN(new_n264));
  OAI21_X1  g0064(.A(G20), .B1(new_n264), .B2(new_n202), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G159), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT74), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n265), .A2(KEYINPUT74), .A3(new_n267), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n249), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n270), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  OAI21_X1  g0074(.A(G33), .B1(new_n251), .B2(new_n252), .ZN(new_n275));
  AOI21_X1  g0075(.A(G20), .B1(new_n275), .B2(new_n257), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT7), .ZN(new_n277));
  OAI21_X1  g0077(.A(G68), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n258), .A2(G33), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(G33), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n281), .A2(KEYINPUT7), .A3(G20), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n274), .B(KEYINPUT16), .C1(new_n278), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n208), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n272), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT8), .B(G58), .Z(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n285), .B1(new_n210), .B2(G20), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(G1), .B(G13), .C1(new_n254), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n210), .C1(G41), .C2(G45), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n295), .A2(G232), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  MUX2_X1   g0106(.A(G223), .B(G226), .S(G1698), .Z(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n281), .B2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n304), .B(KEYINPUT76), .C1(new_n308), .C2(new_n297), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(new_n275), .A3(new_n257), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n297), .B1(new_n312), .B2(new_n305), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n300), .A2(new_n303), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n309), .A2(new_n310), .A3(new_n315), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n314), .A2(KEYINPUT75), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  INV_X1    g0118(.A(new_n313), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(KEYINPUT75), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n248), .B1(new_n293), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n316), .A2(new_n321), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n286), .A2(new_n292), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT18), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n309), .A2(new_n327), .A3(new_n315), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n317), .A2(new_n329), .A3(new_n319), .A4(new_n320), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT17), .B1(new_n332), .B2(new_n325), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT17), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n331), .A2(new_n334), .A3(new_n286), .A4(new_n292), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n323), .A2(new_n326), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n279), .A2(new_n255), .ZN(new_n337));
  INV_X1    g0137(.A(G1698), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G222), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G77), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(G1698), .ZN(new_n341));
  INV_X1    g0141(.A(G223), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n339), .B1(new_n340), .B2(new_n337), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n295), .A2(new_n299), .A3(new_n297), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n302), .B1(new_n346), .B2(G226), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G200), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(G190), .A3(new_n347), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n266), .A2(G150), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n207), .A2(G33), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n288), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n201), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n207), .B1(new_n354), .B2(new_n202), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n285), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n289), .A2(G50), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n291), .B2(G50), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT9), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(KEYINPUT9), .A3(new_n358), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n349), .A2(new_n350), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT10), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n361), .A2(new_n362), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n350), .A4(new_n349), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n348), .A2(new_n310), .B1(new_n356), .B2(new_n358), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(G179), .B2(new_n348), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n337), .A2(G232), .A3(new_n338), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  INV_X1    g0172(.A(G238), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n371), .B1(new_n372), .B2(new_n337), .C1(new_n341), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n344), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n302), .B1(new_n346), .B2(G244), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G200), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n291), .A2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT68), .ZN(new_n380));
  INV_X1    g0180(.A(new_n289), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n340), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n287), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n352), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n285), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n380), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n378), .B(new_n388), .C1(new_n329), .C2(new_n377), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n377), .A2(new_n310), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n375), .A2(new_n318), .A3(new_n376), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n368), .A2(new_n370), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT69), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n368), .A2(new_n393), .A3(KEYINPUT69), .A4(new_n370), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT12), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n381), .B(new_n250), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n291), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n402), .B1(new_n250), .B2(new_n403), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n352), .A2(new_n340), .B1(new_n207), .B2(G68), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT71), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(new_n406), .B1(G50), .B2(new_n266), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n406), .B2(new_n405), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n285), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT11), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT11), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n411), .A3(new_n285), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n404), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n302), .B1(new_n346), .B2(G238), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n257), .A2(new_n259), .A3(G232), .A4(G1698), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n257), .A2(new_n259), .A3(G226), .A4(new_n338), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT70), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT70), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(G33), .A3(G97), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n416), .A2(new_n417), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n344), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n414), .A2(new_n415), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n415), .B1(new_n414), .B2(new_n423), .ZN(new_n426));
  OAI21_X1  g0226(.A(G200), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n414), .A2(new_n423), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT13), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(G190), .A3(new_n424), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n413), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n425), .B2(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n310), .B1(new_n429), .B2(new_n424), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n429), .A2(G179), .A3(new_n424), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n413), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n431), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND4_X1   g0240(.A1(new_n336), .A2(new_n396), .A3(new_n397), .A4(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n210), .B(G45), .C1(new_n296), .C2(KEYINPUT5), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n296), .A2(KEYINPUT5), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G274), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n297), .B(G257), .C1(new_n442), .C2(new_n443), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT4), .A2(G244), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n257), .A2(new_n259), .A3(new_n447), .A4(new_n338), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n257), .A2(new_n259), .A3(G250), .A4(G1698), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n450));
  AND3_X1   g0250(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT4), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n275), .A2(G244), .A3(new_n338), .A4(new_n257), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n445), .B(new_n446), .C1(new_n455), .C2(new_n297), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n454), .A2(new_n453), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n344), .B1(new_n458), .B2(new_n452), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(G190), .A3(new_n445), .A4(new_n446), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n372), .A2(KEYINPUT77), .A3(KEYINPUT6), .A4(G97), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT77), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT6), .A2(G97), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(G107), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n372), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G97), .A2(G107), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n461), .B(new_n464), .C1(new_n468), .C2(KEYINPUT6), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G20), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n266), .A2(G77), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n372), .B1(new_n256), .B2(new_n262), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n285), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n381), .A2(new_n465), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n475), .B(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n289), .B1(G1), .B2(new_n254), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n285), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(G97), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n457), .A2(new_n460), .A3(new_n474), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n474), .A2(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n456), .A2(new_n310), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n459), .A2(new_n318), .A3(new_n445), .A4(new_n446), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n275), .A2(G244), .A3(G1698), .A4(new_n257), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G116), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n373), .A2(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n275), .A2(new_n257), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n344), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n210), .A2(G45), .A3(G274), .ZN(new_n493));
  INV_X1    g0293(.A(G45), .ZN(new_n494));
  OAI21_X1  g0294(.A(G250), .B1(new_n494), .B2(G1), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n344), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n493), .B(KEYINPUT80), .C1(new_n344), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n492), .A2(G190), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n491), .A2(new_n344), .B1(new_n498), .B2(new_n499), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(KEYINPUT83), .A3(G190), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n492), .A2(new_n500), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G200), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n384), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(new_n289), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n479), .ZN(new_n512));
  INV_X1    g0312(.A(G87), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n352), .A2(new_n465), .ZN(new_n516));
  XNOR2_X1  g0316(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n275), .A2(new_n207), .A3(G68), .A4(new_n257), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n467), .A2(new_n513), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n419), .A2(new_n421), .ZN(new_n522));
  AOI21_X1  g0322(.A(G20), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n523), .B2(KEYINPUT82), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT82), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n525), .B(G20), .C1(new_n522), .C2(new_n517), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n520), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n285), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n511), .B(new_n515), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n512), .A2(new_n384), .ZN(new_n531));
  AOI211_X1 g0331(.A(new_n510), .B(new_n531), .C1(new_n527), .C2(new_n285), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n504), .A2(new_n318), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G169), .B2(new_n504), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n508), .A2(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n486), .A2(new_n535), .ZN(new_n536));
  MUX2_X1   g0336(.A(G250), .B(G257), .S(G1698), .Z(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n275), .A3(new_n257), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G294), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n297), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n297), .B(G264), .C1(new_n442), .C2(new_n443), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n445), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT87), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n540), .B2(new_n542), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n310), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n540), .A2(new_n542), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n318), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n513), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n281), .A2(new_n207), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n207), .A2(G87), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n550), .B1(new_n260), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n488), .A2(G20), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT23), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n207), .B2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n372), .A2(KEYINPUT23), .A3(G20), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n552), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n529), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n552), .A2(KEYINPUT24), .A3(new_n554), .A4(new_n559), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT25), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n289), .A2(new_n565), .A3(G107), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n289), .B2(G107), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n479), .A2(G107), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n547), .A2(new_n549), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n562), .B2(new_n563), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n327), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT88), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n540), .A2(new_n542), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(G200), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n546), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n578), .A2(G190), .A3(new_n544), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n572), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n289), .A2(G116), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n479), .B2(G116), .ZN(new_n583));
  AOI21_X1  g0383(.A(G20), .B1(new_n254), .B2(G97), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n451), .B2(new_n450), .ZN(new_n585));
  INV_X1    g0385(.A(G116), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n284), .A2(new_n208), .B1(G20), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(KEYINPUT20), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT20), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(KEYINPUT84), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n591), .B(KEYINPUT20), .C1(new_n585), .C2(new_n587), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n583), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  MUX2_X1   g0393(.A(G257), .B(G264), .S(G1698), .Z(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n275), .A3(new_n257), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n260), .A2(G303), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n344), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n297), .B(G270), .C1(new_n442), .C2(new_n443), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n445), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n329), .ZN(new_n603));
  AOI211_X1 g0403(.A(new_n593), .B(new_n603), .C1(G200), .C2(new_n602), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n297), .B1(new_n595), .B2(new_n596), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n605), .A2(new_n600), .A3(new_n318), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n593), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT85), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n593), .A2(KEYINPUT85), .A3(new_n606), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n310), .B1(new_n598), .B2(new_n601), .ZN(new_n611));
  NOR2_X1   g0411(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(new_n593), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n611), .B2(new_n593), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n609), .B(new_n610), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n604), .A2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n441), .A2(new_n536), .A3(new_n581), .A4(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n370), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n323), .A2(new_n326), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n333), .A2(new_n335), .ZN(new_n620));
  INV_X1    g0420(.A(new_n431), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n392), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n438), .B2(new_n439), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n619), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n618), .B1(new_n625), .B2(new_n368), .ZN(new_n626));
  INV_X1    g0426(.A(new_n441), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n535), .B2(new_n485), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n510), .B(new_n514), .C1(new_n527), .C2(new_n285), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n505), .A3(new_n507), .A4(new_n503), .ZN(new_n632));
  AOI21_X1  g0432(.A(G169), .B1(new_n492), .B2(new_n500), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n318), .B2(new_n504), .ZN(new_n634));
  INV_X1    g0434(.A(new_n531), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n511), .B(new_n635), .C1(new_n528), .C2(new_n529), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n630), .A2(new_n632), .A3(KEYINPUT26), .A4(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n629), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(G169), .B1(new_n578), .B2(new_n544), .ZN(new_n640));
  INV_X1    g0440(.A(new_n549), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n572), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n580), .B1(new_n615), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n632), .A2(new_n637), .A3(new_n481), .A4(new_n485), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n626), .B1(new_n627), .B2(new_n646), .ZN(G369));
  AND2_X1   g0447(.A1(new_n207), .A2(G13), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n210), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n593), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n616), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n615), .A2(new_n593), .A3(new_n654), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT89), .B1(new_n658), .B2(G330), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(KEYINPUT89), .A3(G330), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n654), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n581), .B1(new_n572), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n571), .B2(new_n663), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n615), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n581), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n642), .A2(new_n663), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n213), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n521), .A2(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n206), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n663), .B1(new_n639), .B2(new_n645), .ZN(new_n680));
  AND2_X1   g0480(.A1(KEYINPUT90), .A2(KEYINPUT29), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(KEYINPUT90), .A2(KEYINPUT29), .ZN(new_n684));
  OAI221_X1 g0484(.A(new_n663), .B1(new_n681), .B2(new_n684), .C1(new_n639), .C2(new_n645), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n459), .A2(new_n446), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n506), .A2(new_n548), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(new_n606), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n687), .A2(new_n688), .A3(KEYINPUT30), .A4(new_n606), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n575), .A2(G179), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n456), .A2(new_n693), .A3(new_n506), .A4(new_n602), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n695), .A2(new_n696), .A3(new_n654), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n536), .A2(new_n581), .A3(new_n616), .A4(new_n663), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n696), .B1(new_n695), .B2(new_n654), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n686), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n679), .B1(new_n703), .B2(G1), .ZN(G364));
  INV_X1    g0504(.A(new_n661), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n659), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT91), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n662), .A2(KEYINPUT91), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n210), .B1(new_n648), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n674), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n710), .B(new_n714), .C1(G330), .C2(new_n658), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n208), .B1(G20), .B2(new_n310), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n207), .A2(G190), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n719), .A2(new_n318), .A3(G200), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G311), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n327), .A2(G179), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n718), .ZN(new_n724));
  INV_X1    g0524(.A(G283), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n721), .A2(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n207), .A2(new_n329), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n723), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n337), .B(new_n726), .C1(G303), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n318), .A2(new_n327), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n718), .ZN(new_n732));
  XOR2_X1   g0532(.A(KEYINPUT33), .B(G317), .Z(new_n733));
  NAND2_X1  g0533(.A1(new_n727), .A2(new_n731), .ZN(new_n734));
  INV_X1    g0534(.A(G326), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n727), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n737), .A2(new_n318), .A3(G200), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G322), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n718), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n736), .B(new_n741), .C1(G329), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G294), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n207), .B1(new_n742), .B2(G190), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n730), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G50), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n337), .B1(new_n734), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G58), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n739), .A2(new_n751), .B1(new_n728), .B2(new_n513), .ZN(new_n752));
  INV_X1    g0552(.A(new_n747), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n750), .B(new_n752), .C1(G97), .C2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT93), .B(G159), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n743), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT32), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n732), .A2(new_n250), .B1(new_n724), .B2(new_n372), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(G77), .B2(new_n720), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n754), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n717), .B1(new_n748), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n716), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n281), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n213), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT92), .Z(new_n769));
  NAND2_X1  g0569(.A1(new_n243), .A2(G45), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(G45), .C2(new_n206), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n673), .A2(new_n260), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n772), .A2(G355), .B1(new_n586), .B2(new_n673), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n766), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n761), .A2(new_n774), .A3(new_n714), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n764), .B(KEYINPUT94), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n775), .B1(new_n658), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n715), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  OAI21_X1  g0579(.A(KEYINPUT99), .B1(new_n388), .B2(new_n663), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT99), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n387), .A2(new_n781), .A3(new_n654), .ZN(new_n782));
  AND3_X1   g0582(.A1(new_n389), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT98), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n392), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n390), .A2(KEYINPUT98), .A3(new_n387), .A4(new_n391), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n663), .B(new_n789), .C1(new_n639), .C2(new_n645), .ZN(new_n790));
  INV_X1    g0590(.A(new_n680), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n788), .B1(new_n392), .B2(new_n663), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n713), .B1(new_n793), .B2(new_n701), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n701), .B2(new_n793), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n717), .A2(new_n763), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n713), .B1(G77), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n724), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G68), .ZN(new_n799));
  INV_X1    g0599(.A(G132), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n749), .B2(new_n728), .C1(new_n800), .C2(new_n743), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n767), .B(new_n801), .C1(G58), .C2(new_n753), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT96), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(KEYINPUT96), .ZN(new_n804));
  INV_X1    g0604(.A(new_n732), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n738), .A2(G143), .B1(G150), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n807), .B2(new_n734), .C1(new_n755), .C2(new_n721), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT34), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n803), .A2(new_n804), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G303), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n734), .A2(new_n811), .B1(new_n732), .B2(new_n725), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G97), .B2(new_n753), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n738), .A2(G294), .B1(G311), .B2(new_n744), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n724), .A2(new_n513), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G116), .B2(new_n720), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n260), .B1(new_n728), .B2(new_n372), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT95), .Z(new_n819));
  OAI21_X1  g0619(.A(new_n810), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT97), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n717), .B1(new_n820), .B2(KEYINPUT97), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n797), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n763), .B2(new_n792), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n795), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  NOR3_X1   g0626(.A1(new_n208), .A2(new_n207), .A3(new_n586), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n469), .B2(KEYINPUT35), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT100), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n469), .A2(KEYINPUT35), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT36), .Z(new_n834));
  OR3_X1    g0634(.A1(new_n206), .A2(new_n340), .A3(new_n264), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n354), .A2(G68), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n210), .B(G13), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n437), .B1(new_n434), .B2(new_n435), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n439), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n654), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n652), .B(KEYINPUT103), .Z(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n325), .B1(new_n324), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n293), .A2(new_n331), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT104), .A4(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n322), .A2(new_n844), .B1(new_n286), .B2(new_n292), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n850), .B2(KEYINPUT104), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n325), .A2(new_n845), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n848), .B(new_n852), .C1(new_n336), .C2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n274), .B1(new_n278), .B2(new_n282), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n859), .A2(new_n249), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n283), .A2(new_n285), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n292), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n652), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n324), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n858), .B1(new_n293), .B2(new_n331), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n849), .A2(new_n858), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n863), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n866), .B(KEYINPUT38), .C1(new_n336), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n856), .A2(new_n857), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n619), .B2(new_n620), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n864), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n332), .A2(new_n325), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n858), .B1(new_n872), .B2(new_n850), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n855), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n868), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n869), .A2(KEYINPUT105), .B1(KEYINPUT39), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT105), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n856), .A2(new_n878), .A3(new_n857), .A4(new_n868), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n843), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n323), .A2(new_n326), .A3(new_n844), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n841), .A2(new_n663), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n439), .A2(new_n654), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n841), .A2(new_n621), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT101), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n440), .A2(KEYINPUT101), .A3(new_n883), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n785), .A2(new_n663), .A3(new_n786), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n790), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n876), .B1(new_n890), .B2(KEYINPUT102), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT102), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n892), .B(new_n888), .C1(new_n790), .C2(new_n889), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n881), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n880), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n441), .A2(new_n685), .A3(new_n683), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n626), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n895), .B(new_n897), .Z(new_n898));
  NAND2_X1  g0698(.A1(new_n441), .A2(new_n700), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT106), .Z(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  INV_X1    g0701(.A(new_n882), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n884), .A2(new_n885), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT101), .B1(new_n440), .B2(new_n883), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n700), .A3(new_n792), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n875), .A2(new_n868), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n901), .B1(new_n856), .B2(new_n868), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n700), .A2(new_n792), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n900), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n900), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(G330), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n898), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n210), .B2(new_n648), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n898), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n838), .B1(new_n917), .B2(new_n918), .ZN(G367));
  NOR2_X1   g0719(.A1(new_n631), .A2(new_n663), .ZN(new_n920));
  MUX2_X1   g0720(.A(new_n535), .B(new_n637), .S(new_n920), .Z(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n922), .A2(new_n776), .ZN(new_n923));
  INV_X1    g0723(.A(new_n769), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n765), .B1(new_n213), .B2(new_n384), .C1(new_n924), .C2(new_n239), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n713), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n724), .A2(new_n340), .ZN(new_n927));
  INV_X1    g0727(.A(G150), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n739), .A2(new_n928), .B1(new_n721), .B2(new_n354), .ZN(new_n929));
  INV_X1    g0729(.A(new_n734), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n927), .B(new_n929), .C1(G143), .C2(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n732), .A2(new_n755), .B1(new_n743), .B2(new_n807), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n260), .B(new_n932), .C1(G58), .C2(new_n729), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n931), .B(new_n933), .C1(new_n250), .C2(new_n747), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n767), .B1(new_n465), .B2(new_n724), .C1(new_n722), .C2(new_n734), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n728), .A2(new_n586), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT46), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n738), .A2(G303), .B1(G317), .B2(new_n744), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n938), .B(new_n939), .C1(new_n746), .C2(new_n732), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n720), .A2(G283), .B1(G107), .B2(new_n753), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT110), .Z(new_n942));
  OAI21_X1  g0742(.A(new_n934), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT47), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n717), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n926), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n923), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n486), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n482), .A2(new_n654), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT107), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT107), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n630), .A2(new_n654), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT108), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(new_n666), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n959), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n581), .A3(new_n667), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT42), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n485), .B1(new_n960), .B2(new_n571), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n663), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n965), .A2(new_n967), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n921), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n965), .A2(new_n967), .A3(new_n969), .A4(new_n921), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n961), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n961), .A3(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n665), .A2(new_n667), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n708), .A2(new_n709), .B1(new_n668), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n668), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n706), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n703), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT45), .B1(new_n962), .B2(new_n671), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n962), .A2(KEYINPUT45), .A3(new_n671), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n958), .A2(new_n670), .A3(new_n959), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n958), .A2(KEYINPUT44), .A3(new_n670), .A4(new_n959), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n985), .A2(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n666), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n983), .B1(new_n992), .B2(KEYINPUT109), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT109), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n666), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n989), .A2(new_n990), .ZN(new_n996));
  INV_X1    g0796(.A(new_n986), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n984), .ZN(new_n998));
  INV_X1    g0798(.A(new_n666), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n994), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n703), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n674), .B(KEYINPUT41), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n712), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n948), .B1(new_n976), .B2(new_n1004), .ZN(G387));
  NOR2_X1   g0805(.A1(new_n983), .A2(new_n675), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n703), .B2(new_n981), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n738), .A2(G317), .B1(G311), .B2(new_n805), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n811), .B2(new_n721), .C1(new_n740), .C2(new_n734), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT48), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n725), .B2(new_n747), .C1(new_n746), .C2(new_n728), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT49), .Z(new_n1012));
  OAI22_X1  g0812(.A1(new_n724), .A2(new_n586), .B1(new_n743), .B2(new_n735), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1012), .A2(new_n281), .A3(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G77), .A2(new_n729), .B1(new_n805), .B2(new_n287), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n465), .B2(new_n724), .C1(new_n749), .C2(new_n739), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n930), .A2(G159), .B1(new_n744), .B2(G150), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n250), .B2(new_n721), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n747), .A2(new_n384), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n1016), .A2(new_n1018), .A3(new_n767), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n716), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n665), .A2(new_n776), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n287), .A2(new_n749), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT111), .Z(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n676), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1027), .C1(G68), .C2(G77), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n236), .A2(G45), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n1030), .A3(new_n769), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n772), .A2(new_n1027), .B1(new_n372), .B2(new_n673), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n766), .B1(new_n1033), .B2(KEYINPUT112), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(KEYINPUT112), .B2(new_n1033), .ZN(new_n1035));
  AND4_X1   g0835(.A1(new_n713), .A2(new_n1021), .A3(new_n1022), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n981), .B2(new_n712), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1007), .A2(new_n1037), .ZN(G393));
  NAND3_X1  g0838(.A1(new_n995), .A2(new_n712), .A3(new_n1000), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n260), .B1(new_n724), .B2(new_n372), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n721), .A2(new_n746), .B1(new_n725), .B2(new_n728), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G322), .C2(new_n744), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n738), .A2(G311), .B1(new_n930), .B2(G317), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  OAI22_X1  g0844(.A1(new_n732), .A2(new_n811), .B1(new_n747), .B2(new_n586), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT114), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1042), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n738), .A2(G159), .B1(new_n930), .B2(G150), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT51), .Z(new_n1049));
  INV_X1    g0849(.A(G143), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n354), .A2(new_n732), .B1(new_n743), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G68), .B2(new_n729), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n753), .A2(G77), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n815), .B(new_n767), .C1(new_n287), .C2(new_n720), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1049), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n717), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n769), .A2(new_n246), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n766), .B1(G97), .B2(new_n673), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n714), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1056), .B1(KEYINPUT113), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n764), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1061), .B1(KEYINPUT113), .B2(new_n1060), .C1(new_n962), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1039), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n998), .A2(new_n999), .ZN(new_n1065));
  OAI21_X1  g0865(.A(KEYINPUT109), .B1(new_n992), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n982), .B1(new_n1000), .B2(new_n994), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n995), .A2(new_n1000), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n675), .B1(new_n1069), .B2(new_n982), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1064), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(G390));
  OAI211_X1 g0872(.A(new_n877), .B(new_n879), .C1(new_n842), .C2(new_n890), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n790), .A2(new_n889), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT115), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n790), .A2(KEYINPUT115), .A3(new_n889), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n905), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT116), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n842), .B1(new_n856), .B2(new_n868), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1079), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1073), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n905), .A2(G330), .A3(new_n700), .A4(new_n792), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1073), .B(new_n1084), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n441), .A2(G330), .A3(new_n700), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n896), .A2(new_n1089), .A3(new_n626), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT117), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT117), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n896), .A2(new_n1089), .A3(new_n1092), .A4(new_n626), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n792), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n888), .B1(new_n701), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1096), .A2(new_n1084), .B1(new_n790), .B2(new_n889), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1084), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n701), .A2(KEYINPUT118), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1095), .B1(new_n701), .B2(KEYINPUT118), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n905), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1098), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1094), .A2(KEYINPUT119), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT119), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n701), .A2(KEYINPUT118), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n792), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n888), .B1(new_n1109), .B2(new_n1101), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1085), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1097), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1107), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1088), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1086), .A2(new_n1087), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n674), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1086), .A2(new_n1087), .A3(new_n712), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n713), .B1(new_n287), .B2(new_n796), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n930), .A2(G283), .B1(new_n744), .B2(G294), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n372), .B2(new_n732), .C1(new_n465), .C2(new_n721), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n738), .A2(G116), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n337), .B1(new_n729), .B2(G87), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n799), .A4(new_n1053), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT120), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n720), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n738), .A2(G132), .B1(new_n201), .B2(new_n798), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G128), .A2(new_n930), .B1(new_n805), .B2(G137), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  OR3_X1    g0932(.A1(new_n728), .A2(KEYINPUT53), .A3(new_n928), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n260), .B1(new_n744), .B2(G125), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n753), .A2(G159), .ZN(new_n1135));
  OAI21_X1  g0935(.A(KEYINPUT53), .B1(new_n728), .B2(new_n928), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1123), .A2(new_n1126), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1121), .B1(new_n1138), .B2(new_n716), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n869), .A2(KEYINPUT105), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n879), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(new_n763), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1120), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1119), .A2(new_n1144), .ZN(G378));
  AND3_X1   g0945(.A1(new_n908), .A2(new_n911), .A3(G330), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n880), .B2(new_n894), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1142), .A2(new_n842), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n908), .A2(new_n911), .A3(G330), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1074), .A2(new_n905), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n892), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n890), .A2(KEYINPUT102), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n876), .A3(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1148), .A2(new_n881), .A3(new_n1149), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1147), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n368), .A2(new_n370), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n359), .A2(new_n863), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1158), .B(new_n1159), .Z(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1155), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1147), .A2(new_n1154), .A3(new_n1160), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1160), .A2(new_n762), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n713), .B1(new_n201), .B2(new_n796), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n749), .B1(G33), .B2(G41), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n767), .B2(new_n296), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G97), .A2(new_n805), .B1(new_n744), .B2(G283), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n372), .B2(new_n739), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1170), .A2(G41), .A3(new_n281), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n724), .A2(new_n751), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n734), .A2(new_n586), .B1(new_n728), .B2(new_n340), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n509), .C2(new_n720), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1171), .B(new_n1174), .C1(new_n250), .C2(new_n747), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1168), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G128), .A2(new_n738), .B1(new_n720), .B2(G137), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1128), .A2(new_n729), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n753), .A2(G150), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G125), .A2(new_n930), .B1(new_n805), .B2(G132), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n744), .C2(G124), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n755), .B2(new_n724), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1177), .B1(new_n1176), .B2(new_n1175), .C1(new_n1184), .C2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1166), .B1(new_n1187), .B2(new_n716), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1164), .A2(new_n712), .B1(new_n1165), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1118), .A2(new_n1094), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(KEYINPUT57), .A3(new_n1164), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n674), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1118), .A2(new_n1094), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT57), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1189), .B1(new_n1192), .B2(new_n1194), .ZN(G375));
  NAND2_X1  g0995(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1115), .A2(new_n1003), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT122), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1112), .B2(new_n711), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1105), .A2(KEYINPUT122), .A3(new_n712), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n713), .B1(G68), .B2(new_n796), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n734), .A2(new_n800), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n739), .A2(new_n807), .B1(new_n721), .B2(new_n928), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G159), .C2(new_n729), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n753), .A2(G50), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1172), .B(new_n767), .C1(G128), .C2(new_n744), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1128), .A2(new_n805), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n721), .A2(new_n372), .B1(new_n746), .B2(new_n734), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G116), .B2(new_n805), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT123), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n927), .A2(new_n1019), .A3(new_n337), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G97), .A2(new_n729), .B1(new_n744), .B2(G303), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n725), .C2(new_n739), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1208), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1201), .B1(new_n1215), .B2(new_n716), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n905), .B2(new_n763), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1199), .A2(new_n1200), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1197), .A2(new_n1219), .ZN(G381));
  NAND2_X1  g1020(.A1(new_n1164), .A2(new_n712), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1165), .A2(new_n1188), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n675), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1190), .A2(new_n1164), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1223), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1071), .A2(new_n1231), .A3(new_n825), .ZN(new_n1232));
  OR4_X1    g1032(.A1(G387), .A2(new_n1230), .A3(G381), .A4(new_n1232), .ZN(G407));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1230), .ZN(G409));
  AOI21_X1  g1034(.A(new_n778), .B1(new_n1007), .B2(new_n1037), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n702), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1003), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n711), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n971), .A2(new_n961), .A3(new_n972), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(new_n973), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G390), .B1(new_n1243), .B2(new_n948), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n948), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1245), .B(new_n1071), .C1(new_n1240), .C2(new_n1242), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1237), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(new_n1071), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1243), .A2(new_n948), .A3(G390), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1236), .A3(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT62), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1190), .A2(new_n1003), .A3(new_n1164), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1254), .A2(new_n1189), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT124), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1119), .A2(new_n1256), .A3(new_n1144), .ZN(new_n1257));
  INV_X1    g1057(.A(G213), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1255), .A2(new_n1257), .B1(new_n1258), .B2(G343), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1254), .A2(new_n1189), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(G378), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G375), .B2(G378), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1260), .B1(new_n1263), .B2(new_n1256), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT126), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1266), .B(new_n1260), .C1(new_n1263), .C2(new_n1256), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1269), .A2(new_n1117), .A3(new_n675), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1112), .A2(new_n1113), .A3(KEYINPUT60), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1218), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(G384), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1253), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n653), .A2(G213), .A3(G2897), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1273), .B(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1265), .A2(new_n1267), .A3(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1254), .A2(new_n1189), .A3(new_n1119), .A4(new_n1144), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n1273), .B(new_n1259), .C1(new_n1280), .C2(KEYINPUT124), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1281), .B2(new_n1253), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1252), .B1(new_n1275), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1274), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1247), .A2(new_n1250), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1287), .B(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1264), .B2(new_n1277), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1285), .B(new_n1289), .C1(new_n1281), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1284), .A2(new_n1292), .ZN(G405));
  XNOR2_X1  g1093(.A(new_n1228), .B(G378), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1251), .A2(KEYINPUT127), .B1(new_n1274), .B2(new_n1294), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1294), .A2(new_n1274), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1251), .A2(KEYINPUT127), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1297), .B(new_n1298), .ZN(G402));
endmodule


