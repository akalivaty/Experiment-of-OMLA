//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n195), .B2(new_n189), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G104), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(G104), .A3(new_n197), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n201), .A2(new_n202), .A3(new_n204), .A4(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n198), .A2(new_n206), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G101), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n196), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n207), .A2(new_n209), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n193), .A2(KEYINPUT64), .A3(G143), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n218), .B(KEYINPUT1), .C1(new_n213), .C2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n192), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n210), .B1(new_n211), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(G137), .ZN(new_n228));
  INV_X1    g042(.A(G137), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT11), .A3(G134), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n227), .A2(new_n230), .A3(new_n233), .A4(new_n228), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n224), .A2(KEYINPUT12), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n224), .A2(new_n235), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n224), .A2(KEYINPUT82), .A3(KEYINPUT12), .A4(new_n235), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n211), .A2(new_n223), .A3(new_n244), .A4(KEYINPUT10), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(G128), .A3(new_n219), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n248), .A2(new_n217), .B1(new_n189), .B2(new_n191), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n207), .A2(KEYINPUT10), .A3(new_n209), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT81), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g066(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n253), .A2(new_n203), .B1(G104), .B2(new_n197), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n204), .A2(new_n206), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT80), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n201), .A2(new_n257), .A3(new_n204), .A4(new_n206), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(G101), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n207), .A2(KEYINPUT4), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n256), .A2(new_n262), .A3(G101), .A4(new_n258), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n217), .A2(new_n266), .B1(new_n189), .B2(new_n264), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n235), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT10), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n210), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n252), .A2(new_n268), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G227), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n273), .B(new_n275), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n243), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n252), .A2(new_n268), .A3(new_n271), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n235), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n277), .B1(new_n281), .B2(new_n272), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n187), .B(new_n188), .C1(new_n279), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n272), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n217), .A2(new_n266), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n189), .A2(new_n264), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n259), .B2(new_n260), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n290), .A2(new_n263), .B1(new_n270), .B2(new_n210), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n269), .B1(new_n291), .B2(new_n252), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n276), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(new_n272), .A3(new_n277), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT83), .A3(new_n187), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n277), .B1(new_n294), .B2(new_n272), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n278), .A2(new_n292), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n188), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n285), .A2(new_n297), .B1(new_n300), .B2(G469), .ZN(new_n301));
  OAI21_X1  g115(.A(G214), .B1(G237), .B2(G902), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n302), .B(KEYINPUT84), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G116), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT66), .B1(new_n305), .B2(G119), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G116), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT2), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G113), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n308), .B2(G116), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n305), .A2(KEYINPUT67), .A3(G119), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n310), .A2(new_n315), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n317), .A2(new_n318), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT68), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n315), .A4(new_n310), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n310), .ZN(new_n325));
  INV_X1    g139(.A(new_n315), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n324), .A2(new_n327), .B1(new_n259), .B2(new_n260), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n321), .A2(KEYINPUT5), .A3(new_n310), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n305), .A2(KEYINPUT5), .A3(G119), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(new_n311), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n320), .A2(new_n323), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n328), .A2(new_n263), .B1(new_n211), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT85), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n333), .A2(new_n336), .B1(KEYINPUT86), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(KEYINPUT6), .A3(new_n334), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n324), .A2(new_n327), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n263), .A3(new_n261), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n332), .A2(new_n211), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n337), .A2(KEYINPUT86), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n335), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n338), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n289), .A2(G125), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(G125), .B2(new_n223), .ZN(new_n348));
  INV_X1    g162(.A(G224), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G953), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G210), .B1(G237), .B2(G902), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n334), .B(KEYINPUT8), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n329), .A2(new_n331), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n324), .A2(new_n211), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n211), .B1(new_n324), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT87), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n360), .B(new_n354), .C1(new_n356), .C2(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT7), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n348), .B1(new_n363), .B2(new_n350), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n350), .A2(new_n363), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n347), .B(new_n365), .C1(G125), .C2(new_n223), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n334), .B2(new_n333), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n352), .A2(new_n353), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n353), .B1(new_n352), .B2(new_n369), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n304), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G221), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n375), .B2(new_n188), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n301), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n235), .A2(new_n267), .ZN(new_n378));
  INV_X1    g192(.A(new_n228), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n226), .A2(G137), .ZN(new_n380));
  OAI21_X1  g194(.A(G131), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n234), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n378), .B1(new_n249), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(new_n340), .ZN(new_n384));
  XOR2_X1   g198(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n385));
  NOR2_X1   g199(.A1(G237), .A2(G953), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G210), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n385), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT26), .B(G101), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n388), .B(new_n389), .Z(new_n390));
  NOR2_X1   g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT70), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n320), .A2(new_n323), .B1(new_n326), .B2(new_n325), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n383), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n378), .B(KEYINPUT30), .C1(new_n249), .C2(new_n382), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT69), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n382), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n223), .A2(new_n399), .B1(new_n235), .B2(new_n267), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT69), .B1(new_n400), .B2(KEYINPUT30), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n392), .B(new_n395), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n397), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(KEYINPUT69), .A3(KEYINPUT30), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n392), .B1(new_n406), .B2(new_n395), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n391), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT31), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT28), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n383), .A2(new_n340), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n400), .A2(new_n393), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT28), .B1(new_n400), .B2(new_n393), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n390), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT31), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n416), .B(new_n391), .C1(new_n403), .C2(new_n407), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n409), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G472), .A2(G902), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT32), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT72), .B1(new_n413), .B2(new_n414), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n400), .A2(new_n393), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT28), .B1(new_n384), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT72), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n390), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n428), .A2(KEYINPUT29), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n188), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT73), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n433), .A3(new_n188), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n412), .B(new_n390), .C1(new_n403), .C2(new_n407), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n428), .B1(new_n413), .B2(new_n414), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT29), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G472), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n418), .A2(KEYINPUT32), .A3(new_n419), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n422), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G137), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n274), .A2(G221), .A3(G234), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT74), .B1(new_n190), .B2(G119), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT74), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n308), .A3(G128), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n446), .B(new_n448), .C1(new_n308), .C2(G128), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT24), .B(G110), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT16), .ZN(new_n454));
  INV_X1    g268(.A(G140), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(G125), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(G125), .ZN(new_n457));
  INV_X1    g271(.A(G125), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G140), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n456), .B1(new_n460), .B2(new_n454), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(G146), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n464), .A2(new_n308), .A3(G128), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n190), .A2(G119), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT23), .B1(new_n190), .B2(G119), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G110), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n453), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n461), .A2(new_n193), .ZN(new_n472));
  INV_X1    g286(.A(new_n460), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n193), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n468), .A2(new_n469), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n449), .A2(new_n450), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT76), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT76), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n445), .B1(new_n471), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n453), .A2(new_n463), .A3(new_n470), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n444), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n486), .A3(new_n188), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT25), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G217), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(G234), .B2(new_n188), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n483), .A2(new_n486), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n495), .B(KEYINPUT77), .Z(new_n496));
  NOR2_X1   g310(.A1(new_n493), .A2(G902), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT78), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n386), .A2(G143), .A3(G214), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(G143), .B1(new_n386), .B2(G214), .ZN(new_n504));
  OAI21_X1  g318(.A(G131), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n233), .A3(new_n502), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT91), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n502), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT17), .A3(G131), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n511), .A2(new_n462), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n513), .B(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n460), .A2(KEYINPUT88), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n460), .A2(KEYINPUT88), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(G146), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n474), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G113), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT90), .B(G104), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n515), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n505), .A2(new_n507), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n518), .A2(KEYINPUT19), .A3(new_n519), .ZN(new_n528));
  OR3_X1    g342(.A1(new_n460), .A2(KEYINPUT89), .A3(KEYINPUT19), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT89), .B1(new_n460), .B2(KEYINPUT19), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n472), .B(new_n527), .C1(new_n531), .C2(G146), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n525), .B1(new_n532), .B2(new_n522), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n535));
  NOR2_X1   g349(.A1(G475), .A2(G902), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n526), .A2(new_n533), .ZN(new_n538));
  INV_X1    g352(.A(new_n536), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT20), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n525), .B1(new_n515), .B2(new_n522), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n188), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT92), .B(new_n188), .C1(new_n526), .C2(new_n542), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(G475), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G122), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT93), .B1(new_n549), .B2(G116), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n305), .A3(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n553), .A2(KEYINPUT14), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n553), .A2(KEYINPUT14), .B1(G116), .B2(new_n549), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n197), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n549), .A2(G116), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n197), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G128), .B(G143), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n559), .A2(G134), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(G134), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n190), .A2(G143), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(G134), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n559), .A2(new_n565), .A3(G134), .A4(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(new_n558), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n197), .B1(new_n553), .B2(new_n557), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n374), .A2(new_n492), .A3(G953), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n563), .A2(new_n571), .A3(new_n573), .ZN(new_n576));
  AOI21_X1  g390(.A(G902), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G478), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT15), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n577), .B(new_n579), .Z(new_n580));
  NAND2_X1  g394(.A1(G234), .A2(G237), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(G952), .A3(new_n274), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(KEYINPUT94), .Z(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT21), .B(G898), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(G902), .A3(G953), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n584), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n548), .A2(new_n580), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n377), .A2(new_n441), .A3(new_n501), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  INV_X1    g405(.A(new_n588), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n304), .B(new_n592), .C1(new_n370), .C2(new_n371), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n578), .A2(new_n188), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n577), .B2(new_n578), .ZN(new_n595));
  INV_X1    g409(.A(new_n576), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n573), .B1(new_n563), .B2(new_n571), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT33), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n575), .A2(new_n599), .A3(new_n576), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(G478), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n541), .B2(new_n547), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n593), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n285), .A2(new_n297), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n300), .A2(G469), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n376), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n418), .A2(new_n188), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n609), .A2(G472), .B1(new_n419), .B2(new_n418), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n605), .A2(new_n608), .A3(new_n610), .A4(new_n501), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND3_X1  g427(.A1(new_n580), .A2(new_n547), .A3(new_n541), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n593), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n615), .A2(new_n608), .A3(new_n610), .A4(new_n501), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT95), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n484), .A2(new_n485), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n445), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n498), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n494), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n493), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n489), .B2(new_n490), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n623), .A2(new_n498), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT96), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n377), .A2(new_n589), .A3(new_n610), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  NAND2_X1  g448(.A1(new_n441), .A2(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n352), .A2(new_n369), .ZN(new_n636));
  INV_X1    g450(.A(new_n353), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n352), .A2(new_n369), .A3(new_n353), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n303), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n583), .B1(G900), .B2(new_n586), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n614), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n608), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT97), .B(G128), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G30));
  XOR2_X1   g461(.A(new_n641), .B(KEYINPUT39), .Z(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n608), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n370), .A2(new_n371), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT38), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n548), .A2(new_n580), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n654), .A2(new_n494), .A3(new_n304), .A4(new_n624), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n428), .A2(new_n384), .A3(new_n424), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n412), .B1(new_n403), .B2(new_n407), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(new_n428), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n188), .B1(new_n660), .B2(new_n661), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n440), .A3(new_n422), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n651), .A2(new_n656), .A3(new_n657), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  NAND4_X1  g481(.A1(new_n625), .A2(new_n629), .A3(new_n603), .A4(new_n641), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n377), .A2(new_n441), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n377), .A2(new_n441), .A3(new_n669), .A4(KEYINPUT99), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  NOR2_X1   g489(.A1(new_n279), .A2(new_n282), .ZN(new_n676));
  OAI211_X1 g490(.A(KEYINPUT100), .B(G469), .C1(new_n676), .C2(G902), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n296), .B2(new_n187), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n376), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n606), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n441), .A2(new_n683), .A3(new_n605), .A4(new_n501), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND4_X1  g500(.A1(new_n441), .A2(new_n683), .A3(new_n615), .A4(new_n501), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT101), .B(G116), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G18));
  NAND3_X1  g503(.A1(new_n441), .A2(new_n589), .A3(new_n631), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n682), .B2(new_n372), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n679), .A2(new_n677), .B1(new_n285), .B2(new_n297), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(KEYINPUT102), .A3(new_n681), .A4(new_n640), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n690), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n308), .ZN(G21));
  AND3_X1   g510(.A1(new_n640), .A2(new_n592), .A3(new_n654), .ZN(new_n697));
  INV_X1    g511(.A(G472), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n418), .B2(new_n188), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n423), .A2(new_n427), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n409), .B(new_n417), .C1(new_n428), .C2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n699), .B1(new_n419), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n697), .A2(new_n683), .A3(new_n702), .A4(new_n501), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  NAND2_X1  g518(.A1(new_n692), .A2(new_n694), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n494), .A2(new_n624), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n603), .A2(new_n641), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n702), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  NOR2_X1   g525(.A1(new_n283), .A2(new_n284), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT83), .B1(new_n296), .B2(new_n187), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n607), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n370), .A2(new_n371), .A3(new_n303), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n681), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(KEYINPUT103), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n608), .B2(new_n715), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n440), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n418), .A2(KEYINPUT104), .A3(KEYINPUT32), .A4(new_n419), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n422), .A3(new_n439), .A4(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n501), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n707), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n720), .A2(new_n725), .A3(new_n726), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n716), .A2(KEYINPUT103), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n608), .A2(new_n718), .A3(new_n715), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n724), .A2(new_n501), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT105), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n436), .A2(new_n437), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n432), .B(new_n434), .C1(new_n735), .C2(KEYINPUT29), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n736), .A2(G472), .B1(new_n420), .B2(new_n421), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n500), .B1(new_n737), .B2(new_n440), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n730), .A3(new_n708), .A4(new_n731), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n729), .A2(new_n734), .B1(new_n727), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n233), .ZN(G33));
  NAND3_X1  g555(.A1(new_n720), .A2(new_n738), .A3(new_n643), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  INV_X1    g557(.A(new_n602), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n541), .A3(new_n547), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT43), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT43), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n610), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT44), .A4(new_n706), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n746), .B1(new_n548), .B2(new_n602), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT43), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n420), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n706), .B1(new_n758), .B2(new_n699), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n752), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n751), .A2(new_n760), .A3(new_n715), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n187), .A2(new_n188), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n276), .B1(new_n243), .B2(new_n286), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n281), .A2(new_n272), .A3(new_n277), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(KEYINPUT45), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n298), .B2(new_n299), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n768), .A3(G469), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n766), .A2(KEYINPUT106), .A3(new_n768), .A4(G469), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n762), .B(new_n763), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n606), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT107), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n763), .B1(new_n771), .B2(new_n772), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(new_n606), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n761), .A2(new_n781), .A3(new_n681), .A4(new_n649), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n681), .ZN(new_n784));
  NOR2_X1   g598(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n715), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n441), .A2(new_n788), .A3(new_n501), .A4(new_n707), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n787), .B(new_n789), .C1(new_n784), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  XNOR2_X1  g607(.A(new_n693), .B(KEYINPUT49), .ZN(new_n794));
  INV_X1    g608(.A(new_n665), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n500), .A2(new_n745), .A3(new_n376), .A4(new_n303), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n653), .A4(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT110), .Z(new_n798));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n645), .B1(new_n672), .B2(new_n673), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n640), .A2(new_n654), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n494), .A2(new_n624), .A3(new_n641), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n802), .A2(new_n376), .A3(new_n301), .A4(new_n803), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n705), .A2(new_n709), .B1(new_n804), .B2(new_n665), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n800), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n668), .B1(new_n737), .B2(new_n440), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT99), .B1(new_n808), .B2(new_n377), .ZN(new_n809));
  INV_X1    g623(.A(new_n673), .ZN(new_n810));
  OAI22_X1  g624(.A1(new_n809), .A2(new_n810), .B1(new_n635), .B2(new_n644), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n804), .A2(new_n665), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n710), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n807), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n801), .A2(KEYINPUT114), .A3(new_n805), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n806), .B1(new_n816), .B2(new_n800), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n729), .A2(new_n734), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n739), .A2(new_n727), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n441), .A2(new_n501), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n608), .A2(new_n640), .A3(new_n589), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n611), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n590), .A2(KEYINPUT111), .A3(new_n611), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n632), .A2(new_n703), .A3(new_n616), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n684), .A2(new_n687), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n828), .A2(new_n695), .A3(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n548), .A2(new_n580), .A3(new_n642), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT112), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n635), .A2(new_n832), .A3(new_n716), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n720), .A2(new_n709), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n742), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n820), .A2(new_n827), .A3(new_n830), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n828), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n695), .A2(new_n829), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n827), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(KEYINPUT113), .A3(new_n820), .A4(new_n835), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n817), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n742), .A2(new_n833), .A3(new_n834), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n841), .A2(new_n740), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n801), .A2(KEYINPUT114), .A3(new_n805), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT114), .B1(new_n801), .B2(new_n805), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n800), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n814), .A2(KEYINPUT52), .A3(new_n815), .ZN(new_n852));
  AND4_X1   g666(.A1(KEYINPUT53), .A2(new_n848), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n799), .B1(new_n846), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n749), .A2(new_n584), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n683), .A2(new_n715), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n733), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT48), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n702), .A2(new_n501), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n705), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT118), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n274), .A2(G952), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n857), .A2(new_n665), .A3(new_n500), .A4(new_n583), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n603), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n860), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(new_n547), .A3(new_n541), .A4(new_n602), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT117), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n702), .A2(new_n706), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n858), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n304), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n653), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n862), .A2(new_n683), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n870), .A2(new_n880), .A3(KEYINPUT51), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n693), .A2(new_n376), .ZN(new_n882));
  INV_X1    g696(.A(new_n787), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n784), .A2(new_n791), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n856), .A2(new_n861), .A3(new_n788), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n868), .B1(new_n881), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n870), .A2(new_n880), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n883), .B2(new_n884), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n787), .B(KEYINPUT115), .C1(new_n784), .C2(new_n791), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n892), .A3(new_n882), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n889), .B1(new_n893), .B2(new_n886), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n888), .B1(new_n894), .B2(KEYINPUT51), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n845), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n836), .A2(new_n845), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n817), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n897), .A2(new_n899), .A3(new_n799), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n855), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n798), .B1(new_n901), .B2(new_n902), .ZN(G75));
  NAND2_X1  g717(.A1(new_n897), .A2(new_n899), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(G210), .A3(G902), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n346), .B(KEYINPUT119), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n351), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n274), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(new_n763), .B(KEYINPUT57), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n799), .B1(new_n897), .B2(new_n899), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n900), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n676), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n904), .A2(G902), .A3(new_n771), .A4(new_n772), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n912), .B1(new_n918), .B2(new_n919), .ZN(G54));
  AND2_X1   g734(.A1(KEYINPUT58), .A2(G475), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n904), .A2(G902), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n538), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n922), .B2(new_n538), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n904), .A2(G902), .A3(new_n534), .A4(new_n921), .ZN(new_n926));
  INV_X1    g740(.A(new_n912), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(G60));
  NAND2_X1  g743(.A1(new_n598), .A2(new_n600), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n896), .A2(new_n845), .B1(new_n898), .B2(new_n817), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n799), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n853), .B1(new_n845), .B2(new_n844), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n799), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n594), .B(KEYINPUT59), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n930), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n598), .B2(new_n600), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n900), .B2(new_n915), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n927), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n937), .A2(new_n940), .ZN(G63));
  XNOR2_X1  g755(.A(new_n496), .B(KEYINPUT122), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n492), .A2(new_n188), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n942), .B1(new_n931), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n904), .A2(new_n623), .A3(new_n945), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n948), .A3(new_n927), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT61), .A4(new_n927), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G66));
  NAND2_X1  g767(.A1(new_n841), .A2(new_n274), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT123), .Z(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n585), .B2(new_n349), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n907), .B1(G898), .B2(new_n274), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G69));
  NOR2_X1   g773(.A1(new_n733), .A2(new_n802), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n781), .A2(new_n681), .A3(new_n960), .A4(new_n649), .ZN(new_n961));
  AND4_X1   g775(.A1(new_n820), .A2(new_n792), .A3(new_n742), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n801), .A2(new_n710), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n782), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(KEYINPUT127), .A3(new_n782), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n962), .A2(new_n969), .A3(new_n274), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n406), .B1(KEYINPUT30), .B2(new_n400), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(new_n531), .ZN(new_n972));
  NAND2_X1  g786(.A1(G900), .A2(G953), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  INV_X1    g790(.A(new_n666), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n963), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n801), .A2(new_n666), .A3(KEYINPUT62), .A4(new_n710), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n792), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n788), .B1(new_n604), .B2(new_n614), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n738), .A2(new_n982), .A3(new_n608), .A4(new_n649), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n782), .A2(KEYINPUT124), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT124), .B1(new_n782), .B2(new_n983), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n975), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n986), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n984), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(KEYINPUT125), .A3(new_n792), .A4(new_n980), .ZN(new_n991));
  AOI21_X1  g805(.A(G953), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n974), .B1(new_n992), .B2(new_n972), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n274), .B1(G227), .B2(G900), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n974), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  OAI221_X1 g811(.A(new_n974), .B1(new_n995), .B2(new_n994), .C1(new_n992), .C2(new_n972), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n997), .A2(new_n998), .ZN(G72));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n962), .A2(new_n969), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n842), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n927), .B1(new_n1004), .B2(new_n436), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n659), .A2(new_n428), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n988), .A2(new_n842), .A3(new_n991), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n1001), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1006), .A2(new_n436), .A3(new_n1001), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n933), .A2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1005), .A2(new_n1008), .A3(new_n1010), .ZN(G57));
endmodule


