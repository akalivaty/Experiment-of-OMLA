//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G113), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G113), .A3(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n464), .B(new_n466), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G137), .B1(G101), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n472), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n480), .B1(new_n469), .B2(G2105), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT69), .Z(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n463), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n473), .B2(new_n474), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n485), .A2(new_n487), .B1(G124), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n483), .A2(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G138), .B(new_n488), .C1(new_n467), .C2(new_n468), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n494), .A2(new_n495), .A3(G138), .A4(new_n488), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n488), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n489), .A2(G126), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(G62), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n508), .A2(new_n518), .A3(G62), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n513), .B1(new_n520), .B2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  OR2_X1    g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n524), .A2(new_n525), .B1(new_n506), .B2(new_n507), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n526), .A2(G89), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n510), .A2(KEYINPUT71), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n524), .A2(new_n533), .A3(new_n525), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n532), .A2(G51), .A3(G543), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT72), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(KEYINPUT72), .A3(new_n536), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n531), .B1(new_n538), .B2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n521), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n526), .A2(G90), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n532), .A2(G52), .A3(G543), .A4(new_n534), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND3_X1  g122(.A1(new_n532), .A2(G543), .A3(new_n534), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G43), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n521), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n526), .A2(G81), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n532), .A2(G53), .A3(G543), .A4(new_n534), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT73), .B(G65), .Z(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(new_n508), .ZN(new_n563));
  INV_X1    g138(.A(G78), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n564), .B2(new_n505), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(G91), .B2(new_n526), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n506), .A2(new_n569), .A3(new_n507), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n526), .A2(G87), .B1(G651), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n532), .A2(G49), .A3(G543), .A4(new_n534), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  OAI21_X1  g148(.A(G61), .B1(new_n514), .B2(new_n515), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G48), .A2(G543), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(G651), .B1(new_n510), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n508), .A2(new_n510), .A3(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT74), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n526), .A2(new_n581), .A3(G86), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(G305));
  XOR2_X1   g158(.A(KEYINPUT75), .B(G85), .Z(new_n584));
  NAND2_X1  g159(.A1(new_n526), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n585), .B1(new_n586), .B2(new_n521), .C1(new_n548), .C2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NOR2_X1   g164(.A1(G301), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n549), .A2(G54), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n508), .A2(new_n510), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n521), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n591), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT76), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n590), .B1(new_n601), .B2(new_n589), .ZN(G284));
  AOI21_X1  g177(.A(new_n590), .B1(new_n601), .B2(new_n589), .ZN(G321));
  NAND2_X1  g178(.A1(G299), .A2(new_n589), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n589), .B2(G168), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(new_n589), .B2(G168), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n601), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND3_X1  g183(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n607), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT77), .ZN(new_n611));
  MUX2_X1   g186(.A(new_n609), .B(new_n611), .S(G868), .Z(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n494), .A2(new_n476), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n489), .A2(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n488), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n479), .A2(new_n481), .ZN(new_n624));
  INV_X1    g199(.A(G135), .ZN(new_n625));
  OAI221_X1 g200(.A(new_n621), .B1(new_n622), .B2(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT80), .B(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n619), .A2(new_n620), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(KEYINPUT14), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT81), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n634), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n642), .A2(new_n645), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  INV_X1    g232(.A(new_n650), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n657), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n521), .B1(new_n517), .B2(new_n519), .ZN(new_n681));
  OAI21_X1  g256(.A(G16), .B1(new_n681), .B2(new_n512), .ZN(new_n682));
  INV_X1    g257(.A(G1971), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G22), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G6), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(G16), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G305), .B2(G16), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AOI211_X1 g267(.A(new_n688), .B(new_n690), .C1(G305), .C2(G16), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n686), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n682), .A2(new_n685), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G1971), .ZN(new_n696));
  AND4_X1   g271(.A1(G49), .A2(new_n532), .A3(G543), .A4(new_n534), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n570), .A2(G651), .ZN(new_n698));
  INV_X1    g273(.A(G87), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n593), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(G16), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n684), .A2(G23), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n703), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n684), .B1(new_n571), .B2(new_n572), .ZN(new_n706));
  INV_X1    g281(.A(new_n702), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n696), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n680), .B1(new_n694), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n689), .B(new_n691), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n704), .A2(new_n708), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n683), .B1(new_n682), .B2(new_n685), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n711), .A2(new_n714), .A3(KEYINPUT86), .A4(new_n686), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(new_n717), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT84), .B(G29), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n489), .A2(G119), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n488), .A2(G107), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n482), .A2(KEYINPUT85), .A3(G131), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n728));
  INV_X1    g303(.A(G131), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n624), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n726), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n722), .B1(new_n731), .B2(new_n721), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n734), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n684), .A2(G24), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G290), .B2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1986), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n735), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(KEYINPUT87), .B1(new_n720), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT34), .B1(new_n710), .B2(new_n715), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n743), .A2(new_n744), .A3(new_n740), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n719), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT88), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(new_n719), .C1(new_n742), .C2(new_n745), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n747), .A2(KEYINPUT89), .A3(KEYINPUT36), .A4(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G32), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G105), .ZN(new_n756));
  INV_X1    g331(.A(new_n476), .ZN(new_n757));
  INV_X1    g332(.A(G129), .ZN(new_n758));
  INV_X1    g333(.A(new_n489), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n755), .B1(new_n756), .B2(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G141), .B2(new_n482), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n752), .B1(new_n761), .B2(new_n751), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT27), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(KEYINPUT27), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G1996), .ZN(new_n766));
  INV_X1    g341(.A(G1996), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n763), .A2(new_n767), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n684), .A2(G5), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G301), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT97), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT30), .B(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n775), .A2(new_n751), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G34), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(KEYINPUT24), .ZN(new_n780));
  INV_X1    g355(.A(new_n721), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(KEYINPUT24), .B2(new_n779), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n780), .B1(new_n782), .B2(KEYINPUT95), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(KEYINPUT95), .B2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(G160), .A2(G29), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G2084), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n778), .B1(new_n626), .B2(new_n721), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n772), .B2(new_n771), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G19), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n554), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT92), .B(G1341), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n774), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n781), .A2(G35), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G162), .B2(new_n781), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT29), .ZN(new_n797));
  INV_X1    g372(.A(G2090), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n786), .A2(new_n787), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT98), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n488), .A2(G103), .A3(G2104), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT25), .Z(new_n803));
  AOI22_X1  g378(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n804));
  INV_X1    g379(.A(G139), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n803), .B1(new_n488), .B2(new_n804), .C1(new_n624), .C2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G33), .B(new_n806), .S(G29), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2072), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n781), .A2(G27), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n781), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2078), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n801), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n769), .A2(new_n794), .A3(new_n799), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n684), .A2(G21), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G168), .B2(new_n684), .ZN(new_n815));
  INV_X1    g390(.A(G1966), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n684), .A2(G20), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT23), .Z(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G299), .B2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1956), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n721), .A2(G26), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT28), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n482), .A2(G140), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n489), .A2(G128), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n488), .A2(G116), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n825), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(G29), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT94), .ZN(new_n833));
  INV_X1    g408(.A(G2067), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(G4), .A2(G16), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT90), .Z(new_n837));
  INV_X1    g412(.A(new_n601), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n684), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT91), .B(G1348), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NOR4_X1   g416(.A1(new_n813), .A2(new_n822), .A3(new_n835), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n750), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT89), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n746), .B2(KEYINPUT36), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n746), .B2(KEYINPUT88), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n845), .B1(new_n749), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n843), .A2(new_n848), .ZN(G311));
  OAI21_X1  g424(.A(KEYINPUT99), .B1(new_n843), .B2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n749), .ZN(new_n851));
  INV_X1    g426(.A(new_n845), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n750), .A4(new_n842), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n850), .A2(new_n855), .ZN(G150));
  NAND2_X1  g431(.A1(new_n508), .A2(G67), .ZN(new_n857));
  NAND2_X1  g432(.A1(G80), .A2(G543), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n521), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT100), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(new_n593), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT101), .B(G55), .Z(new_n863));
  OAI22_X1  g438(.A1(new_n859), .A2(KEYINPUT100), .B1(new_n548), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n867), .A3(new_n609), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n554), .A2(KEYINPUT102), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n609), .A2(new_n867), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n870), .A3(new_n865), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n601), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT104), .ZN(new_n879));
  AOI21_X1  g454(.A(G860), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n866), .A2(G860), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT37), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(G145));
  NAND2_X1  g459(.A1(new_n489), .A2(G130), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n488), .A2(G118), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  INV_X1    g462(.A(G142), .ZN(new_n888));
  OAI221_X1 g463(.A(new_n885), .B1(new_n886), .B2(new_n887), .C1(new_n624), .C2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n617), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n731), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT105), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT105), .B1(new_n493), .B2(new_n496), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n501), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n831), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n806), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(new_n761), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n761), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n892), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n626), .B(G160), .Z(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(G162), .Z(new_n903));
  NOR2_X1   g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n898), .A2(new_n899), .A3(new_n892), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n903), .B1(new_n901), .B2(new_n905), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g487(.A1(new_n866), .A2(new_n589), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n611), .B(new_n872), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n591), .A2(new_n599), .A3(new_n597), .ZN(new_n915));
  NAND2_X1  g490(.A1(G299), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n600), .A2(new_n561), .A3(new_n566), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  OR3_X1    g495(.A1(G299), .A2(new_n915), .A3(KEYINPUT107), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(KEYINPUT107), .A3(new_n917), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT41), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(KEYINPUT41), .B2(new_n918), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n920), .B1(new_n914), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(G303), .B(G305), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  OR2_X1    g502(.A1(G290), .A2(G288), .ZN(new_n928));
  NAND2_X1  g503(.A1(G290), .A2(G288), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n926), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n930), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n926), .A3(KEYINPUT108), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n934), .A2(KEYINPUT109), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT109), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n935), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(KEYINPUT42), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n925), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n913), .B1(new_n942), .B2(new_n589), .ZN(G295));
  OAI21_X1  g518(.A(new_n913), .B1(new_n942), .B2(new_n589), .ZN(G331));
  NAND2_X1  g519(.A1(G301), .A2(KEYINPUT110), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n542), .A2(new_n545), .A3(new_n946), .A4(new_n543), .ZN(new_n947));
  INV_X1    g522(.A(new_n539), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n947), .B(new_n530), .C1(new_n948), .C2(new_n537), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  NAND3_X1  g526(.A1(G168), .A2(new_n951), .A3(new_n947), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n945), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n868), .A2(new_n871), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n952), .A3(new_n945), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n956), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n872), .B1(new_n958), .B2(new_n953), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n919), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n957), .A2(new_n959), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n924), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n936), .A2(new_n937), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n964), .B(new_n965), .C1(new_n963), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n957), .A2(new_n959), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n918), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n924), .A2(new_n957), .A3(new_n959), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n909), .B1(new_n970), .B2(new_n938), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT41), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n921), .B2(new_n922), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(new_n918), .B2(new_n972), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AOI211_X1 g551(.A(new_n974), .B(new_n972), .C1(new_n921), .C2(new_n922), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT113), .B1(new_n978), .B2(new_n967), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(KEYINPUT112), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n973), .B2(new_n975), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n957), .A4(new_n959), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n983), .A3(new_n968), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n971), .B1(new_n938), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n966), .B(KEYINPUT44), .C1(new_n985), .C2(new_n965), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n938), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(new_n964), .A3(new_n965), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT43), .B1(new_n971), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI211_X1 g569(.A(KEYINPUT114), .B(KEYINPUT44), .C1(new_n989), .C2(new_n991), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n986), .B1(new_n994), .B2(new_n995), .ZN(G397));
  XOR2_X1   g571(.A(KEYINPUT119), .B(G8), .Z(new_n997));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n497), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT105), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n1001), .B2(new_n501), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n472), .A2(G40), .A3(new_n477), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n997), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n510), .A2(new_n577), .ZN(new_n1006));
  INV_X1    g581(.A(new_n575), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n508), .B2(G61), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1006), .B(new_n579), .C1(new_n1008), .C2(new_n521), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(G1981), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n578), .A2(new_n1012), .A3(new_n580), .A4(new_n582), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(new_n1009), .B2(G1981), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1005), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n997), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1009), .A2(G1981), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT121), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(KEYINPUT49), .A3(new_n1013), .A4(new_n1011), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n895), .A2(new_n1021), .A3(new_n1003), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1016), .A2(new_n1017), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT122), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT122), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1004), .A2(new_n1025), .A3(new_n1020), .A4(new_n1016), .ZN(new_n1026));
  AOI211_X1 g601(.A(G1976), .B(G288), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1013), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1004), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n895), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n502), .A2(new_n1021), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1034), .A3(new_n1003), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n683), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1384), .B1(new_n497), .B2(new_n501), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1003), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1002), .B2(new_n1037), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1036), .A2(KEYINPUT117), .B1(new_n798), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(new_n1042), .A3(new_n683), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1030), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G303), .A2(G8), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT55), .Z(new_n1046));
  NOR2_X1   g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT45), .B1(new_n895), .B2(new_n1021), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1003), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n816), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n895), .A2(new_n1037), .A3(new_n1021), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n472), .A2(G40), .A3(new_n477), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1032), .B2(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1053), .A3(new_n787), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1017), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(G286), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1022), .B(new_n1017), .C1(new_n1058), .C2(G288), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1976), .B1(new_n571), .B2(new_n572), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT120), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1059), .A2(new_n1066), .A3(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1057), .A2(new_n1063), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT63), .B1(new_n1047), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1036), .A2(KEYINPUT117), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1040), .A2(new_n798), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1043), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(G8), .A3(new_n1046), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1044), .A2(KEYINPUT118), .A3(new_n1046), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1037), .B1(new_n895), .B2(new_n1021), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1003), .B1(new_n1032), .B2(KEYINPUT50), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT123), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1052), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1081), .B(new_n1082), .C1(new_n1002), .C2(new_n1037), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1083), .A3(new_n798), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n997), .B1(new_n1084), .B2(new_n1036), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(new_n1046), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1056), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1076), .A2(new_n1077), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1029), .B(new_n1070), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1063), .B(new_n1068), .C1(new_n1085), .C2(new_n1046), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT118), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT126), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1093), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1035), .A2(G2078), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1040), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1102), .A2(new_n1103), .B1(new_n772), .B2(new_n1104), .ZN(new_n1105));
  OR4_X1    g680(.A1(new_n1103), .A2(new_n1048), .A3(new_n1049), .A4(G2078), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(G301), .B(KEYINPUT54), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1048), .A2(new_n1103), .A3(G2078), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1052), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1107), .A2(new_n1108), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1030), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G168), .A2(new_n997), .ZN(new_n1114));
  OAI221_X1 g689(.A(KEYINPUT51), .B1(new_n1113), .B2(new_n1114), .C1(new_n1056), .C2(G168), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(KEYINPUT51), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1056), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n840), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n1121));
  AND4_X1   g696(.A1(new_n1021), .A2(new_n895), .A3(new_n834), .A4(new_n1003), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n915), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1002), .A2(new_n834), .A3(new_n1003), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT60), .B(new_n1127), .C1(new_n1040), .C2(new_n1119), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n600), .B1(new_n1128), .B2(KEYINPUT125), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1125), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1121), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1022), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1035), .B2(G1996), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n554), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT59), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G299), .B(KEYINPUT57), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT56), .B(G2072), .Z(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1031), .A2(new_n1034), .A3(new_n1003), .A4(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1142));
  OAI22_X1  g717(.A1(KEYINPUT124), .A2(new_n1141), .B1(new_n1142), .B2(G1956), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(KEYINPUT124), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1138), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1141), .A2(KEYINPUT124), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1142), .A2(G1956), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1138), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1144), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1146), .A2(new_n1150), .A3(KEYINPUT61), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1132), .A2(new_n1137), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1146), .B1(new_n600), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1150), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1118), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1091), .B1(new_n1101), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT62), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1056), .A2(G168), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT51), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1117), .B(KEYINPUT62), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1107), .A2(G171), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1161), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(KEYINPUT126), .B(new_n1092), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1099), .B1(new_n1098), .B2(new_n1093), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1101), .A2(KEYINPUT127), .A3(new_n1167), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1160), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1048), .A2(new_n1003), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1175), .A2(G1996), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT116), .ZN(new_n1177));
  INV_X1    g752(.A(new_n761), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(G1996), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n831), .B(new_n834), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n1177), .A2(new_n1178), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1175), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n731), .B(new_n734), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1182), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(G290), .A2(G1986), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT115), .Z(new_n1188));
  AND2_X1   g763(.A1(G290), .A2(G1986), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1183), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1174), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1177), .B(KEYINPUT46), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1180), .A2(new_n761), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1193), .B1(new_n1175), .B2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT47), .ZN(new_n1196));
  INV_X1    g771(.A(new_n731), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1182), .A2(new_n734), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n831), .A2(G2067), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1183), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1188), .A2(new_n1183), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT48), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1186), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1196), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1192), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g781(.A1(G401), .A2(new_n460), .A3(G227), .A4(G229), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n1208), .A2(new_n911), .A3(new_n992), .ZN(G225));
  INV_X1    g783(.A(G225), .ZN(G308));
endmodule


