//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n209), .B1(new_n212), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XNOR2_X1  g0032(.A(G50), .B(G68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  XOR2_X1   g0034(.A(G58), .B(G77), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  XOR2_X1   g0040(.A(KEYINPUT8), .B(G58), .Z(new_n241));
  INV_X1    g0041(.A(G20), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n242), .A2(G1), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  OR2_X1    g0045(.A1(new_n245), .A2(KEYINPUT76), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n210), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n252), .B1(new_n245), .B2(KEYINPUT76), .ZN(new_n253));
  INV_X1    g0053(.A(new_n251), .ZN(new_n254));
  INV_X1    g0054(.A(new_n241), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n246), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G58), .ZN(new_n257));
  INV_X1    g0057(.A(G68), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(G20), .B1(new_n259), .B2(new_n201), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G159), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT7), .B1(new_n268), .B2(new_n242), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  AOI211_X1 g0070(.A(new_n270), .B(G20), .C1(new_n265), .C2(new_n267), .ZN(new_n271));
  OAI21_X1  g0071(.A(G68), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT75), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n263), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n270), .B1(new_n275), .B2(G20), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n242), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n258), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT75), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT16), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n263), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n272), .A2(KEYINPUT16), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n248), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n256), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT18), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n265), .A2(new_n267), .A3(G226), .A4(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n265), .A2(new_n267), .A3(G223), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G87), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT77), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n211), .B2(new_n295), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  INV_X1    g0102(.A(G45), .ZN(new_n303));
  AOI21_X1  g0103(.A(G1), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n299), .A2(G232), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT77), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n290), .A2(new_n306), .A3(new_n291), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n293), .A2(new_n294), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n292), .A2(new_n305), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n284), .A2(new_n285), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n256), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT16), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n281), .B1(new_n278), .B2(KEYINPUT75), .ZN(new_n317));
  AOI211_X1 g0117(.A(new_n273), .B(new_n258), .C1(new_n276), .C2(new_n277), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n278), .A2(new_n263), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n249), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT18), .B1(new_n322), .B2(new_n312), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n304), .A2(new_n296), .A3(G274), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n225), .B2(new_n298), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(G190), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n293), .A2(new_n307), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n309), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n256), .B(new_n331), .C1(new_n280), .C2(new_n283), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n322), .A2(KEYINPUT17), .A3(new_n331), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n275), .A2(G232), .A3(new_n287), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n275), .A2(G238), .A3(G1698), .ZN(new_n340));
  INV_X1    g0140(.A(G107), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n339), .B(new_n340), .C1(new_n341), .C2(new_n275), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n342), .A2(KEYINPUT66), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n296), .B1(new_n342), .B2(KEYINPUT66), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G244), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n325), .B1(new_n346), .B2(new_n298), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT67), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n251), .B(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n248), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(G77), .A3(new_n244), .ZN(new_n353));
  INV_X1    g0153(.A(G13), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(G1), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(new_n350), .A3(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(G77), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n241), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n264), .A2(G20), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT15), .B(G87), .Z(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n360), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n359), .B1(new_n365), .B2(new_n248), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n349), .A2(new_n310), .B1(new_n353), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n347), .B1(new_n343), .B2(new_n344), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n294), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n353), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n368), .B2(G190), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n349), .A2(G200), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n254), .A2(new_n248), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n243), .A2(new_n202), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(new_n202), .B2(new_n254), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n241), .A2(new_n361), .B1(G150), .B2(new_n261), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n203), .A2(G20), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n378), .B1(new_n381), .B2(new_n249), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n275), .A2(G1698), .ZN(new_n383));
  XOR2_X1   g0183(.A(KEYINPUT65), .B(G223), .Z(new_n384));
  INV_X1    g0184(.A(G77), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n383), .A2(new_n384), .B1(new_n385), .B2(new_n275), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n275), .A2(G222), .A3(new_n287), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n291), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n299), .A2(G226), .B1(new_n301), .B2(new_n304), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n382), .B1(new_n391), .B2(G169), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n390), .A2(G179), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n375), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT73), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n243), .A2(new_n258), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n352), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n358), .A2(new_n249), .A3(new_n398), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT12), .B1(new_n358), .B2(G68), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT12), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n355), .A2(new_n403), .A3(G20), .A4(new_n258), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n399), .A2(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n261), .A2(G50), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT72), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n362), .A2(new_n385), .B1(new_n242), .B2(G68), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n248), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT11), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT11), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(new_n248), .C1(new_n407), .C2(new_n408), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n405), .A2(new_n413), .A3(KEYINPUT74), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT74), .B1(new_n405), .B2(new_n413), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n296), .A2(G238), .A3(new_n297), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n325), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT71), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT71), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n325), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n275), .A2(G232), .A3(G1698), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n275), .A2(G226), .A3(new_n287), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT70), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT70), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G33), .A3(G97), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n291), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n424), .A2(new_n425), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n425), .B1(new_n424), .B2(new_n434), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n418), .B(G169), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n437), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(G179), .A3(new_n435), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n435), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n418), .B1(new_n442), .B2(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n417), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n436), .A2(new_n437), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G190), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(G200), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n447), .C1(new_n415), .C2(new_n416), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(KEYINPUT9), .B(new_n378), .C1(new_n381), .C2(new_n249), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n388), .A2(G190), .A3(new_n389), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT9), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n249), .B1(new_n379), .B2(new_n380), .ZN(new_n453));
  INV_X1    g0253(.A(new_n378), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT68), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n390), .B2(G200), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n390), .A2(new_n457), .A3(G200), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT10), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n450), .A2(new_n451), .A3(new_n455), .A4(KEYINPUT69), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n462), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(new_n459), .A3(new_n460), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR4_X1   g0267(.A1(new_n338), .A2(new_n396), .A3(new_n449), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n303), .A2(G1), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G257), .A3(new_n296), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(G274), .A3(new_n296), .A4(new_n470), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n265), .A2(new_n267), .A3(G244), .A4(new_n287), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n479), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n275), .A2(G244), .A3(new_n287), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n275), .A2(G250), .A3(G1698), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n480), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  AOI211_X1 g0285(.A(KEYINPUT80), .B(new_n477), .C1(new_n485), .C2(new_n291), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n291), .ZN(new_n488));
  INV_X1    g0288(.A(new_n477), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G190), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n486), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G200), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  AND2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G97), .A2(G107), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n341), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n341), .B1(new_n276), .B2(new_n277), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(KEYINPUT78), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT78), .ZN(new_n504));
  AOI211_X1 g0304(.A(new_n504), .B(new_n341), .C1(new_n276), .C2(new_n277), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n248), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n251), .A2(G97), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n249), .B(new_n251), .C1(G1), .C2(new_n264), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n509), .B2(G97), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n494), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n469), .B1(new_n492), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n493), .A2(KEYINPUT80), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n477), .B1(new_n485), .B2(new_n291), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n487), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(G190), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n510), .ZN(new_n517));
  OAI21_X1  g0317(.A(G107), .B1(new_n269), .B2(new_n271), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n504), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n502), .A2(KEYINPUT78), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(new_n501), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n517), .B1(new_n521), .B2(new_n248), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n516), .A2(new_n522), .A3(KEYINPUT81), .A4(new_n494), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n310), .B1(new_n486), .B2(new_n490), .ZN(new_n524));
  AOI211_X1 g0324(.A(G179), .B(new_n477), .C1(new_n485), .C2(new_n291), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n506), .B2(new_n510), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n512), .A2(new_n523), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n265), .A2(new_n267), .A3(G244), .A4(G1698), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n265), .A2(new_n267), .A3(G238), .A4(new_n287), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n291), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n296), .A2(G274), .A3(new_n470), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n250), .A2(G45), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n296), .A2(G250), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n532), .A2(G190), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT84), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n536), .B1(new_n291), .B2(new_n531), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(KEYINPUT84), .A3(G190), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n358), .A2(new_n363), .ZN(new_n544));
  INV_X1    g0344(.A(G87), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n508), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n429), .B2(new_n431), .ZN(new_n548));
  NOR4_X1   g0348(.A1(KEYINPUT82), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT82), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G87), .A2(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(new_n341), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n548), .A2(G20), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n265), .A2(new_n267), .A3(new_n242), .A4(G68), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n554), .A2(KEYINPUT83), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n361), .A2(G97), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n554), .A2(KEYINPUT83), .B1(new_n556), .B2(new_n547), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n544), .B(new_n546), .C1(new_n558), .C2(new_n248), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n532), .A2(new_n537), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n543), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n475), .A2(new_n470), .B1(new_n211), .B2(new_n295), .ZN(new_n563));
  INV_X1    g0363(.A(new_n472), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT5), .A2(G41), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n534), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n563), .A2(G270), .B1(new_n301), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n266), .A2(G33), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n569));
  OAI21_X1  g0369(.A(G303), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n265), .A2(new_n267), .A3(G264), .A4(G1698), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n265), .A2(new_n267), .A3(G257), .A4(new_n287), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n291), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G200), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n250), .B2(G33), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n350), .B1(new_n355), .B2(G20), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n249), .B(new_n578), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n356), .A2(new_n577), .A3(new_n357), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n247), .A2(new_n210), .B1(G20), .B2(new_n577), .ZN(new_n583));
  INV_X1    g0383(.A(G97), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n483), .B(new_n242), .C1(G33), .C2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n583), .A2(KEYINPUT20), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT20), .B1(new_n583), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n581), .B(new_n582), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n576), .B(new_n589), .C1(new_n491), .C2(new_n575), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n341), .A2(KEYINPUT23), .A3(G20), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT23), .B1(new_n341), .B2(G20), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n591), .A2(new_n592), .B1(G20), .B2(new_n530), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n265), .A2(new_n267), .A3(new_n242), .A4(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT22), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT22), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n275), .A2(new_n596), .A3(new_n242), .A4(G87), .ZN(new_n597));
  AOI211_X1 g0397(.A(KEYINPUT24), .B(new_n593), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n597), .ZN(new_n600));
  INV_X1    g0400(.A(new_n593), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n248), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n254), .A2(new_n341), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT25), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(G107), .B2(new_n509), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n265), .A2(new_n267), .A3(G257), .A4(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n265), .A2(new_n267), .A3(G250), .A4(new_n287), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G294), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n291), .B1(new_n563), .B2(G264), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(G190), .A3(new_n476), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n291), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n563), .A2(G264), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n476), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n603), .A2(new_n606), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n558), .A2(new_n248), .ZN(new_n618));
  INV_X1    g0418(.A(new_n544), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n509), .A2(new_n363), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n541), .A2(new_n294), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n560), .A2(new_n310), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n562), .A2(new_n590), .A3(new_n617), .A4(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT85), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n575), .A2(new_n588), .A3(G169), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n588), .A2(G179), .A3(new_n574), .A4(new_n567), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n310), .B1(new_n567), .B2(new_n574), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n627), .B1(new_n631), .B2(new_n588), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n603), .A2(new_n606), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n615), .A2(G179), .ZN(new_n635));
  AOI21_X1  g0435(.A(G169), .B1(new_n611), .B2(new_n476), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n625), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n468), .A2(new_n527), .A3(new_n640), .ZN(G372));
  AND3_X1   g0441(.A1(new_n448), .A2(new_n334), .A3(new_n335), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n444), .A2(new_n370), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n324), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT89), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT89), .B1(new_n464), .B2(new_n466), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n394), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n468), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT86), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n541), .B2(G169), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n560), .A2(KEYINPUT86), .A3(new_n310), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n621), .A2(new_n622), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n562), .A2(new_n654), .A3(new_n617), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n633), .B2(new_n638), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n527), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT87), .B1(new_n526), .B2(new_n524), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n562), .A2(new_n654), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n526), .A2(new_n524), .A3(KEYINPUT87), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT26), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n562), .A2(new_n526), .A3(new_n524), .A4(new_n624), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n664), .A2(KEYINPUT88), .B1(KEYINPUT26), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT88), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n526), .A2(new_n524), .A3(KEYINPUT87), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n669), .A2(new_n660), .A3(new_n661), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n670), .B2(KEYINPUT26), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n659), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n649), .B1(new_n650), .B2(new_n672), .ZN(G369));
  NAND2_X1  g0473(.A1(new_n355), .A2(new_n242), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G343), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n588), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n633), .B(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n590), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n634), .A2(new_n680), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n617), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n638), .ZN(new_n687));
  INV_X1    g0487(.A(new_n638), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n679), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n679), .B1(new_n630), .B2(new_n632), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n689), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(G399));
  OR3_X1    g0496(.A1(new_n549), .A2(new_n552), .A3(G116), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT90), .Z(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n207), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n214), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n654), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n526), .A2(new_n524), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT87), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n562), .A2(new_n654), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n663), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n706), .B1(KEYINPUT26), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT92), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n656), .B1(new_n639), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n633), .A2(new_n638), .A3(KEYINPUT92), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n527), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n679), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT26), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n711), .A2(KEYINPUT88), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT88), .B1(new_n711), .B2(new_n720), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n658), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n679), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT91), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n719), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT29), .B1(new_n726), .B2(KEYINPUT91), .ZN(new_n729));
  INV_X1    g0529(.A(G330), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n575), .A2(new_n294), .A3(new_n560), .ZN(new_n732));
  INV_X1    g0532(.A(new_n615), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n732), .A2(new_n514), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n541), .A2(new_n611), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n567), .A2(new_n574), .A3(G179), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n513), .A2(new_n737), .A3(new_n515), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n513), .A2(new_n737), .A3(KEYINPUT30), .A4(new_n515), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n731), .B(new_n679), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n739), .ZN(new_n743));
  INV_X1    g0543(.A(new_n734), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT31), .B1(new_n745), .B2(new_n680), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n512), .A2(new_n523), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n640), .A2(new_n748), .A3(new_n707), .A4(new_n679), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n730), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n728), .A2(new_n729), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n705), .B1(new_n751), .B2(G1), .ZN(G364));
  INV_X1    g0552(.A(new_n684), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n683), .A2(G330), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n354), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n250), .B1(new_n755), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n701), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n753), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT93), .Z(new_n760));
  OR2_X1    g0560(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n275), .A2(G355), .A3(new_n207), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n236), .A2(new_n303), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n700), .A2(new_n275), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G45), .B2(new_n214), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n764), .B1(G116), .B2(new_n207), .C1(new_n765), .C2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n210), .B1(G20), .B2(new_n310), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n763), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n772), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n491), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n294), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G97), .ZN(new_n780));
  NAND2_X1  g0580(.A1(G20), .A2(G179), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT96), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n329), .A2(G190), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n780), .B1(new_n790), .B2(new_n258), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT101), .Z(new_n792));
  NOR2_X1   g0592(.A1(new_n491), .A2(new_n329), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n784), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G190), .A2(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n784), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G50), .A2(new_n795), .B1(new_n798), .B2(G77), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n242), .A2(G179), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n785), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G107), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n793), .A2(new_n800), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n268), .B1(new_n805), .B2(G87), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n784), .A2(new_n777), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G58), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n799), .A2(new_n803), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n800), .A2(new_n796), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT97), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT97), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G159), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT98), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT32), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n810), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT33), .B(G317), .Z(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n790), .A2(new_n821), .B1(new_n822), .B2(new_n807), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT102), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n275), .B1(new_n805), .B2(G303), .ZN(new_n825));
  INV_X1    g0625(.A(G294), .ZN(new_n826));
  INV_X1    g0626(.A(new_n779), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G311), .B2(new_n798), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G329), .A2(new_n815), .B1(new_n802), .B2(G283), .ZN(new_n830));
  INV_X1    g0630(.A(G326), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n794), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n792), .A2(new_n820), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT103), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n773), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n775), .B1(new_n683), .B2(new_n776), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n760), .A2(new_n838), .ZN(G396));
  NAND3_X1  g0639(.A1(new_n671), .A2(new_n722), .A3(new_n721), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n680), .B1(new_n840), .B2(new_n658), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n371), .A2(new_n680), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n374), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n370), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n370), .A2(new_n680), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n375), .A2(new_n679), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n841), .A2(new_n847), .B1(new_n672), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n750), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n758), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n268), .B1(new_n805), .B2(G50), .ZN(new_n853));
  INV_X1    g0653(.A(new_n802), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n257), .B2(new_n827), .C1(new_n854), .C2(new_n258), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G137), .A2(new_n795), .B1(new_n798), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G143), .ZN(new_n857));
  INV_X1    g0657(.A(G150), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n856), .B1(new_n857), .B2(new_n807), .C1(new_n790), .C2(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT34), .Z(new_n860));
  AOI211_X1 g0660(.A(new_n855), .B(new_n860), .C1(G132), .C2(new_n815), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n275), .B1(new_n805), .B2(G107), .ZN(new_n862));
  INV_X1    g0662(.A(G303), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n780), .B(new_n862), .C1(new_n794), .C2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n815), .A2(G311), .B1(new_n798), .B2(G116), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n802), .A2(G87), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n826), .C2(new_n807), .ZN(new_n867));
  INV_X1    g0667(.A(new_n790), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n864), .B(new_n867), .C1(G283), .C2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n773), .B1(new_n861), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n773), .A2(new_n770), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n763), .B1(new_n385), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n870), .B(new_n872), .C1(new_n847), .C2(new_n771), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n852), .A2(new_n873), .ZN(G384));
  OAI21_X1  g0674(.A(new_n332), .B1(new_n322), .B2(new_n312), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n322), .A2(new_n677), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n284), .A2(new_n313), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n284), .A2(new_n678), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n332), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n876), .B1(new_n324), .B2(new_n336), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n316), .B1(new_n278), .B2(new_n263), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n282), .A2(new_n887), .A3(new_n248), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n677), .B1(new_n888), .B2(new_n256), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n324), .B2(new_n336), .ZN(new_n890));
  INV_X1    g0690(.A(new_n332), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n312), .A2(new_n677), .B1(new_n888), .B2(new_n256), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n890), .A2(KEYINPUT38), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT39), .B1(new_n886), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n890), .A2(KEYINPUT38), .A3(new_n894), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n890), .B2(new_n894), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT14), .B1(new_n445), .B2(new_n310), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n440), .A3(new_n438), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n417), .A3(new_n679), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n901), .A2(new_n905), .B1(new_n324), .B2(new_n677), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT106), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n405), .A2(new_n413), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT74), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n414), .A3(new_n680), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT105), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n910), .A2(new_n913), .A3(new_n414), .A4(new_n680), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n444), .A2(new_n448), .A3(new_n912), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n903), .A2(new_n417), .A3(new_n680), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n898), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n895), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n848), .B1(new_n840), .B2(new_n658), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n917), .B(new_n919), .C1(new_n920), .C2(new_n846), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n906), .A2(new_n907), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n918), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n882), .B2(new_n883), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n897), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n905), .C1(new_n925), .C2(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n324), .A2(new_n677), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n921), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT106), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n649), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT29), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n841), .B2(new_n727), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n680), .B1(new_n712), .B2(new_n716), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n841), .B2(KEYINPUT91), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n932), .B1(new_n938), .B2(new_n468), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n931), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n745), .A2(new_n680), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n731), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n749), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n917), .A3(new_n847), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n925), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT108), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n944), .A2(new_n917), .A3(new_n847), .A4(KEYINPUT108), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(new_n919), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n947), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n468), .A2(new_n944), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n730), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n940), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n958), .A2(KEYINPUT109), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(KEYINPUT109), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n940), .A2(new_n957), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n755), .A2(new_n250), .ZN(new_n962));
  NOR4_X1   g0762(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n212), .A2(new_n577), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n500), .B(KEYINPUT104), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT35), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT36), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n214), .A2(new_n385), .A3(new_n259), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n202), .A2(G68), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n250), .B(G13), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n963), .A2(new_n970), .A3(new_n973), .ZN(G367));
  OR2_X1    g0774(.A1(new_n522), .A2(new_n679), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n527), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT110), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n527), .A2(KEYINPUT110), .A3(new_n975), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n707), .B1(new_n980), .B2(new_n638), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n526), .A2(new_n524), .A3(new_n680), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(new_n982), .A3(new_n979), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n690), .A2(new_n693), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n981), .A2(new_n679), .B1(KEYINPUT42), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(KEYINPUT42), .B2(new_n985), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n559), .A2(new_n679), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n710), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n654), .B2(new_n988), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n987), .A2(KEYINPUT43), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n691), .A2(new_n983), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n987), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n991), .A2(new_n992), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n992), .B1(new_n991), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n701), .B(KEYINPUT41), .Z(new_n1000));
  NAND2_X1  g0800(.A1(new_n983), .A2(new_n695), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT45), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n978), .A2(new_n694), .A3(new_n982), .A4(new_n979), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n691), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT45), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1001), .B(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1003), .B(KEYINPUT44), .Z(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n1008), .A3(new_n692), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n690), .B(new_n693), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(KEYINPUT111), .B2(new_n684), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n684), .B(KEYINPUT111), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n1010), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1005), .A2(new_n751), .A3(new_n1009), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1000), .B1(new_n1014), .B2(new_n751), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT112), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n756), .B1(new_n1015), .B2(KEYINPUT112), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n999), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n231), .A2(new_n766), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n774), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n700), .B2(new_n363), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n763), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(G283), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n797), .A2(new_n1023), .B1(new_n341), .B2(new_n827), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT113), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n868), .A2(G294), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT46), .B1(new_n805), .B2(G116), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n268), .C1(new_n584), .C2(new_n801), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G303), .A2(new_n808), .B1(new_n795), .B2(G311), .ZN(new_n1031));
  INV_X1    g0831(.A(G317), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n814), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(G159), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n790), .A2(new_n1035), .B1(new_n202), .B2(new_n797), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT114), .Z(new_n1037));
  AOI22_X1  g0837(.A1(new_n815), .A2(G137), .B1(new_n795), .B2(G143), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n858), .B2(new_n807), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n827), .A2(new_n258), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n801), .A2(new_n385), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n275), .B1(new_n804), .B2(new_n257), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1034), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n773), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1022), .B1(new_n776), .B2(new_n990), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1018), .A2(new_n1047), .ZN(G387));
  NAND2_X1  g0848(.A1(new_n690), .A2(new_n772), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n763), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n698), .A2(new_n207), .A3(new_n275), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(G107), .B2(new_n207), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n699), .A2(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n699), .A2(KEYINPUT115), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n241), .A2(new_n202), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n1056), .C1(G68), .C2(G77), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1053), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n700), .B(new_n275), .C1(new_n228), .C2(G45), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1052), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1050), .B1(new_n1060), .B2(new_n1020), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n808), .A2(G50), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n779), .A2(new_n363), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n805), .A2(G77), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1062), .A2(new_n275), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G97), .A2(new_n802), .B1(new_n798), .B2(G68), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n858), .B2(new_n814), .C1(new_n1035), .C2(new_n794), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(new_n241), .C2(new_n868), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT116), .Z(new_n1069));
  INV_X1    g0869(.A(new_n801), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n275), .B1(new_n1070), .B2(G116), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n827), .A2(new_n1023), .B1(new_n804), .B2(new_n826), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G317), .A2(new_n808), .B1(new_n795), .B2(G322), .ZN(new_n1073));
  INV_X1    g0873(.A(G311), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1073), .B1(new_n863), .B2(new_n797), .C1(new_n790), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT48), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT49), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1071), .B1(new_n831), .B2(new_n814), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1069), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1061), .B1(new_n1082), .B2(new_n773), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1013), .A2(new_n757), .B1(new_n1049), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n751), .A2(new_n1013), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n701), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n751), .A2(new_n1013), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(G393));
  NAND2_X1  g0888(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1085), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n701), .A3(new_n1014), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1005), .A2(new_n757), .A3(new_n1009), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n239), .A2(new_n766), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1093), .B(new_n774), .C1(new_n584), .C2(new_n207), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1074), .A2(new_n807), .B1(new_n794), .B2(new_n1032), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n814), .A2(new_n822), .B1(new_n797), .B2(new_n826), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n275), .B1(new_n805), .B2(G283), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n803), .B(new_n1098), .C1(new_n577), .C2(new_n827), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1097), .B(new_n1099), .C1(new_n868), .C2(G303), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n814), .A2(new_n857), .B1(new_n797), .B2(new_n255), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n268), .B1(new_n805), .B2(G68), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n866), .B(new_n1102), .C1(new_n385), .C2(new_n827), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n868), .C2(G50), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n858), .A2(new_n794), .B1(new_n807), .B2(new_n1035), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT51), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1096), .A2(new_n1100), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1050), .B(new_n1094), .C1(new_n1107), .C2(new_n1046), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT117), .Z(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n776), .B2(new_n983), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1091), .A2(new_n1092), .A3(new_n1110), .ZN(G390));
  OAI21_X1  g0911(.A(new_n468), .B1(new_n728), .B2(new_n729), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n917), .B1(new_n750), .B2(new_n847), .ZN(new_n1113));
  AND4_X1   g0913(.A1(G330), .A2(new_n944), .A3(new_n847), .A4(new_n917), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1113), .A2(new_n1114), .B1(new_n920), .B2(new_n846), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n944), .A2(new_n847), .A3(G330), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n917), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT118), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n846), .B1(new_n935), .B2(new_n844), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n750), .A2(new_n847), .A3(new_n917), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1115), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n650), .A2(new_n850), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1112), .A2(new_n1124), .A3(new_n649), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT119), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n917), .B1(new_n920), .B2(new_n846), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n901), .B1(new_n1129), .B2(new_n904), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n886), .A2(new_n895), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1131), .B(new_n904), .C1(new_n1120), .C2(new_n1117), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1114), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n672), .A2(new_n848), .B1(new_n370), .B2(new_n680), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n905), .B1(new_n1135), .B2(new_n917), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1132), .B(new_n1121), .C1(new_n1136), .C2(new_n901), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT119), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n939), .A2(new_n1139), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1128), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1128), .A2(new_n1138), .A3(new_n1140), .A4(KEYINPUT120), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n650), .B1(new_n934), .B2(new_n937), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1146), .A2(new_n932), .A3(new_n1125), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n1134), .A3(new_n1137), .A4(new_n1124), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1148), .A2(new_n701), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n763), .B1(new_n255), .B2(new_n871), .ZN(new_n1151));
  OR3_X1    g0951(.A1(new_n804), .A2(KEYINPUT53), .A3(new_n858), .ZN(new_n1152));
  OAI21_X1  g0952(.A(KEYINPUT53), .B1(new_n804), .B2(new_n858), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n1035), .C2(new_n827), .ZN(new_n1154));
  XOR2_X1   g0954(.A(KEYINPUT54), .B(G143), .Z(new_n1155));
  AOI22_X1  g0955(.A1(G132), .A2(new_n808), .B1(new_n798), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n794), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1154), .B(new_n1158), .C1(G137), .C2(new_n868), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n275), .B1(new_n801), .B2(new_n202), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n815), .B2(G125), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT121), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n868), .A2(G107), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n854), .A2(new_n258), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n577), .A2(new_n807), .B1(new_n794), .B2(new_n1023), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n814), .A2(new_n826), .B1(new_n797), .B2(new_n584), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n268), .B1(new_n804), .B2(new_n545), .C1(new_n827), .C2(new_n385), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1159), .A2(new_n1162), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1151), .B1(new_n1046), .B2(new_n1169), .C1(new_n901), .C2(new_n771), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1138), .B2(new_n756), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1150), .A2(new_n1172), .ZN(G378));
  NAND2_X1  g0973(.A1(new_n951), .A2(new_n953), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n947), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(G330), .A3(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n395), .B1(new_n646), .B2(new_n647), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n382), .A2(new_n678), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1178), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1184), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n1182), .A3(new_n1177), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1176), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n954), .B2(G330), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n907), .B1(new_n906), .B2(new_n921), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n907), .A2(new_n921), .A3(new_n927), .A4(new_n926), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1190), .A2(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1176), .A2(new_n1189), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n954), .A2(G330), .A3(new_n1188), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1195), .A2(new_n922), .A3(new_n930), .A4(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1194), .A2(new_n1197), .A3(KEYINPUT57), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT123), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1148), .A2(new_n1199), .A3(new_n1147), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1148), .B2(new_n1147), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1147), .B1(new_n1138), .B2(new_n1127), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT123), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1148), .A2(new_n1199), .A3(new_n1147), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1203), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n701), .B(new_n1202), .C1(new_n1207), .C2(KEYINPUT57), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1203), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1189), .A2(new_n770), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n871), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n758), .B1(new_n1211), .B2(G50), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n275), .A2(G41), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G50), .B(new_n1213), .C1(new_n264), .C2(new_n302), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G116), .A2(new_n795), .B1(new_n798), .B2(new_n363), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1023), .B2(new_n814), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1064), .B(new_n1213), .C1(new_n257), .C2(new_n801), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1216), .A2(new_n1040), .A3(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n807), .A2(new_n341), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT122), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n584), .C2(new_n790), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1214), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G128), .A2(new_n808), .B1(new_n798), .B2(G137), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n795), .A2(G125), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n779), .A2(G150), .B1(new_n805), .B2(new_n1155), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G132), .B2(new_n868), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n815), .A2(G124), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G33), .B(G41), .C1(new_n1070), .C2(G159), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT59), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1231), .B(new_n1232), .C1(new_n1228), .C2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1223), .B1(new_n1222), .B2(new_n1221), .C1(new_n1230), .C2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1212), .B1(new_n1235), .B2(new_n773), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1209), .A2(new_n757), .B1(new_n1210), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1208), .A2(new_n1237), .ZN(G375));
  AOI21_X1  g1038(.A(new_n275), .B1(new_n805), .B2(G97), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1063), .B(new_n1239), .C1(new_n807), .C2(new_n1023), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G107), .A2(new_n798), .B1(new_n795), .B2(G294), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n385), .B2(new_n854), .C1(new_n863), .C2(new_n814), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(G116), .C2(new_n868), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n268), .B1(new_n1070), .B2(G58), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n1035), .B2(new_n804), .C1(new_n202), .C2(new_n827), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n815), .A2(G128), .B1(new_n795), .B2(G132), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G137), .A2(new_n808), .B1(new_n798), .B2(G150), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1245), .B(new_n1248), .C1(new_n868), .C2(new_n1155), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n773), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n1050), .C1(G68), .C2(new_n1211), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1117), .B2(new_n770), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1124), .B2(new_n757), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1147), .A2(KEYINPUT124), .A3(new_n1124), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1112), .A2(new_n649), .A3(new_n1126), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1124), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1000), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1128), .A2(new_n1261), .A3(new_n1140), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1253), .B1(new_n1260), .B2(new_n1262), .ZN(G381));
  OR4_X1    g1063(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1264), .A2(G387), .A3(G381), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1171), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1208), .A4(new_n1237), .ZN(G407));
  INV_X1    g1067(.A(G213), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(G343), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G375), .C2(new_n1270), .ZN(G409));
  NAND3_X1  g1071(.A1(new_n1208), .A2(G378), .A3(new_n1237), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1209), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1237), .B1(new_n1273), .B2(new_n1000), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1266), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1269), .ZN(new_n1277));
  INV_X1    g1077(.A(G384), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n701), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1127), .A2(KEYINPUT60), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1259), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1253), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1278), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1258), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1256), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1282), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1281), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(G384), .A3(new_n1253), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1285), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1276), .A2(new_n1277), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1269), .A2(G2897), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1285), .B2(new_n1291), .ZN(new_n1297));
  INV_X1    g1097(.A(G2897), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1277), .B1(KEYINPUT126), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(KEYINPUT126), .B2(new_n1298), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1285), .A2(new_n1291), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1285), .A2(new_n1291), .A3(KEYINPUT127), .A4(new_n1300), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1297), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1295), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1269), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n1292), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1294), .A2(new_n1306), .A3(new_n1307), .A4(new_n1310), .ZN(new_n1311));
  XOR2_X1   g1111(.A(G393), .B(G396), .Z(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1018), .A2(new_n1047), .A3(G390), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G390), .B1(new_n1018), .B2(new_n1047), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(G390), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G387), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1018), .A2(new_n1047), .A3(G390), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1312), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1316), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1311), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1316), .A2(new_n1320), .A3(new_n1307), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1293), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1308), .A2(KEYINPUT63), .A3(new_n1292), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1308), .A2(KEYINPUT125), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1305), .B1(new_n1308), .B2(KEYINPUT125), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1325), .B(new_n1326), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1322), .A2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1266), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1272), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1332), .A2(new_n1292), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1292), .ZN(new_n1334));
  OR3_X1    g1134(.A1(new_n1333), .A2(new_n1334), .A3(new_n1321), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1321), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(G402));
endmodule


