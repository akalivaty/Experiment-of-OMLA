//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2106), .ZN(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(G2104), .ZN(new_n469));
  OAI22_X1  g044(.A1(new_n466), .A2(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  AOI21_X1  g049(.A(new_n465), .B1(new_n462), .B2(new_n463), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n465), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  OAI221_X1 g054(.A(new_n476), .B1(new_n477), .B2(new_n478), .C1(new_n479), .C2(new_n466), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT67), .Z(G162));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n483), .B(KEYINPUT69), .C1(new_n485), .C2(new_n484), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n488), .A2(KEYINPUT70), .A3(KEYINPUT4), .A4(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n465), .B2(G114), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(G126), .B2(new_n475), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n483), .B(new_n499), .C1(new_n485), .C2(new_n484), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n499), .B1(new_n486), .B2(new_n487), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(new_n489), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n498), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT71), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(G543), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(new_n513), .A3(new_n511), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n506), .A2(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(G62), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(KEYINPUT72), .B1(G75), .B2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n510), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n516), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  XNOR2_X1  g097(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n525), .B1(new_n513), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(new_n529), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G51), .A3(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(G89), .A3(new_n513), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n527), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n510), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n530), .A2(G52), .A3(G543), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n530), .A2(G90), .A3(new_n513), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n537), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(KEYINPUT75), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(KEYINPUT75), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(G651), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  INV_X1    g125(.A(new_n512), .ZN(new_n551));
  INV_X1    g126(.A(new_n514), .ZN(new_n552));
  AOI22_X1  g127(.A1(G43), .A2(new_n551), .B1(new_n552), .B2(G81), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT77), .Z(G188));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT78), .B1(new_n514), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n530), .A2(new_n564), .A3(G91), .A4(new_n513), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n512), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n530), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g146(.A(KEYINPUT79), .B(G65), .Z(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(new_n513), .B1(G78), .B2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n510), .B1(new_n573), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n566), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT81), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n568), .A2(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(new_n581), .A3(new_n566), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(new_n542), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n585), .A2(new_n540), .B1(new_n510), .B2(new_n535), .ZN(G301));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n533), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n527), .A2(KEYINPUT82), .A3(new_n531), .A4(new_n532), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G286));
  NAND3_X1  g166(.A1(new_n530), .A2(G49), .A3(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n514), .C2(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(new_n552), .A2(G86), .ZN(new_n596));
  INV_X1    g171(.A(G48), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n510), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n599), .A2(KEYINPUT83), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(KEYINPUT83), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n596), .B1(new_n597), .B2(new_n512), .C1(new_n600), .C2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n552), .A2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n551), .A2(G47), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(new_n510), .C2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n552), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n514), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n512), .A2(new_n613), .B1(new_n510), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n607), .B1(G868), .B2(new_n616), .ZN(G284));
  OAI21_X1  g192(.A(new_n607), .B1(G868), .B2(new_n616), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G286), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(new_n583), .ZN(G297));
  AOI21_X1  g196(.A(new_n620), .B1(new_n619), .B2(new_n583), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT84), .ZN(G148));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n623), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XOR2_X1   g204(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n466), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G135), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n465), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n475), .A2(KEYINPUT86), .A3(G123), .ZN(new_n639));
  AOI21_X1  g214(.A(KEYINPUT86), .B1(new_n475), .B2(G123), .ZN(new_n640));
  OAI221_X1 g215(.A(new_n636), .B1(new_n637), .B2(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n634), .A2(G2100), .B1(new_n641), .B2(G2096), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n642), .B(new_n643), .C1(G2100), .C2(new_n634), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT87), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(G14), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT88), .Z(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT89), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(KEYINPUT17), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n662), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n664), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n669), .A3(new_n662), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g253(.A1(new_n670), .A2(new_n673), .A3(new_n674), .A4(new_n676), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT91), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n684), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(new_n686), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n690), .A3(new_n686), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G1981), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT20), .B1(new_n688), .B2(new_n693), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n695), .A2(new_n700), .A3(new_n685), .A4(new_n687), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n697), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n698), .B1(new_n697), .B2(new_n702), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n683), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n697), .A2(new_n702), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G1981), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n697), .A2(new_n698), .A3(new_n702), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n707), .A2(G1986), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT92), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n705), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n705), .B2(new_n709), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n682), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n703), .A2(new_n704), .A3(new_n683), .ZN(new_n716));
  AOI21_X1  g291(.A(G1986), .B1(new_n707), .B2(new_n708), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n705), .A2(new_n709), .A3(new_n712), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n681), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(G229));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n723), .A2(G6), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G305), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT32), .B(G1981), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT97), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n723), .A2(G23), .ZN(new_n729));
  NAND2_X1  g304(.A1(G288), .A2(KEYINPUT98), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n552), .A2(G87), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT98), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n731), .A2(new_n732), .A3(new_n592), .A4(new_n593), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n729), .B1(new_n734), .B2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT33), .B(G1976), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n728), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n727), .A2(KEYINPUT97), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n735), .A2(new_n737), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n723), .A2(G22), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G166), .B2(new_n723), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1971), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT34), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G25), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n475), .A2(G119), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT93), .Z(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G107), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n635), .B2(G131), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(new_n749), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT94), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n759), .B(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(G16), .A2(G24), .ZN(new_n763));
  XNOR2_X1  g338(.A(G290), .B(KEYINPUT95), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n723), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n762), .B1(new_n766), .B2(G1986), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G1986), .B2(new_n766), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n747), .A2(new_n748), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT36), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT104), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n749), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n749), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT29), .Z(new_n774));
  INV_X1    g349(.A(G2090), .ZN(new_n775));
  INV_X1    g350(.A(G1341), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n555), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G16), .B2(G19), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G4), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n616), .B2(G16), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G1348), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n782), .A2(G1348), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  NAND2_X1  g360(.A1(G164), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G27), .B2(G29), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G29), .A2(G33), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT25), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n635), .A2(G139), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n464), .A2(G127), .ZN(new_n795));
  AND2_X1   g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  OAI21_X1  g371(.A(G2105), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n789), .B1(new_n799), .B2(G29), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G2072), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n749), .A2(G32), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT102), .B(KEYINPUT26), .Z(new_n804));
  NAND3_X1  g379(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G105), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n469), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n475), .A2(G129), .ZN(new_n809));
  INV_X1    g384(.A(G141), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n466), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n803), .B1(new_n812), .B2(new_n749), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT27), .B(G1996), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n801), .A2(new_n802), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G2084), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n749), .ZN(new_n820));
  INV_X1    g395(.A(G160), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n749), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n816), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n723), .A2(G21), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G168), .B2(new_n723), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(G1966), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(G1966), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n823), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT31), .B(G11), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT30), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(G28), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n749), .B1(new_n831), .B2(G28), .ZN(new_n833));
  OAI221_X1 g408(.A(new_n830), .B1(new_n832), .B2(new_n833), .C1(new_n641), .C2(new_n749), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n817), .B2(new_n822), .ZN(new_n835));
  OAI221_X1 g410(.A(new_n835), .B1(new_n802), .B2(new_n801), .C1(new_n813), .C2(new_n815), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n787), .A2(new_n785), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT100), .B(KEYINPUT28), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n749), .A2(G26), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n475), .A2(G128), .ZN(new_n841));
  INV_X1    g416(.A(G140), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n466), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n844));
  OR3_X1    g419(.A1(KEYINPUT99), .A2(G104), .A3(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT99), .B1(G104), .B2(G2105), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n840), .B1(new_n848), .B2(new_n749), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G2067), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n836), .A2(new_n837), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n780), .A2(new_n788), .A3(new_n829), .A4(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT103), .B(KEYINPUT23), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n723), .A2(G20), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n583), .B2(new_n723), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G1956), .ZN(new_n857));
  NOR2_X1   g432(.A1(G171), .A2(new_n723), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G5), .B2(new_n723), .ZN(new_n859));
  INV_X1    g434(.A(G1961), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n778), .A2(new_n776), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n774), .A2(new_n775), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n861), .B(new_n862), .C1(new_n860), .C2(new_n859), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n852), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n770), .A2(new_n771), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n771), .B1(new_n770), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(G311));
  NAND2_X1  g442(.A1(new_n770), .A2(new_n864), .ZN(G150));
  NAND4_X1  g443(.A1(new_n509), .A2(G55), .A3(G543), .A4(new_n511), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n513), .A2(G67), .ZN(new_n870));
  NAND2_X1  g445(.A1(G80), .A2(G543), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G651), .ZN(new_n873));
  INV_X1    g448(.A(G93), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n869), .B(new_n873), .C1(new_n514), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT105), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(G860), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n554), .A2(new_n876), .ZN(new_n879));
  INV_X1    g454(.A(new_n875), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n549), .A2(new_n550), .A3(new_n553), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT38), .Z(new_n883));
  INV_X1    g458(.A(new_n616), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(new_n623), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n883), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT106), .Z(new_n889));
  INV_X1    g464(.A(G860), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n887), .B2(KEYINPUT39), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n878), .B1(new_n889), .B2(new_n891), .ZN(G145));
  XNOR2_X1  g467(.A(new_n480), .B(KEYINPUT67), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G160), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n641), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n475), .A2(G130), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n465), .A2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(G142), .B2(new_n635), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n632), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n758), .ZN(new_n902));
  INV_X1    g477(.A(new_n812), .ZN(new_n903));
  NAND2_X1  g478(.A1(G164), .A2(new_n848), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n843), .A2(new_n847), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n504), .B2(new_n498), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n906), .A3(new_n798), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n798), .B1(new_n904), .B2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n812), .A3(new_n907), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n902), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n895), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n912), .ZN(new_n915));
  INV_X1    g490(.A(new_n902), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n913), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(KEYINPUT107), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n921), .A3(new_n916), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n918), .B1(new_n923), .B2(new_n895), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g500(.A(new_n882), .B(new_n626), .Z(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n580), .A2(new_n581), .A3(new_n566), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n581), .B1(new_n580), .B2(new_n566), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n579), .A2(KEYINPUT108), .A3(new_n582), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n884), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n583), .A2(new_n927), .A3(new_n616), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT41), .B1(new_n932), .B2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n926), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n933), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n939), .B2(new_n926), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n734), .B(G305), .ZN(new_n942));
  XOR2_X1   g517(.A(G303), .B(G290), .Z(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n944), .A2(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n941), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n941), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n876), .A2(new_n619), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(G295));
  NAND2_X1  g526(.A1(G295), .A2(KEYINPUT110), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(G331));
  NAND2_X1  g530(.A1(new_n590), .A2(G171), .ZN(new_n956));
  NAND2_X1  g531(.A1(G301), .A2(new_n533), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n882), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n879), .A3(new_n881), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n935), .A2(new_n961), .A3(new_n936), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n958), .A2(new_n960), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n938), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n944), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT41), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n938), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n967), .A3(new_n934), .ZN(new_n968));
  INV_X1    g543(.A(new_n944), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n939), .A2(new_n961), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G37), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n965), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n970), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n975), .B2(new_n944), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n977), .A3(new_n971), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(KEYINPUT44), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n977), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n973), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n978), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n979), .B1(new_n983), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n498), .B2(new_n504), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT112), .B(G40), .Z(new_n989));
  NOR3_X1   g564(.A1(new_n988), .A2(new_n821), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n758), .A2(new_n760), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n812), .B(G1996), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n905), .A2(G2067), .ZN(new_n993));
  INV_X1    g568(.A(G2067), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n848), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n758), .A2(new_n760), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n991), .A2(new_n992), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(G290), .B(G1986), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n821), .A2(new_n989), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT45), .B(new_n985), .C1(new_n498), .C2(new_n504), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n988), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1001), .B1(new_n1004), .B2(G2078), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1007), .B(new_n985), .C1(new_n498), .C2(new_n504), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1002), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT121), .B(G1961), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n988), .A2(new_n1003), .ZN(new_n1012));
  NAND4_X1  g587(.A1(G160), .A2(KEYINPUT53), .A3(G40), .A4(new_n785), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1005), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G171), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n785), .A2(KEYINPUT53), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1004), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT122), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n1011), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1005), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT54), .B(new_n1015), .C1(new_n1021), .C2(G171), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n596), .B1(new_n597), .B2(new_n512), .ZN(new_n1023));
  OAI21_X1  g598(.A(G1981), .B1(new_n1023), .B2(new_n599), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(G305), .B2(G1981), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n986), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1002), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1024), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n730), .A2(new_n733), .A3(G1976), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT114), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(G8), .B(new_n1029), .C1(new_n1033), .C2(KEYINPUT114), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1033), .A2(KEYINPUT114), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(new_n1034), .A3(new_n1030), .A4(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1032), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G303), .A2(G8), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1043), .B(KEYINPUT55), .Z(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT113), .B(G1971), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n1004), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(G2090), .B2(new_n1009), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1044), .A2(G8), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1044), .B1(G8), .B2(new_n1047), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1042), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1022), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1021), .A2(G171), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1014), .A2(G171), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT54), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1966), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1004), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1006), .A2(new_n817), .A3(new_n1002), .A4(new_n1008), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(KEYINPUT117), .A3(new_n1058), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n533), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT118), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1057), .A2(KEYINPUT117), .A3(new_n1058), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT117), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1067));
  OAI21_X1  g642(.A(G168), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1059), .A2(G8), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1059), .A2(KEYINPUT119), .A3(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT51), .B1(new_n533), .B2(G8), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1065), .A2(new_n1070), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1061), .A2(G8), .A3(new_n533), .A4(new_n1062), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1078), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1055), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1055), .B(KEYINPUT123), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1029), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1086), .A2(new_n994), .B1(new_n1009), .B2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(new_n884), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n884), .A2(KEYINPUT60), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1089), .A2(KEYINPUT60), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT56), .B(G2072), .Z(new_n1093));
  OR2_X1    g668(.A1(new_n1004), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1956), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1009), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n578), .B(KEYINPUT57), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1098), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(new_n1096), .A3(new_n1094), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT61), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT58), .B(G1341), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n1086), .A2(new_n1104), .B1(new_n1004), .B2(G1996), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n555), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT59), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1092), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1102), .A2(KEYINPUT61), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1107), .B(new_n1092), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1091), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1088), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1101), .A2(new_n616), .A3(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1116), .A2(new_n1099), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1084), .A2(new_n1085), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1071), .A2(G286), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1050), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT63), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G288), .A2(G1976), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT115), .Z(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G305), .A2(G1981), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1030), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1048), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(new_n1042), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1122), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT62), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1131));
  NOR4_X1   g706(.A1(new_n1052), .A2(new_n1049), .A3(new_n1042), .A4(new_n1048), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1080), .A2(new_n1081), .A3(KEYINPUT62), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1000), .B1(new_n1119), .B2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(G290), .A2(G1986), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n990), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT124), .B(KEYINPUT48), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1140), .B(new_n1141), .C1(new_n990), .C2(new_n998), .ZN(new_n1142));
  INV_X1    g717(.A(new_n996), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n990), .B1(new_n1143), .B2(new_n903), .ZN(new_n1144));
  INV_X1    g719(.A(G1996), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n990), .A2(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1146), .A2(KEYINPUT46), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(KEYINPUT46), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT47), .Z(new_n1150));
  NAND2_X1  g725(.A1(new_n992), .A2(new_n996), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n995), .B1(new_n1151), .B2(new_n997), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1142), .B(new_n1150), .C1(new_n990), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1136), .A2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1156));
  NAND4_X1  g730(.A1(new_n660), .A2(new_n678), .A3(G319), .A4(new_n679), .ZN(new_n1157));
  INV_X1    g731(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n721), .B2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g733(.A(KEYINPUT125), .B(new_n1157), .C1(new_n715), .C2(new_n720), .ZN(new_n1160));
  OAI21_X1  g734(.A(new_n924), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g735(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g736(.A(KEYINPUT126), .B1(new_n982), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1164));
  AOI211_X1 g738(.A(new_n1164), .B(new_n1161), .C1(new_n981), .C2(new_n978), .ZN(new_n1165));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n1166));
  NOR3_X1   g740(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n973), .A2(new_n980), .ZN(new_n1168));
  AOI21_X1  g742(.A(new_n977), .B1(new_n976), .B2(new_n971), .ZN(new_n1169));
  OAI21_X1  g743(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1170), .A2(new_n1164), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n982), .A2(KEYINPUT126), .A3(new_n1162), .ZN(new_n1172));
  AOI21_X1  g746(.A(KEYINPUT127), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g747(.A1(new_n1167), .A2(new_n1173), .ZN(G308));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1172), .ZN(G225));
endmodule


