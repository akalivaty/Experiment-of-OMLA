//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT97), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G128), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT97), .A3(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT13), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n190), .A2(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT98), .ZN(new_n196));
  OAI22_X1  g010(.A1(new_n195), .A2(new_n196), .B1(new_n194), .B2(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(new_n192), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(new_n194), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n198), .A2(new_n196), .A3(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(G134), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT99), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT99), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n203), .B(G134), .C1(new_n197), .C2(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n198), .A2(new_n193), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G134), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G122), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n209), .A2(G122), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n208), .A2(new_n213), .A3(new_n210), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n206), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n202), .A2(new_n204), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n205), .B(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n210), .B1(new_n208), .B2(KEYINPUT14), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n208), .A2(KEYINPUT14), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT100), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT100), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n208), .A2(new_n221), .A3(KEYINPUT14), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n214), .B(new_n217), .C1(new_n223), .C2(new_n213), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT9), .B(G234), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT83), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n226), .A2(new_n227), .A3(G953), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n216), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n216), .B2(new_n224), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n187), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G478), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT15), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(G234), .A2(G237), .ZN(new_n235));
  INV_X1    g049(.A(G953), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n235), .A2(G952), .A3(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n235), .A2(G902), .A3(G953), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT21), .B(G898), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI221_X1 g055(.A(new_n187), .B1(KEYINPUT15), .B2(new_n232), .C1(new_n229), .C2(new_n230), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n234), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G113), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(G104), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n189), .A2(KEYINPUT92), .ZN(new_n247));
  NOR2_X1   g061(.A1(G237), .A2(G953), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n247), .A2(G214), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT92), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n251), .A2(new_n247), .B1(new_n248), .B2(G214), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT18), .A2(G131), .ZN(new_n254));
  XNOR2_X1  g068(.A(G125), .B(G140), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G140), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G125), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G140), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n253), .A2(new_n254), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G214), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n265), .A2(G237), .A3(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n247), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT92), .B(G143), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n254), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n269), .A2(KEYINPUT93), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT93), .B1(new_n269), .B2(new_n270), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n264), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G131), .B1(new_n249), .B2(new_n252), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n267), .B(new_n275), .C1(new_n266), .C2(new_n268), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT17), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT95), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT95), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n274), .A2(new_n276), .A3(new_n280), .A4(new_n277), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT16), .ZN(new_n284));
  OR3_X1    g098(.A1(new_n260), .A2(KEYINPUT16), .A3(G140), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n260), .A2(KEYINPUT16), .A3(G140), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(KEYINPUT78), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n256), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n283), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n255), .B2(KEYINPUT16), .ZN(new_n291));
  OAI211_X1 g105(.A(G146), .B(new_n290), .C1(new_n291), .C2(new_n283), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n269), .A2(KEYINPUT17), .A3(G131), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n246), .B(new_n273), .C1(new_n282), .C2(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT19), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT19), .B1(new_n259), .B2(new_n261), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT94), .B1(new_n298), .B2(G146), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n274), .A2(new_n276), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT94), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n301), .B(new_n256), .C1(new_n296), .C2(new_n297), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n299), .A2(new_n300), .A3(new_n292), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n273), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n246), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n295), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G475), .A2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT96), .B1(new_n295), .B2(new_n306), .ZN(new_n311));
  OAI22_X1  g125(.A1(new_n308), .A2(new_n310), .B1(new_n311), .B2(KEYINPUT20), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT96), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT20), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n310), .B1(new_n295), .B2(new_n306), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n295), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n289), .A2(new_n292), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n319), .A2(new_n279), .A3(new_n293), .A4(new_n281), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n246), .B1(new_n320), .B2(new_n273), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n187), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n312), .A2(new_n317), .B1(G475), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n243), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G221), .B1(new_n226), .B2(G902), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT84), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G469), .ZN(new_n328));
  AND2_X1   g142(.A1(KEYINPUT0), .A2(G128), .ZN(new_n329));
  XNOR2_X1  g143(.A(G143), .B(G146), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(KEYINPUT64), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n256), .A2(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n189), .A2(G146), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT0), .A2(G128), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT64), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT69), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n331), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n331), .B2(new_n338), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT3), .B1(new_n245), .B2(G107), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n213), .A3(G104), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n245), .A2(G107), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT87), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT87), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n343), .A2(new_n345), .A3(new_n349), .A4(new_n346), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(G101), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G101), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n343), .A2(new_n345), .A3(new_n352), .A4(new_n346), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(KEYINPUT4), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n347), .B2(KEYINPUT87), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n350), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n342), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n189), .A2(G146), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n256), .A2(G143), .ZN(new_n361));
  OAI211_X1 g175(.A(G128), .B(new_n359), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n245), .A2(G107), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n213), .A2(G104), .ZN(new_n364));
  OAI21_X1  g178(.A(G101), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n332), .B(new_n333), .C1(KEYINPUT1), .C2(new_n191), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n362), .A2(new_n353), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n367), .A2(KEYINPUT10), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(KEYINPUT10), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n358), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT70), .ZN(new_n372));
  INV_X1    g186(.A(G134), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT65), .B1(new_n373), .B2(G137), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT11), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT11), .ZN(new_n376));
  OAI211_X1 g190(.A(KEYINPUT65), .B(new_n376), .C1(new_n373), .C2(G137), .ZN(new_n377));
  INV_X1    g191(.A(G137), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G134), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AND4_X1   g194(.A1(new_n275), .A2(new_n375), .A3(new_n377), .A4(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n379), .B1(new_n374), .B2(KEYINPUT11), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n275), .B1(new_n382), .B2(new_n377), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n372), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n375), .A2(new_n377), .A3(new_n380), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G131), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n275), .A3(new_n377), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(KEYINPUT70), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n371), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n381), .A2(new_n383), .A3(new_n372), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT70), .B1(new_n386), .B2(new_n387), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n358), .A2(new_n393), .A3(new_n370), .ZN(new_n394));
  XNOR2_X1  g208(.A(G110), .B(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n236), .A2(G227), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n390), .A2(new_n394), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n401));
  INV_X1    g215(.A(new_n367), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n366), .A2(new_n362), .B1(new_n353), .B2(new_n365), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n362), .A2(new_n366), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n353), .A2(new_n365), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT89), .A3(new_n367), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n389), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n386), .B2(new_n387), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n367), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(new_n412), .B2(new_n413), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n331), .A2(new_n338), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT69), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n331), .A2(new_n338), .A3(new_n339), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n419), .A2(new_n357), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n421), .A2(new_n354), .B1(new_n369), .B2(new_n368), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n411), .A2(new_n417), .B1(new_n422), .B2(new_n393), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n400), .B1(new_n423), .B2(new_n399), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n328), .B1(new_n424), .B2(new_n187), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT90), .B(G469), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n401), .A2(new_n413), .B1(new_n384), .B2(new_n388), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT12), .B1(new_n427), .B2(new_n408), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n412), .A2(new_n413), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT88), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n394), .B(new_n399), .C1(new_n428), .C2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n399), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n358), .A2(new_n393), .A3(new_n370), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n393), .B1(new_n358), .B2(new_n370), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(G902), .B(new_n426), .C1(new_n433), .C2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n327), .B1(new_n425), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G214), .B1(G237), .B2(G902), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n209), .A2(G119), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n209), .A2(KEYINPUT68), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G116), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n446), .A3(G119), .ZN(new_n447));
  INV_X1    g261(.A(new_n441), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(G113), .B(new_n443), .C1(new_n449), .C2(new_n442), .ZN(new_n450));
  NOR2_X1   g264(.A1(KEYINPUT2), .A2(G113), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT2), .A2(G113), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n447), .A3(new_n456), .A4(new_n448), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n450), .A2(new_n457), .A3(new_n353), .A4(new_n365), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n457), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n357), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n353), .A2(KEYINPUT4), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n355), .B2(new_n350), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n458), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G122), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n458), .B(new_n466), .C1(new_n462), .C2(new_n464), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n471), .A3(new_n467), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n331), .A2(new_n338), .A3(G125), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n362), .A2(new_n260), .A3(new_n366), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n236), .A2(G224), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n466), .B(KEYINPUT8), .Z(new_n479));
  NAND2_X1  g293(.A1(new_n443), .A2(G113), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n441), .B1(new_n207), .B2(G119), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(KEYINPUT5), .ZN(new_n482));
  INV_X1    g296(.A(new_n457), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n406), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n479), .B1(new_n484), .B2(new_n458), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n476), .A2(KEYINPUT7), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n486), .A2(KEYINPUT91), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(KEYINPUT91), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n475), .B2(new_n489), .ZN(new_n490));
  AOI211_X1 g304(.A(KEYINPUT91), .B(new_n486), .C1(new_n473), .C2(new_n474), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n485), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G902), .B1(new_n492), .B2(new_n469), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n478), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n478), .B2(new_n493), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n440), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n324), .A2(new_n439), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT32), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n248), .A2(G210), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT27), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(G101), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n378), .A3(G134), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT66), .B1(new_n378), .B2(G134), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n373), .A2(G137), .ZN(new_n508));
  OAI211_X1 g322(.A(G131), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n387), .A2(new_n509), .A3(new_n366), .A4(new_n362), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n389), .B2(new_n342), .ZN(new_n512));
  INV_X1    g326(.A(new_n461), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(KEYINPUT28), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n381), .A2(new_n383), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n510), .B1(new_n515), .B2(new_n418), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n461), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n342), .B1(new_n391), .B2(new_n392), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n513), .A3(new_n510), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n504), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n461), .B(new_n511), .C1(new_n389), .C2(new_n342), .ZN(new_n524));
  INV_X1    g338(.A(new_n504), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n386), .A2(new_n387), .ZN(new_n527));
  INV_X1    g341(.A(new_n418), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n509), .A2(new_n362), .A3(new_n366), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n527), .A2(new_n528), .B1(new_n387), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n461), .B1(new_n530), .B2(KEYINPUT30), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n510), .A2(KEYINPUT30), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n389), .B2(new_n342), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n519), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n513), .B1(new_n516), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT71), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n526), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT31), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n534), .B1(new_n531), .B2(new_n533), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n539), .A3(KEYINPUT71), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT31), .A3(new_n526), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n523), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT72), .Z(new_n550));
  OAI21_X1  g364(.A(new_n500), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT29), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n522), .A2(new_n504), .A3(new_n514), .A4(new_n517), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n524), .B1(new_n544), .B2(new_n545), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n552), .B(new_n553), .C1(new_n554), .C2(new_n504), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT73), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n519), .A2(new_n556), .A3(new_n513), .A4(new_n510), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n513), .B2(new_n512), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n512), .B2(new_n513), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT28), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI211_X1 g374(.A(KEYINPUT74), .B(KEYINPUT28), .C1(new_n512), .C2(new_n513), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT74), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n520), .B2(new_n521), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n525), .A2(new_n552), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n555), .A2(new_n566), .A3(new_n187), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G472), .ZN(new_n568));
  INV_X1    g382(.A(new_n522), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n514), .A2(new_n517), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n525), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n520), .A2(new_n504), .ZN(new_n572));
  AOI211_X1 g386(.A(new_n542), .B(new_n572), .C1(new_n544), .C2(new_n545), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT31), .B1(new_n546), .B2(new_n526), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n550), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n551), .A2(new_n568), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n289), .A2(new_n292), .ZN(new_n580));
  INV_X1    g394(.A(G110), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT76), .ZN(new_n582));
  OAI211_X1 g396(.A(G119), .B(new_n191), .C1(new_n582), .C2(KEYINPUT23), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT23), .ZN(new_n584));
  INV_X1    g398(.A(G119), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n585), .B2(G128), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT76), .B1(new_n585), .B2(G128), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT77), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n581), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(KEYINPUT77), .B(new_n583), .C1(new_n586), .C2(new_n587), .ZN(new_n591));
  XNOR2_X1  g405(.A(G119), .B(G128), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT24), .B(G110), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT75), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n592), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n590), .A2(new_n591), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n580), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n593), .A2(new_n594), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n581), .B(new_n583), .C1(new_n586), .C2(new_n587), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n601), .A2(new_n602), .B1(new_n256), .B2(new_n255), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n292), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT22), .B(G137), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n236), .A2(G221), .A3(G234), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(new_n607));
  AND4_X1   g421(.A1(new_n579), .A2(new_n600), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n580), .A2(new_n599), .B1(new_n292), .B2(new_n603), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n579), .B1(new_n609), .B2(new_n607), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n590), .A2(new_n591), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n595), .A2(new_n598), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n604), .B1(new_n319), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT79), .ZN(new_n616));
  INV_X1    g430(.A(new_n607), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT79), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT80), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n616), .A2(KEYINPUT80), .A3(new_n619), .A4(new_n617), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n611), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n227), .B1(G234), .B2(new_n187), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(G902), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n611), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n600), .A2(new_n618), .A3(new_n604), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n618), .B1(new_n600), .B2(new_n604), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT80), .B1(new_n633), .B2(new_n617), .ZN(new_n634));
  INV_X1    g448(.A(new_n623), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n187), .B(new_n630), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT25), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(G902), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n608), .B2(new_n610), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(new_n634), .B2(new_n635), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT82), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n622), .A2(new_n623), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(KEYINPUT82), .A3(new_n641), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n638), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n629), .B1(new_n647), .B2(new_n626), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n499), .A2(new_n578), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G101), .ZN(G3));
  INV_X1    g464(.A(G472), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n575), .B2(new_n187), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n543), .A2(new_n547), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n550), .B1(new_n653), .B2(new_n571), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n440), .B(new_n241), .C1(new_n496), .C2(new_n497), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n439), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n232), .A2(new_n187), .ZN(new_n658));
  INV_X1    g472(.A(new_n230), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n216), .A2(new_n224), .A3(new_n228), .ZN(new_n660));
  AOI21_X1  g474(.A(G902), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n658), .B1(new_n661), .B2(new_n232), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT33), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n659), .A2(new_n663), .A3(new_n660), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT33), .B1(new_n229), .B2(new_n230), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n665), .A3(G478), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n323), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n656), .A2(new_n648), .A3(new_n657), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT34), .B(G104), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  INV_X1    g485(.A(new_n656), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n648), .A2(new_n657), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n234), .A2(new_n242), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n316), .B(new_n315), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n322), .A2(G475), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n672), .A2(new_n673), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT35), .B(G107), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  OR2_X1    g494(.A1(new_n617), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n633), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n628), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT25), .B1(new_n624), .B2(new_n187), .ZN(new_n685));
  AOI211_X1 g499(.A(new_n643), .B(new_n640), .C1(new_n622), .C2(new_n623), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT82), .B1(new_n645), .B2(new_n641), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n626), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n652), .A2(new_n654), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n499), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT101), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n692), .B(new_n694), .ZN(G12));
  NOR2_X1   g509(.A1(new_n439), .A2(new_n498), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n237), .B1(new_n238), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n677), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n690), .A2(new_n578), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G128), .ZN(G30));
  XOR2_X1   g515(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n698), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n657), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT40), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n686), .A2(new_n687), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n689), .B1(new_n706), .B2(new_n638), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n683), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n496), .A2(new_n497), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT38), .Z(new_n710));
  INV_X1    g524(.A(new_n674), .ZN(new_n711));
  INV_X1    g525(.A(new_n440), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n323), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n708), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n558), .A2(new_n504), .A3(new_n559), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(G902), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n554), .A2(new_n525), .ZN(new_n717));
  OAI21_X1  g531(.A(G472), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n551), .A2(new_n577), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n705), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT103), .B(G143), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G45));
  AOI21_X1  g537(.A(new_n316), .B1(new_n314), .B2(new_n315), .ZN(new_n724));
  AND4_X1   g538(.A1(KEYINPUT96), .A2(new_n307), .A3(new_n315), .A4(new_n309), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n676), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n698), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n666), .A3(new_n662), .A4(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n690), .A2(new_n578), .A3(new_n696), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  NAND2_X1  g545(.A1(new_n433), .A2(new_n437), .ZN(new_n732));
  INV_X1    g546(.A(new_n426), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n187), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(G902), .B1(new_n433), .B2(new_n437), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n734), .B(new_n327), .C1(new_n328), .C2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n655), .A2(new_n667), .A3(new_n323), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n578), .A3(new_n648), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NOR2_X1   g556(.A1(new_n655), .A2(new_n677), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n578), .A3(new_n648), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  INV_X1    g559(.A(new_n324), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n736), .A2(new_n498), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n690), .A2(new_n578), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  AOI211_X1 g563(.A(new_n629), .B(new_n240), .C1(new_n647), .C2(new_n626), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n560), .A2(new_n564), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n525), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n550), .B1(new_n752), .B2(new_n653), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n652), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n498), .A2(new_n323), .A3(new_n711), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n750), .A2(new_n738), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n747), .B1(new_n707), .B2(new_n683), .ZN(new_n759));
  INV_X1    g573(.A(new_n753), .ZN(new_n760));
  OAI21_X1  g574(.A(G472), .B1(new_n548), .B2(G902), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n729), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n478), .A2(new_n493), .ZN(new_n764));
  INV_X1    g578(.A(new_n494), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n712), .B1(new_n766), .B2(new_n495), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n735), .A2(new_n328), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n327), .A3(new_n734), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n647), .A2(new_n626), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(new_n684), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n652), .A2(new_n728), .A3(new_n753), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(KEYINPUT105), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n763), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  NAND3_X1  g589(.A1(new_n766), .A2(new_n440), .A3(new_n495), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n728), .A2(new_n439), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n578), .A3(new_n648), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT106), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n777), .A2(new_n578), .A3(new_n648), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n551), .A2(KEYINPUT107), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n551), .A2(KEYINPUT107), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n577), .A3(new_n568), .A4(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(KEYINPUT42), .A3(new_n648), .A4(new_n777), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  NOR2_X1   g603(.A1(new_n439), .A2(new_n776), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n578), .A2(new_n648), .A3(new_n699), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n373), .ZN(G36));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n424), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT108), .B1(new_n424), .B2(new_n793), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n424), .A2(KEYINPUT108), .A3(new_n793), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n328), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n328), .A2(new_n187), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n734), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n327), .A3(new_n703), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT109), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n803), .A2(new_n806), .A3(new_n327), .A4(new_n703), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OAI22_X1  g622(.A1(new_n707), .A2(new_n683), .B1(new_n654), .B2(new_n652), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT111), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n667), .A2(new_n726), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n812), .B2(KEYINPUT43), .ZN(new_n813));
  XNOR2_X1  g627(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n813), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n776), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n816), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT112), .B1(new_n819), .B2(KEYINPUT44), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n816), .A2(new_n821), .A3(new_n817), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n808), .B(new_n818), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  NAND2_X1  g638(.A1(new_n802), .A2(new_n734), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n327), .B1(new_n825), .B2(new_n800), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n803), .A2(KEYINPUT47), .A3(new_n327), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n578), .A2(new_n648), .A3(new_n728), .A4(new_n776), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G140), .ZN(G42));
  NOR4_X1   g647(.A1(new_n667), .A2(new_n726), .A3(new_n326), .A4(new_n712), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n768), .A2(new_n734), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n648), .B(new_n834), .C1(new_n835), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT113), .Z(new_n839));
  AOI21_X1  g653(.A(new_n710), .B1(new_n835), .B2(new_n837), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n720), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n690), .A2(new_n790), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n676), .A2(new_n711), .A3(new_n675), .A4(new_n727), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n578), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n762), .B2(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n791), .B(new_n845), .C1(new_n783), .C2(new_n787), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n711), .B2(new_n726), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n323), .A2(new_n674), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n656), .A2(new_n648), .A3(new_n657), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n692), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n649), .A3(new_n669), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n852), .B1(new_n851), .B2(new_n692), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n756), .A2(new_n740), .A3(new_n744), .A4(new_n748), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n759), .A2(new_n758), .A3(new_n762), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT105), .B1(new_n771), .B2(new_n772), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n700), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n657), .A2(new_n727), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n708), .A2(new_n863), .A3(new_n719), .A4(new_n755), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n730), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n860), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n690), .A2(new_n578), .A3(new_n696), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n763), .A2(new_n773), .B1(new_n867), .B2(new_n699), .ZN(new_n868));
  INV_X1    g682(.A(new_n865), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT52), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n846), .B(new_n857), .C1(new_n866), .C2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n861), .B1(new_n860), .B2(new_n865), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT52), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n854), .A2(new_n872), .A3(new_n855), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n856), .B(KEYINPUT116), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n846), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n876), .B1(KEYINPUT54), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n815), .A2(new_n648), .A3(new_n237), .A4(new_n754), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n736), .A2(new_n440), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n710), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT50), .Z(new_n891));
  INV_X1    g705(.A(new_n237), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n736), .A2(new_n776), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n815), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n894), .A2(new_n690), .A3(new_n754), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT118), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n720), .A2(new_n648), .A3(new_n893), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT119), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n323), .A3(new_n667), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n830), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n327), .B1(new_n837), .B2(KEYINPUT117), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(KEYINPUT117), .B2(new_n837), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n776), .B(new_n886), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n885), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n902), .A2(new_n904), .ZN(new_n907));
  INV_X1    g721(.A(new_n886), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n907), .A2(new_n440), .A3(new_n709), .A4(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n897), .A3(KEYINPUT51), .A4(new_n900), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n899), .A2(new_n668), .ZN(new_n911));
  INV_X1    g725(.A(G952), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n912), .B(G953), .C1(new_n908), .C2(new_n747), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n894), .A2(new_n648), .A3(new_n786), .ZN(new_n916));
  NOR2_X1   g730(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n906), .A2(new_n910), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n884), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(G952), .A2(G953), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n841), .B1(new_n921), .B2(new_n922), .ZN(G75));
  NAND2_X1  g737(.A1(new_n912), .A2(G953), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT123), .Z(new_n925));
  NAND4_X1  g739(.A1(new_n883), .A2(KEYINPUT122), .A3(G210), .A4(G902), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n470), .A2(new_n472), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n477), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n187), .B1(new_n873), .B2(new_n882), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT122), .B1(new_n932), .B2(G210), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n925), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT56), .B1(new_n932), .B2(G210), .ZN(new_n935));
  INV_X1    g749(.A(new_n929), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT121), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n932), .A2(G210), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n938), .B(new_n929), .C1(new_n939), .C2(KEYINPUT56), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n934), .B1(new_n937), .B2(new_n940), .ZN(G51));
  INV_X1    g755(.A(new_n925), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n883), .B(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n799), .B(KEYINPUT57), .Z(new_n945));
  OAI21_X1  g759(.A(new_n732), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n932), .A2(new_n797), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(G54));
  AND2_X1   g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  AND4_X1   g763(.A1(G902), .A2(new_n883), .A3(new_n308), .A4(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n308), .B1(new_n932), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n925), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(KEYINPUT124), .B(new_n925), .C1(new_n950), .C2(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(G60));
  AND2_X1   g770(.A1(new_n664), .A2(new_n665), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n658), .B(KEYINPUT59), .Z(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n884), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n925), .B1(new_n944), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(G63));
  XNOR2_X1  g777(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n227), .A2(new_n187), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n883), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n625), .ZN(new_n968));
  INV_X1    g782(.A(new_n682), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n883), .A2(new_n969), .A3(new_n966), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n925), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n968), .A2(KEYINPUT61), .A3(new_n925), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(G66));
  INV_X1    g789(.A(new_n239), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n236), .B1(new_n976), .B2(G224), .ZN(new_n977));
  INV_X1    g791(.A(new_n857), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n236), .ZN(new_n979));
  INV_X1    g793(.A(G898), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n927), .B1(new_n980), .B2(G953), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n979), .B(new_n981), .ZN(G69));
  INV_X1    g796(.A(G227), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n983), .B2(new_n697), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n868), .A2(new_n730), .ZN(new_n985));
  INV_X1    g799(.A(new_n791), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n788), .A2(new_n986), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n985), .B(new_n987), .C1(new_n830), .C2(new_n831), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n808), .A2(new_n648), .A3(new_n755), .A4(new_n786), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n823), .A2(new_n988), .A3(new_n236), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n537), .B1(KEYINPUT30), .B2(new_n530), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(new_n298), .Z(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(G900), .B2(G953), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n992), .ZN(new_n995));
  OR3_X1    g809(.A1(new_n985), .A2(KEYINPUT62), .A3(new_n721), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT62), .B1(new_n985), .B2(new_n721), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n578), .A2(new_n648), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n850), .A2(new_n668), .ZN(new_n999));
  NOR4_X1   g813(.A1(new_n998), .A2(new_n999), .A3(new_n704), .A4(new_n776), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n830), .B2(new_n831), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n823), .A2(new_n996), .A3(new_n997), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n995), .B1(new_n1002), .B2(new_n236), .ZN(new_n1003));
  OAI211_X1 g817(.A(KEYINPUT126), .B(new_n984), .C1(new_n994), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1002), .A2(new_n236), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n992), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n990), .A2(new_n993), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1004), .A2(new_n1010), .ZN(G72));
  XNOR2_X1  g825(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n651), .A2(new_n187), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1012), .B(new_n1013), .Z(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(new_n1002), .B2(new_n978), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n717), .ZN(new_n1016));
  AND4_X1   g830(.A1(new_n823), .A2(new_n988), .A3(new_n857), .A4(new_n989), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1014), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n525), .B(new_n554), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n541), .B1(new_n554), .B2(new_n504), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1014), .B(new_n1020), .C1(new_n874), .C2(new_n875), .ZN(new_n1021));
  AND4_X1   g835(.A1(new_n925), .A2(new_n1016), .A3(new_n1019), .A4(new_n1021), .ZN(G57));
endmodule


