//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n461), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n465), .B1(new_n470), .B2(KEYINPUT69), .ZN(new_n471));
  OR3_X1    g046(.A1(new_n466), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(G137), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(new_n464), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n469), .B1(new_n475), .B2(new_n461), .ZN(G160));
  NAND3_X1  g051(.A1(new_n471), .A2(G2105), .A3(new_n472), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(new_n461), .A3(new_n472), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n479), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n471), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n471), .A2(new_n461), .A3(new_n472), .A4(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n461), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(G62), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT72), .A4(G62), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n502), .B(new_n504), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT71), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(G88), .A3(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n501), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n511), .A2(new_n520), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  OAI211_X1 g101(.A(G51), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(G76), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n502), .A2(new_n504), .ZN(new_n533));
  INV_X1    g108(.A(G63), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n533), .A2(new_n534), .B1(new_n528), .B2(new_n529), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n532), .B1(G651), .B2(new_n535), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT73), .B(G89), .Z(new_n537));
  NAND3_X1  g112(.A1(new_n516), .A2(new_n519), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G168));
  NAND3_X1  g114(.A1(new_n502), .A2(new_n504), .A3(G64), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G651), .B1(G52), .B2(new_n523), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n516), .A2(G90), .A3(new_n519), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n530), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n516), .A2(G81), .A3(new_n519), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT74), .B(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n523), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n549), .A2(KEYINPUT75), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(KEYINPUT75), .B1(new_n549), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT76), .Z(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND3_X1  g137(.A1(new_n516), .A2(G91), .A3(new_n519), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n518), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n530), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT77), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n567), .A2(new_n568), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n533), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n572), .A2(new_n573), .A3(new_n563), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n543), .A2(new_n544), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G301));
  NAND2_X1  g159(.A1(new_n536), .A2(new_n538), .ZN(G286));
  AND2_X1   g160(.A1(new_n516), .A2(new_n519), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT79), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n523), .A2(G49), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n533), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G48), .B2(new_n523), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n516), .A2(G86), .A3(new_n519), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n533), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G47), .B2(new_n523), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n516), .A2(G85), .A3(new_n519), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n516), .A2(new_n519), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n516), .A2(new_n519), .A3(KEYINPUT10), .A4(G92), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n517), .A2(G66), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT80), .Z(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n523), .A2(G54), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n611), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n605), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n605), .B1(new_n618), .B2(G868), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n579), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n579), .B2(G868), .ZN(G280));
  NOR2_X1   g198(.A1(new_n617), .A2(G559), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G860), .B2(new_n618), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT81), .Z(G148));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n554), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n624), .B2(new_n627), .ZN(G323));
  XOR2_X1   g204(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n630));
  XNOR2_X1  g205(.A(G323), .B(new_n630), .ZN(G282));
  NAND2_X1  g206(.A1(new_n478), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT83), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n656), .A2(KEYINPUT86), .A3(new_n658), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n651), .B(new_n654), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n661), .B1(new_n662), .B2(new_n657), .ZN(new_n663));
  OAI211_X1 g238(.A(G14), .B(new_n659), .C1(new_n660), .C2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(KEYINPUT17), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n675), .A3(new_n669), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n670), .B(KEYINPUT87), .Z(new_n677));
  OAI211_X1 g252(.A(new_n672), .B(new_n676), .C1(new_n674), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n683), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n687), .A2(KEYINPUT20), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n683), .A3(new_n686), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n690), .B(new_n692), .C1(KEYINPUT20), .C2(new_n687), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1986), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1991), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G35), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G162), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT29), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G2090), .ZN(new_n704));
  NOR2_X1   g279(.A1(G29), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n478), .A2(G129), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n481), .A2(G141), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n706), .A2(new_n707), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n705), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(new_n700), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G160), .B2(new_n700), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G2084), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT94), .B1(G29), .B2(G33), .ZN(new_n723));
  OR3_X1    g298(.A1(KEYINPUT94), .A2(G29), .A3(G33), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n471), .A2(G139), .A3(new_n461), .A4(new_n472), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n465), .A2(new_n467), .A3(G127), .ZN(new_n726));
  INV_X1    g301(.A(G115), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n464), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G2105), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n725), .B(new_n729), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n723), .B(new_n724), .C1(new_n736), .C2(new_n700), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT96), .B(G2072), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G168), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G21), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT99), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT30), .B2(new_n746), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n636), .B2(new_n700), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n745), .B(new_n749), .C1(new_n741), .C2(new_n742), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n722), .A2(new_n739), .A3(new_n744), .A4(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G5), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G171), .B2(new_n752), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT100), .B(G1961), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n754), .B(new_n755), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(KEYINPUT23), .A3(G20), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n758));
  INV_X1    g333(.A(G20), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G16), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n760), .C1(new_n579), .C2(new_n752), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1956), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n751), .A2(new_n756), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n703), .A2(G2090), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT101), .ZN(new_n765));
  OAI21_X1  g340(.A(KEYINPUT91), .B1(G4), .B2(G16), .ZN(new_n766));
  OR3_X1    g341(.A1(KEYINPUT91), .A2(G4), .A3(G16), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(new_n617), .C2(new_n752), .ZN(new_n768));
  INV_X1    g343(.A(G1348), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n752), .A2(G19), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n555), .B2(new_n752), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1341), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n700), .A2(G26), .ZN(new_n774));
  INV_X1    g349(.A(G140), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n480), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT92), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT93), .B1(G104), .B2(G2105), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(KEYINPUT93), .A2(G104), .A3(G2105), .ZN(new_n781));
  OAI221_X1 g356(.A(G2104), .B1(G116), .B2(new_n461), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n478), .A2(G128), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n778), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n774), .B1(new_n784), .B2(new_n700), .ZN(new_n785));
  MUX2_X1   g360(.A(new_n774), .B(new_n785), .S(KEYINPUT28), .Z(new_n786));
  AOI211_X1 g361(.A(new_n770), .B(new_n773), .C1(new_n786), .C2(G2067), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(G2067), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n700), .A2(G27), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G164), .B2(new_n700), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n763), .A2(new_n765), .A3(new_n787), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n752), .A2(G23), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n591), .B2(new_n752), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT33), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1976), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n752), .A2(G6), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n596), .A2(new_n597), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n752), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT90), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT32), .B(G1981), .Z(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n752), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n752), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(G1971), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n804), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n798), .B(new_n809), .C1(G1971), .C2(new_n807), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT89), .B(KEYINPUT34), .Z(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n752), .A2(G24), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G290), .B2(G16), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G1986), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT88), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n478), .A2(new_n817), .A3(G119), .ZN(new_n818));
  INV_X1    g393(.A(G119), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT88), .B1(new_n477), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(G95), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n823));
  INV_X1    g398(.A(G131), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n480), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n821), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  MUX2_X1   g402(.A(G25), .B(new_n827), .S(G29), .Z(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G1991), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(G1986), .B2(new_n815), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n829), .B2(new_n828), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n810), .B2(new_n811), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n812), .A2(new_n816), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT36), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(KEYINPUT36), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n704), .B(new_n794), .C1(new_n834), .C2(new_n835), .ZN(G311));
  AOI21_X1  g411(.A(new_n794), .B1(new_n834), .B2(new_n835), .ZN(new_n837));
  INV_X1    g412(.A(new_n704), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(G150));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n533), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G651), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n523), .A2(G55), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n843), .B(new_n844), .C1(new_n607), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n618), .A2(G559), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT39), .Z(new_n850));
  INV_X1    g425(.A(new_n846), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n554), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n548), .B(new_n846), .C1(new_n552), .C2(new_n553), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n850), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n848), .B1(new_n857), .B2(G860), .ZN(G145));
  NAND3_X1  g433(.A1(new_n778), .A2(new_n782), .A3(new_n783), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n734), .A2(new_n735), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n729), .A2(new_n725), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n494), .A2(new_n487), .A3(new_n497), .A4(new_n489), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n736), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n863), .A2(new_n865), .A3(new_n712), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n712), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n859), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n713), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n863), .A2(new_n865), .A3(new_n712), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n784), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n639), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n827), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n478), .A2(G130), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n481), .A2(G142), .ZN(new_n876));
  OR2_X1    g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n825), .B1(new_n818), .B2(new_n820), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n639), .A3(new_n823), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n874), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n880), .B1(new_n874), .B2(new_n882), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n868), .B(new_n872), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n868), .A2(new_n872), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT105), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n888), .B2(KEYINPUT103), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n885), .A2(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n887), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT104), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n889), .A2(new_n890), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n636), .B(G160), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G162), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n885), .A3(new_n891), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g478(.A1(new_n846), .A2(new_n627), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n617), .A2(new_n579), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n609), .A2(new_n610), .B1(G54), .B2(new_n523), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n907), .A2(new_n615), .B1(new_n571), .B2(new_n578), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n905), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n617), .A2(new_n579), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n907), .A2(new_n571), .A3(new_n578), .A4(new_n615), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT41), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n854), .B(new_n624), .ZN(new_n916));
  MUX2_X1   g491(.A(new_n913), .B(new_n915), .S(new_n916), .Z(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n602), .A2(new_n918), .A3(new_n603), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n602), .B2(new_n603), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(G303), .A2(new_n800), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n520), .A2(new_n524), .ZN(new_n923));
  AOI21_X1  g498(.A(G305), .B1(new_n923), .B2(new_n511), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n516), .A2(G85), .A3(new_n519), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n523), .A2(G47), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n530), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT106), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n602), .A2(new_n918), .A3(new_n603), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(G303), .A2(new_n800), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n923), .A2(new_n511), .A3(G305), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n925), .A2(new_n591), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n591), .B1(new_n925), .B2(new_n935), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT42), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n936), .B2(new_n937), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n932), .B1(new_n934), .B2(new_n933), .ZN(new_n942));
  OAI21_X1  g517(.A(G288), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n925), .A2(new_n591), .A3(new_n935), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(KEYINPUT107), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n938), .B1(new_n946), .B2(KEYINPUT42), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n917), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n904), .B1(new_n948), .B2(new_n627), .ZN(G295));
  OAI21_X1  g524(.A(new_n904), .B1(new_n948), .B2(new_n627), .ZN(G331));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n543), .A2(new_n544), .A3(new_n582), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n582), .B1(new_n543), .B2(new_n544), .ZN(new_n953));
  OAI21_X1  g528(.A(G168), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(G171), .A2(G286), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n956), .A2(new_n852), .A3(new_n853), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n853), .B2(new_n852), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n915), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n545), .B1(new_n536), .B2(new_n538), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(G301), .B2(G168), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n549), .A2(new_n551), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT75), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n549), .A2(KEYINPUT75), .A3(new_n551), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n846), .B1(new_n966), .B2(new_n548), .ZN(new_n967));
  INV_X1    g542(.A(new_n853), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n956), .A2(new_n852), .A3(new_n853), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n909), .A2(new_n969), .A3(new_n912), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n959), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G37), .B1(new_n946), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT107), .B1(new_n943), .B2(new_n944), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n914), .B1(new_n969), .B2(new_n970), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n957), .A2(new_n958), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n913), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT108), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n940), .A2(new_n959), .A3(new_n945), .A4(new_n971), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n951), .B(new_n973), .C1(new_n980), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT109), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n973), .A2(new_n981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n976), .A2(KEYINPUT108), .A3(new_n979), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n981), .A2(new_n982), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n951), .A4(new_n973), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n985), .A2(new_n987), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(KEYINPUT43), .A3(new_n973), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n986), .A2(new_n951), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  MUX2_X1   g571(.A(new_n993), .B(new_n996), .S(KEYINPUT44), .Z(G397));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n862), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n475), .A2(new_n461), .ZN(new_n1002));
  INV_X1    g577(.A(new_n469), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(G40), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n492), .B2(new_n498), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1007));
  INV_X1    g582(.A(G1971), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1002), .A2(G40), .A3(new_n1003), .ZN(new_n1010));
  INV_X1    g585(.A(new_n999), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1010), .B(KEYINPUT115), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n862), .B2(new_n998), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1004), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n499), .A2(new_n998), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1014), .B(new_n1017), .C1(new_n1018), .C2(KEYINPUT50), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1009), .B1(new_n1019), .B2(G2090), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G8), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT55), .Z(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1004), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1006), .B2(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1029), .A2(G2090), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1026), .B1(new_n1030), .B2(new_n1009), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1023), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G8), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(G1981), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n800), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G305), .A2(G1981), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1038), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  OAI221_X1 g618(.A(new_n1035), .B1(KEYINPUT49), .B2(new_n1039), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n591), .A2(G1976), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1033), .A2(new_n1045), .A3(G8), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(KEYINPUT112), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  NAND3_X1  g624(.A1(G288), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1047), .A2(KEYINPUT112), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1033), .A2(new_n1045), .A3(G8), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n999), .A2(new_n1000), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1010), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n742), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1027), .B(new_n1060), .C1(new_n1006), .C2(new_n1028), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1026), .B(G286), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1025), .A2(new_n1032), .A3(new_n1055), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT116), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT63), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1054), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n1025), .A4(new_n1062), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(KEYINPUT63), .A3(new_n1062), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1031), .A2(new_n1023), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT117), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1032), .A2(new_n1055), .A3(new_n1062), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1071), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(KEYINPUT63), .A4(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1069), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1019), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1007), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n572), .A2(KEYINPUT118), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1084), .A2(KEYINPUT57), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n572), .A2(new_n563), .A3(new_n577), .ZN(new_n1086));
  XOR2_X1   g661(.A(new_n1085), .B(new_n1086), .Z(new_n1087));
  AND3_X1   g662(.A1(new_n1080), .A2(new_n1083), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1078), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n617), .A2(KEYINPUT121), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1029), .A2(new_n769), .ZN(new_n1093));
  INV_X1    g668(.A(G2067), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1010), .A2(new_n1094), .A3(new_n1011), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1092), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n617), .A2(KEYINPUT121), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1093), .A2(KEYINPUT60), .A3(new_n1095), .A4(new_n1091), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1098), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1019), .A2(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1087), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT61), .ZN(new_n1105));
  INV_X1    g680(.A(G1996), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1005), .B(new_n1106), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT58), .B(G1341), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1033), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n554), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT59), .Z(new_n1111));
  NAND4_X1  g686(.A1(new_n1090), .A2(new_n1102), .A3(new_n1105), .A4(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1103), .A2(KEYINPUT119), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1087), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1103), .A2(KEYINPUT119), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1104), .A2(new_n618), .A3(new_n1096), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1066), .A2(new_n1025), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1007), .B2(G2078), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1010), .B(KEYINPUT123), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1001), .B1(new_n1124), .B2(new_n791), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1122), .A2(new_n1057), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1961), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1029), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1121), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  INV_X1    g705(.A(G301), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1121), .B(new_n1128), .C1(new_n1058), .C2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT54), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1131), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1136), .B(new_n1137), .C1(new_n1131), .C2(new_n1129), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1119), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1059), .A2(G168), .A3(new_n1061), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT51), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(G8), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1146), .A2(G8), .A3(G286), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1144), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1140), .A2(G8), .A3(new_n1142), .A4(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1118), .A2(new_n1139), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1044), .A2(new_n1049), .A3(new_n591), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1034), .B1(new_n1152), .B2(new_n1037), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1032), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n1055), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1150), .A2(KEYINPUT62), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1119), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1136), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1145), .A2(new_n1159), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1077), .A2(new_n1151), .A3(new_n1155), .A4(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1057), .A2(new_n1004), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1164), .A2(new_n1106), .A3(new_n713), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(KEYINPUT110), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1165), .A2(KEYINPUT110), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n859), .B(new_n1094), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(G1996), .B2(new_n712), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1166), .B(new_n1167), .C1(new_n1163), .C2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n827), .B(new_n829), .Z(new_n1171));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n1164), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(G290), .B(G1986), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1163), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1162), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1163), .A2(new_n1106), .ZN(new_n1176));
  NAND2_X1  g751(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1176), .B(new_n1177), .Z(new_n1178));
  AND2_X1   g753(.A1(new_n1168), .A2(new_n713), .ZN(new_n1179));
  OAI221_X1 g754(.A(new_n1178), .B1(KEYINPUT125), .B2(KEYINPUT46), .C1(new_n1179), .C2(new_n1164), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT47), .Z(new_n1181));
  NOR3_X1   g756(.A1(new_n1164), .A2(G1986), .A3(G290), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT48), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1172), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n827), .A2(new_n829), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1170), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n784), .A2(new_n1094), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1164), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1181), .A2(new_n1184), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1175), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g765(.A1(G229), .A2(new_n459), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n664), .A2(new_n680), .ZN(new_n1193));
  AOI21_X1  g767(.A(new_n1193), .B1(new_n898), .B2(new_n901), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n993), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n993), .A2(new_n1194), .A3(new_n1197), .A4(new_n1192), .ZN(new_n1198));
  AND2_X1   g772(.A1(new_n1196), .A2(new_n1198), .ZN(G308));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(G225));
endmodule


