

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739;

  AND2_X1 U366 ( .A1(n604), .A2(n577), .ZN(n571) );
  XNOR2_X1 U367 ( .A(n571), .B(KEYINPUT40), .ZN(n737) );
  INV_X2 U368 ( .A(G143), .ZN(n416) );
  XNOR2_X2 U369 ( .A(n495), .B(KEYINPUT19), .ZN(n574) );
  XNOR2_X2 U370 ( .A(n371), .B(KEYINPUT39), .ZN(n604) );
  XNOR2_X2 U371 ( .A(n463), .B(KEYINPUT10), .ZN(n719) );
  XNOR2_X2 U372 ( .A(n521), .B(G472), .ZN(n559) );
  NOR2_X2 U373 ( .A1(n363), .A2(n588), .ZN(n532) );
  XNOR2_X1 U374 ( .A(n478), .B(n383), .ZN(n372) );
  NAND2_X1 U375 ( .A1(n417), .A2(n351), .ZN(n612) );
  NOR2_X1 U376 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U377 ( .A(n523), .B(KEYINPUT105), .ZN(n734) );
  NOR2_X1 U378 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X1 U379 ( .A(n376), .B(n375), .ZN(n593) );
  NOR2_X1 U380 ( .A1(n570), .A2(n569), .ZN(n591) );
  XNOR2_X1 U381 ( .A(n560), .B(KEYINPUT1), .ZN(n621) );
  XNOR2_X1 U382 ( .A(n404), .B(KEYINPUT102), .ZN(n577) );
  XNOR2_X1 U383 ( .A(n461), .B(n462), .ZN(n537) );
  XNOR2_X1 U384 ( .A(n372), .B(n479), .ZN(n382) );
  XNOR2_X1 U385 ( .A(n366), .B(G104), .ZN(n485) );
  XOR2_X1 U386 ( .A(G137), .B(KEYINPUT69), .Z(n508) );
  XNOR2_X2 U387 ( .A(n400), .B(n530), .ZN(n645) );
  NOR2_X1 U388 ( .A1(G902), .A2(G237), .ZN(n489) );
  INV_X1 U389 ( .A(KEYINPUT6), .ZN(n378) );
  AND2_X1 U390 ( .A1(n608), .A2(n607), .ZN(n724) );
  XOR2_X1 U391 ( .A(KEYINPUT76), .B(G110), .Z(n483) );
  XNOR2_X1 U392 ( .A(n482), .B(n382), .ZN(n423) );
  NOR2_X1 U393 ( .A1(G953), .A2(G237), .ZN(n467) );
  XOR2_X1 U394 ( .A(KEYINPUT68), .B(G131), .Z(n464) );
  NOR2_X1 U395 ( .A1(n734), .A2(n733), .ZN(n533) );
  INV_X1 U396 ( .A(G101), .ZN(n427) );
  NAND2_X1 U397 ( .A1(n711), .A2(n724), .ZN(n657) );
  NOR2_X1 U398 ( .A1(n537), .A2(n529), .ZN(n640) );
  XNOR2_X1 U399 ( .A(n445), .B(G469), .ZN(n446) );
  NOR2_X1 U400 ( .A1(G902), .A2(n694), .ZN(n447) );
  INV_X1 U401 ( .A(G953), .ZN(n725) );
  XNOR2_X1 U402 ( .A(G116), .B(G107), .ZN(n488) );
  INV_X1 U403 ( .A(G122), .ZN(n366) );
  INV_X1 U404 ( .A(KEYINPUT16), .ZN(n365) );
  XNOR2_X1 U405 ( .A(n414), .B(n413), .ZN(n702) );
  XNOR2_X1 U406 ( .A(n456), .B(n345), .ZN(n413) );
  XNOR2_X1 U407 ( .A(n460), .B(n415), .ZN(n414) );
  XNOR2_X1 U408 ( .A(n477), .B(G146), .ZN(n439) );
  XNOR2_X1 U409 ( .A(n438), .B(n440), .ZN(n402) );
  INV_X1 U410 ( .A(G140), .ZN(n440) );
  INV_X1 U411 ( .A(G104), .ZN(n436) );
  XNOR2_X1 U412 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U413 ( .A(KEYINPUT91), .ZN(n490) );
  NAND2_X1 U414 ( .A1(n591), .A2(n638), .ZN(n371) );
  AND2_X1 U415 ( .A1(n557), .A2(n526), .ZN(n425) );
  XNOR2_X1 U416 ( .A(n544), .B(KEYINPUT81), .ZN(n525) );
  NOR2_X1 U417 ( .A1(n537), .A2(n536), .ZN(n404) );
  NAND2_X1 U418 ( .A1(n704), .A2(n350), .ZN(n395) );
  NOR2_X1 U419 ( .A1(n387), .A2(n354), .ZN(n386) );
  INV_X1 U420 ( .A(n392), .ZN(n387) );
  NAND2_X1 U421 ( .A1(n390), .A2(n354), .ZN(n389) );
  NAND2_X1 U422 ( .A1(n395), .A2(n392), .ZN(n390) );
  NOR2_X1 U423 ( .A1(n704), .A2(n398), .ZN(n397) );
  INV_X1 U424 ( .A(n613), .ZN(n398) );
  BUF_X1 U425 ( .A(n725), .Z(n374) );
  NAND2_X1 U426 ( .A1(n704), .A2(n349), .ZN(n408) );
  NOR2_X1 U427 ( .A1(n407), .A2(n708), .ZN(n406) );
  NOR2_X1 U428 ( .A1(n348), .A2(G475), .ZN(n407) );
  NOR2_X1 U429 ( .A1(n634), .A2(n678), .ZN(n586) );
  INV_X1 U430 ( .A(KEYINPUT83), .ZN(n375) );
  XNOR2_X1 U431 ( .A(G116), .B(G137), .ZN(n429) );
  NOR2_X1 U432 ( .A1(n605), .A2(n577), .ZN(n634) );
  INV_X1 U433 ( .A(KEYINPUT70), .ZN(n595) );
  INV_X1 U434 ( .A(KEYINPUT44), .ZN(n534) );
  XOR2_X1 U435 ( .A(G125), .B(G146), .Z(n481) );
  XOR2_X1 U436 ( .A(KEYINPUT8), .B(n455), .Z(n509) );
  NAND2_X1 U437 ( .A1(G234), .A2(n725), .ZN(n455) );
  XOR2_X1 U438 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n451) );
  XNOR2_X1 U439 ( .A(G134), .B(KEYINPUT9), .ZN(n450) );
  XNOR2_X1 U440 ( .A(n453), .B(n454), .ZN(n415) );
  XOR2_X1 U441 ( .A(KEYINPUT96), .B(KEYINPUT99), .Z(n454) );
  INV_X1 U442 ( .A(KEYINPUT100), .ZN(n458) );
  XNOR2_X1 U443 ( .A(G143), .B(G113), .ZN(n465) );
  XOR2_X1 U444 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n469) );
  INV_X1 U445 ( .A(KEYINPUT89), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n481), .B(n381), .ZN(n482) );
  XNOR2_X1 U447 ( .A(KEYINPUT17), .B(KEYINPUT90), .ZN(n381) );
  XNOR2_X1 U448 ( .A(KEYINPUT38), .B(n589), .ZN(n638) );
  NOR2_X1 U449 ( .A1(n566), .A2(n567), .ZN(n568) );
  AND2_X1 U450 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U451 ( .A1(n613), .A2(n396), .ZN(n394) );
  XNOR2_X1 U452 ( .A(G128), .B(G119), .ZN(n505) );
  AND2_X1 U453 ( .A1(n724), .A2(n610), .ZN(n418) );
  NOR2_X1 U454 ( .A1(n544), .A2(n411), .ZN(n410) );
  NAND2_X1 U455 ( .A1(n412), .A2(n637), .ZN(n411) );
  INV_X1 U456 ( .A(n579), .ZN(n412) );
  XNOR2_X1 U457 ( .A(n563), .B(KEYINPUT41), .ZN(n632) );
  XNOR2_X1 U458 ( .A(n621), .B(n368), .ZN(n582) );
  INV_X1 U459 ( .A(KEYINPUT86), .ZN(n368) );
  XNOR2_X1 U460 ( .A(n476), .B(n373), .ZN(n536) );
  XNOR2_X1 U461 ( .A(n475), .B(G475), .ZN(n373) );
  NOR2_X1 U462 ( .A1(n559), .A2(n579), .ZN(n377) );
  INV_X1 U463 ( .A(KEYINPUT104), .ZN(n420) );
  NAND2_X1 U464 ( .A1(n380), .A2(n379), .ZN(n545) );
  INV_X1 U465 ( .A(n621), .ZN(n379) );
  XNOR2_X1 U466 ( .A(n487), .B(n421), .ZN(n714) );
  XNOR2_X1 U467 ( .A(n486), .B(n488), .ZN(n421) );
  XNOR2_X1 U468 ( .A(n485), .B(n365), .ZN(n486) );
  XNOR2_X1 U469 ( .A(n444), .B(n443), .ZN(n694) );
  XNOR2_X1 U470 ( .A(n439), .B(n402), .ZN(n444) );
  INV_X1 U471 ( .A(KEYINPUT116), .ZN(n369) );
  XNOR2_X1 U472 ( .A(n399), .B(KEYINPUT34), .ZN(n363) );
  XNOR2_X1 U473 ( .A(n528), .B(n364), .ZN(n733) );
  INV_X1 U474 ( .A(KEYINPUT64), .ZN(n364) );
  XNOR2_X1 U475 ( .A(n577), .B(n403), .ZN(n679) );
  INV_X1 U476 ( .A(KEYINPUT106), .ZN(n403) );
  OR2_X1 U477 ( .A1(n575), .A2(n574), .ZN(n678) );
  INV_X1 U478 ( .A(n679), .ZN(n681) );
  OR2_X1 U479 ( .A1(n384), .A2(n397), .ZN(n385) );
  AND2_X1 U480 ( .A1(n391), .A2(n389), .ZN(n388) );
  XNOR2_X1 U481 ( .A(n358), .B(n357), .ZN(G63) );
  INV_X1 U482 ( .A(KEYINPUT124), .ZN(n357) );
  NOR2_X1 U483 ( .A1(n409), .A2(n405), .ZN(n701) );
  NOR2_X1 U484 ( .A1(n704), .A2(n348), .ZN(n409) );
  NAND2_X1 U485 ( .A1(n408), .A2(n406), .ZN(n405) );
  XNOR2_X1 U486 ( .A(n356), .B(n355), .ZN(G51) );
  INV_X1 U487 ( .A(KEYINPUT56), .ZN(n355) );
  XOR2_X1 U488 ( .A(n451), .B(n450), .Z(n345) );
  XOR2_X1 U489 ( .A(G113), .B(G119), .Z(n346) );
  XNOR2_X1 U490 ( .A(n559), .B(n378), .ZN(n544) );
  XNOR2_X1 U491 ( .A(n504), .B(KEYINPUT22), .ZN(n524) );
  OR2_X1 U492 ( .A1(n652), .A2(n651), .ZN(n347) );
  XOR2_X1 U493 ( .A(n700), .B(n699), .Z(n348) );
  AND2_X1 U494 ( .A1(n348), .A2(G475), .ZN(n349) );
  NOR2_X1 U495 ( .A1(n613), .A2(n396), .ZN(n350) );
  XOR2_X1 U496 ( .A(n611), .B(KEYINPUT65), .Z(n351) );
  XNOR2_X1 U497 ( .A(n616), .B(n615), .ZN(n352) );
  XNOR2_X1 U498 ( .A(n702), .B(KEYINPUT123), .ZN(n353) );
  NOR2_X1 U499 ( .A1(G952), .A2(n374), .ZN(n708) );
  INV_X1 U500 ( .A(n708), .ZN(n393) );
  XOR2_X1 U501 ( .A(KEYINPUT63), .B(KEYINPUT109), .Z(n354) );
  XNOR2_X1 U502 ( .A(n532), .B(n531), .ZN(n736) );
  NAND2_X1 U503 ( .A1(n359), .A2(n393), .ZN(n356) );
  NAND2_X1 U504 ( .A1(n360), .A2(n393), .ZN(n358) );
  XNOR2_X1 U505 ( .A(n617), .B(n352), .ZN(n359) );
  NAND2_X1 U506 ( .A1(n362), .A2(KEYINPUT2), .ZN(n426) );
  XNOR2_X1 U507 ( .A(n703), .B(n353), .ZN(n360) );
  OR2_X2 U508 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U509 ( .A1(n704), .A2(G210), .ZN(n617) );
  NAND2_X1 U510 ( .A1(n704), .A2(G478), .ZN(n703) );
  INV_X1 U511 ( .A(n657), .ZN(n362) );
  NAND2_X1 U512 ( .A1(n622), .A2(n560), .ZN(n566) );
  XNOR2_X1 U513 ( .A(n439), .B(n361), .ZN(n435) );
  INV_X1 U514 ( .A(n441), .ZN(n361) );
  XNOR2_X1 U515 ( .A(n512), .B(n424), .ZN(n513) );
  INV_X1 U516 ( .A(n559), .ZN(n628) );
  XNOR2_X1 U517 ( .A(n545), .B(n420), .ZN(n419) );
  NAND2_X1 U518 ( .A1(n541), .A2(n503), .ZN(n504) );
  XNOR2_X2 U519 ( .A(n502), .B(n501), .ZN(n541) );
  NAND2_X1 U520 ( .A1(n592), .A2(n677), .ZN(n376) );
  AND2_X1 U521 ( .A1(n632), .A2(n367), .ZN(n564) );
  INV_X1 U522 ( .A(n575), .ZN(n367) );
  XNOR2_X1 U523 ( .A(n370), .B(n369), .ZN(n664) );
  NAND2_X1 U524 ( .A1(n662), .A2(n663), .ZN(n370) );
  XNOR2_X1 U525 ( .A(n377), .B(KEYINPUT28), .ZN(n561) );
  XNOR2_X1 U526 ( .A(n527), .B(KEYINPUT32), .ZN(n528) );
  INV_X1 U527 ( .A(n524), .ZN(n380) );
  NAND2_X1 U528 ( .A1(n681), .A2(n410), .ZN(n600) );
  NOR2_X2 U529 ( .A1(n614), .A2(n610), .ZN(n493) );
  NAND2_X1 U530 ( .A1(n380), .A2(n425), .ZN(n527) );
  NOR2_X1 U531 ( .A1(n600), .A2(n589), .ZN(n581) );
  NAND2_X1 U532 ( .A1(n395), .A2(n386), .ZN(n384) );
  NAND2_X1 U533 ( .A1(n388), .A2(n385), .ZN(G57) );
  NAND2_X1 U534 ( .A1(n397), .A2(n354), .ZN(n391) );
  INV_X1 U535 ( .A(G472), .ZN(n396) );
  NAND2_X1 U536 ( .A1(n645), .A2(n541), .ZN(n399) );
  NAND2_X1 U537 ( .A1(n401), .A2(n578), .ZN(n400) );
  INV_X1 U538 ( .A(n540), .ZN(n401) );
  XNOR2_X2 U539 ( .A(n723), .B(n427), .ZN(n477) );
  XNOR2_X2 U540 ( .A(n493), .B(n492), .ZN(n603) );
  AND2_X4 U541 ( .A1(n426), .A2(n612), .ZN(n704) );
  XNOR2_X2 U542 ( .A(n452), .B(KEYINPUT4), .ZN(n723) );
  XNOR2_X2 U543 ( .A(n416), .B(G128), .ZN(n452) );
  NAND2_X1 U544 ( .A1(n418), .A2(n711), .ZN(n417) );
  XNOR2_X2 U545 ( .A(n551), .B(KEYINPUT45), .ZN(n711) );
  NAND2_X1 U546 ( .A1(n419), .A2(n522), .ZN(n523) );
  XNOR2_X1 U547 ( .A(n422), .B(n714), .ZN(n614) );
  XNOR2_X1 U548 ( .A(n480), .B(n423), .ZN(n422) );
  XNOR2_X1 U549 ( .A(KEYINPUT23), .B(KEYINPUT84), .ZN(n424) );
  XNOR2_X1 U550 ( .A(n596), .B(n595), .ZN(n597) );
  INV_X1 U551 ( .A(n668), .ZN(n547) );
  XNOR2_X1 U552 ( .A(n437), .B(n436), .ZN(n438) );
  INV_X1 U553 ( .A(n689), .ZN(n606) );
  XNOR2_X1 U554 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U555 ( .A1(n690), .A2(n606), .ZN(n607) );
  XNOR2_X1 U556 ( .A(n721), .B(n442), .ZN(n443) );
  XNOR2_X1 U557 ( .A(KEYINPUT36), .B(KEYINPUT108), .ZN(n580) );
  XNOR2_X1 U558 ( .A(n514), .B(n513), .ZN(n706) );
  XNOR2_X1 U559 ( .A(n581), .B(n580), .ZN(n584) );
  XNOR2_X1 U560 ( .A(n667), .B(n666), .ZN(G75) );
  XOR2_X1 U561 ( .A(G134), .B(n464), .Z(n441) );
  XNOR2_X1 U562 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n428) );
  XNOR2_X1 U563 ( .A(n346), .B(n428), .ZN(n484) );
  XOR2_X1 U564 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n430) );
  XNOR2_X1 U565 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U566 ( .A(n484), .B(n431), .Z(n433) );
  NAND2_X1 U567 ( .A1(n467), .A2(G210), .ZN(n432) );
  XNOR2_X1 U568 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U569 ( .A(n435), .B(n434), .ZN(n520) );
  XNOR2_X1 U570 ( .A(n520), .B(KEYINPUT62), .ZN(n613) );
  XOR2_X1 U571 ( .A(G902), .B(KEYINPUT15), .Z(n610) );
  INV_X1 U572 ( .A(n610), .ZN(n609) );
  XNOR2_X1 U573 ( .A(G107), .B(n483), .ZN(n437) );
  XNOR2_X1 U574 ( .A(n508), .B(n441), .ZN(n721) );
  NAND2_X1 U575 ( .A1(G227), .A2(n374), .ZN(n442) );
  XNOR2_X1 U576 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n445) );
  XNOR2_X2 U577 ( .A(n447), .B(n446), .ZN(n560) );
  NAND2_X1 U578 ( .A1(n609), .A2(G234), .ZN(n448) );
  XNOR2_X1 U579 ( .A(n448), .B(KEYINPUT20), .ZN(n515) );
  NAND2_X1 U580 ( .A1(G221), .A2(n515), .ZN(n449) );
  XNOR2_X1 U581 ( .A(KEYINPUT21), .B(n449), .ZN(n556) );
  INV_X1 U582 ( .A(n556), .ZN(n618) );
  XNOR2_X1 U583 ( .A(KEYINPUT101), .B(G478), .ZN(n462) );
  XNOR2_X1 U584 ( .A(n452), .B(KEYINPUT97), .ZN(n453) );
  NAND2_X1 U585 ( .A1(G217), .A2(n509), .ZN(n456) );
  INV_X1 U586 ( .A(n488), .ZN(n457) );
  XNOR2_X1 U587 ( .A(n457), .B(G122), .ZN(n459) );
  NOR2_X1 U588 ( .A1(G902), .A2(n702), .ZN(n461) );
  XNOR2_X1 U589 ( .A(n481), .B(G140), .ZN(n463) );
  XNOR2_X1 U590 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U591 ( .A(n719), .B(n466), .ZN(n474) );
  NAND2_X1 U592 ( .A1(n467), .A2(G214), .ZN(n468) );
  XNOR2_X1 U593 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U594 ( .A(KEYINPUT94), .B(n470), .ZN(n472) );
  INV_X1 U595 ( .A(n485), .ZN(n471) );
  XNOR2_X1 U596 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U597 ( .A(n474), .B(n473), .ZN(n698) );
  NOR2_X1 U598 ( .A1(G902), .A2(n698), .ZN(n476) );
  XNOR2_X1 U599 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n475) );
  INV_X1 U600 ( .A(n536), .ZN(n529) );
  AND2_X1 U601 ( .A1(n618), .A2(n640), .ZN(n503) );
  INV_X1 U602 ( .A(n477), .ZN(n480) );
  XOR2_X1 U603 ( .A(KEYINPUT88), .B(KEYINPUT18), .Z(n479) );
  NAND2_X1 U604 ( .A1(G224), .A2(n725), .ZN(n478) );
  XNOR2_X1 U605 ( .A(n484), .B(n483), .ZN(n487) );
  XOR2_X1 U606 ( .A(KEYINPUT74), .B(n489), .Z(n494) );
  NAND2_X1 U607 ( .A1(n494), .A2(G210), .ZN(n491) );
  NAND2_X1 U608 ( .A1(n494), .A2(G214), .ZN(n637) );
  AND2_X2 U609 ( .A1(n603), .A2(n637), .ZN(n495) );
  NAND2_X1 U610 ( .A1(G234), .A2(G237), .ZN(n496) );
  XNOR2_X1 U611 ( .A(n496), .B(KEYINPUT14), .ZN(n497) );
  NAND2_X1 U612 ( .A1(n497), .A2(G952), .ZN(n652) );
  NOR2_X1 U613 ( .A1(G953), .A2(n652), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G902), .A2(n497), .ZN(n552) );
  OR2_X1 U615 ( .A1(n374), .A2(G898), .ZN(n716) );
  NOR2_X1 U616 ( .A1(n552), .A2(n716), .ZN(n498) );
  NOR2_X1 U617 ( .A1(n555), .A2(n498), .ZN(n499) );
  XNOR2_X1 U618 ( .A(n499), .B(KEYINPUT92), .ZN(n500) );
  NOR2_X2 U619 ( .A1(n574), .A2(n500), .ZN(n502) );
  XNOR2_X1 U620 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n501) );
  XOR2_X1 U621 ( .A(KEYINPUT24), .B(G110), .Z(n506) );
  XNOR2_X1 U622 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U623 ( .A(n507), .B(n719), .ZN(n514) );
  XOR2_X1 U624 ( .A(n508), .B(KEYINPUT79), .Z(n511) );
  NAND2_X1 U625 ( .A1(G221), .A2(n509), .ZN(n510) );
  XNOR2_X1 U626 ( .A(n511), .B(n510), .ZN(n512) );
  NOR2_X1 U627 ( .A1(n706), .A2(G902), .ZN(n519) );
  XOR2_X1 U628 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n517) );
  NAND2_X1 U629 ( .A1(n515), .A2(G217), .ZN(n516) );
  XNOR2_X1 U630 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X2 U631 ( .A(n519), .B(n518), .ZN(n557) );
  INV_X1 U632 ( .A(n557), .ZN(n619) );
  NOR2_X1 U633 ( .A1(n520), .A2(G902), .ZN(n521) );
  NOR2_X1 U634 ( .A1(n619), .A2(n628), .ZN(n522) );
  NOR2_X1 U635 ( .A1(n582), .A2(n525), .ZN(n526) );
  NAND2_X1 U636 ( .A1(n537), .A2(n529), .ZN(n588) );
  XOR2_X1 U637 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n530) );
  NOR2_X1 U638 ( .A1(n556), .A2(n557), .ZN(n622) );
  NAND2_X1 U639 ( .A1(n621), .A2(n622), .ZN(n540) );
  XNOR2_X1 U640 ( .A(KEYINPUT35), .B(KEYINPUT80), .ZN(n531) );
  NAND2_X1 U641 ( .A1(n533), .A2(n736), .ZN(n535) );
  XNOR2_X1 U642 ( .A(n535), .B(n534), .ZN(n550) );
  NAND2_X1 U643 ( .A1(n537), .A2(n536), .ZN(n674) );
  XNOR2_X1 U644 ( .A(KEYINPUT103), .B(n674), .ZN(n605) );
  NOR2_X1 U645 ( .A1(n566), .A2(n628), .ZN(n538) );
  NAND2_X1 U646 ( .A1(n541), .A2(n538), .ZN(n539) );
  XNOR2_X1 U647 ( .A(KEYINPUT93), .B(n539), .ZN(n670) );
  NOR2_X1 U648 ( .A1(n559), .A2(n540), .ZN(n630) );
  NAND2_X1 U649 ( .A1(n630), .A2(n541), .ZN(n542) );
  XNOR2_X1 U650 ( .A(n542), .B(KEYINPUT31), .ZN(n685) );
  NOR2_X1 U651 ( .A1(n670), .A2(n685), .ZN(n543) );
  NOR2_X1 U652 ( .A1(n634), .A2(n543), .ZN(n548) );
  INV_X1 U653 ( .A(n544), .ZN(n578) );
  NOR2_X1 U654 ( .A1(n578), .A2(n545), .ZN(n546) );
  NAND2_X1 U655 ( .A1(n619), .A2(n546), .ZN(n668) );
  NOR2_X1 U656 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U657 ( .A1(n550), .A2(n549), .ZN(n551) );
  OR2_X1 U658 ( .A1(n374), .A2(n552), .ZN(n553) );
  NOR2_X1 U659 ( .A1(G900), .A2(n553), .ZN(n554) );
  NOR2_X1 U660 ( .A1(n555), .A2(n554), .ZN(n567) );
  NOR2_X1 U661 ( .A1(n567), .A2(n556), .ZN(n558) );
  NAND2_X1 U662 ( .A1(n558), .A2(n557), .ZN(n579) );
  NAND2_X1 U663 ( .A1(n561), .A2(n560), .ZN(n575) );
  INV_X1 U664 ( .A(n603), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n638), .A2(n637), .ZN(n562) );
  XNOR2_X1 U666 ( .A(n562), .B(KEYINPUT107), .ZN(n636) );
  NAND2_X1 U667 ( .A1(n640), .A2(n636), .ZN(n563) );
  XNOR2_X1 U668 ( .A(n564), .B(KEYINPUT42), .ZN(n738) );
  NAND2_X1 U669 ( .A1(n628), .A2(n637), .ZN(n565) );
  XNOR2_X1 U670 ( .A(KEYINPUT30), .B(n565), .ZN(n570) );
  XNOR2_X1 U671 ( .A(n568), .B(KEYINPUT77), .ZN(n569) );
  NOR2_X1 U672 ( .A1(n738), .A2(n737), .ZN(n573) );
  XNOR2_X1 U673 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n572) );
  XNOR2_X1 U674 ( .A(n573), .B(n572), .ZN(n598) );
  XNOR2_X1 U675 ( .A(KEYINPUT67), .B(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U676 ( .A1(n576), .A2(n586), .ZN(n585) );
  INV_X1 U677 ( .A(n582), .ZN(n583) );
  NAND2_X1 U678 ( .A1(n584), .A2(n583), .ZN(n688) );
  NAND2_X1 U679 ( .A1(n585), .A2(n688), .ZN(n594) );
  INV_X1 U680 ( .A(KEYINPUT47), .ZN(n587) );
  OR2_X1 U681 ( .A1(n587), .A2(n586), .ZN(n592) );
  NOR2_X1 U682 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n677) );
  XNOR2_X1 U684 ( .A(n599), .B(KEYINPUT48), .ZN(n608) );
  NOR2_X1 U685 ( .A1(n621), .A2(n600), .ZN(n601) );
  XNOR2_X1 U686 ( .A(n601), .B(KEYINPUT43), .ZN(n602) );
  NOR2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n690) );
  NAND2_X1 U688 ( .A1(n605), .A2(n604), .ZN(n689) );
  NAND2_X1 U689 ( .A1(KEYINPUT2), .A2(n610), .ZN(n611) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n656) );
  XNOR2_X1 U691 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT55), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n657), .B(n656), .ZN(n655) );
  NAND2_X1 U694 ( .A1(n632), .A2(n645), .ZN(n653) );
  XNOR2_X1 U695 ( .A(KEYINPUT52), .B(KEYINPUT115), .ZN(n650) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U697 ( .A(KEYINPUT49), .B(n620), .ZN(n626) );
  OR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT50), .ZN(n624) );
  XNOR2_X1 U700 ( .A(KEYINPUT112), .B(n624), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n631), .B(KEYINPUT51), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n648) );
  INV_X1 U706 ( .A(n634), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n644) );
  NOR2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U709 ( .A(KEYINPUT113), .B(n639), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U711 ( .A(KEYINPUT114), .B(n642), .ZN(n643) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U714 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n650), .B(n649), .ZN(n651) );
  AND2_X1 U716 ( .A1(n653), .A2(n347), .ZN(n658) );
  AND2_X1 U717 ( .A1(KEYINPUT82), .A2(n658), .ZN(n654) );
  NAND2_X1 U718 ( .A1(n655), .A2(n654), .ZN(n663) );
  AND2_X1 U719 ( .A1(n657), .A2(n656), .ZN(n661) );
  INV_X1 U720 ( .A(KEYINPUT82), .ZN(n659) );
  NAND2_X1 U721 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U722 ( .A1(G953), .A2(n664), .ZN(n667) );
  INV_X1 U723 ( .A(KEYINPUT53), .ZN(n665) );
  XNOR2_X1 U724 ( .A(n665), .B(KEYINPUT117), .ZN(n666) );
  XNOR2_X1 U725 ( .A(G101), .B(n668), .ZN(G3) );
  NAND2_X1 U726 ( .A1(n670), .A2(n681), .ZN(n669) );
  XNOR2_X1 U727 ( .A(n669), .B(G104), .ZN(G6) );
  XOR2_X1 U728 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n672) );
  INV_X1 U729 ( .A(n674), .ZN(n684) );
  NAND2_X1 U730 ( .A1(n670), .A2(n684), .ZN(n671) );
  XNOR2_X1 U731 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U732 ( .A(G107), .B(n673), .ZN(G9) );
  NOR2_X1 U733 ( .A1(n674), .A2(n678), .ZN(n676) );
  XNOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .ZN(n675) );
  XNOR2_X1 U735 ( .A(n676), .B(n675), .ZN(G30) );
  XNOR2_X1 U736 ( .A(G143), .B(n677), .ZN(G45) );
  NOR2_X1 U737 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U738 ( .A(G146), .B(n680), .Z(G48) );
  XOR2_X1 U739 ( .A(G113), .B(KEYINPUT111), .Z(n683) );
  NAND2_X1 U740 ( .A1(n685), .A2(n681), .ZN(n682) );
  XNOR2_X1 U741 ( .A(n683), .B(n682), .ZN(G15) );
  NAND2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U743 ( .A(n686), .B(G116), .ZN(G18) );
  XOR2_X1 U744 ( .A(G125), .B(KEYINPUT37), .Z(n687) );
  XNOR2_X1 U745 ( .A(n688), .B(n687), .ZN(G27) );
  XNOR2_X1 U746 ( .A(G134), .B(n689), .ZN(G36) );
  XOR2_X1 U747 ( .A(G140), .B(n690), .Z(G42) );
  XOR2_X1 U748 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n692) );
  XNOR2_X1 U749 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n691) );
  XNOR2_X1 U750 ( .A(n692), .B(n691), .ZN(n693) );
  XOR2_X1 U751 ( .A(n694), .B(n693), .Z(n696) );
  NAND2_X1 U752 ( .A1(n704), .A2(G469), .ZN(n695) );
  XNOR2_X1 U753 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U754 ( .A1(n708), .A2(n697), .ZN(G54) );
  XNOR2_X1 U755 ( .A(KEYINPUT59), .B(KEYINPUT122), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n698), .B(KEYINPUT121), .ZN(n699) );
  XNOR2_X1 U757 ( .A(KEYINPUT60), .B(n701), .ZN(G60) );
  NAND2_X1 U758 ( .A1(G217), .A2(n704), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(G66) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n709) );
  XNOR2_X1 U762 ( .A(KEYINPUT61), .B(n709), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n710), .A2(G898), .ZN(n713) );
  NAND2_X1 U764 ( .A1(n711), .A2(n374), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n718) );
  XNOR2_X1 U766 ( .A(n714), .B(G101), .ZN(n715) );
  NAND2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U768 ( .A(n718), .B(n717), .Z(G69) );
  XOR2_X1 U769 ( .A(n719), .B(KEYINPUT125), .Z(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U771 ( .A(n723), .B(n722), .Z(n727) );
  XOR2_X1 U772 ( .A(n727), .B(n724), .Z(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(n374), .ZN(n732) );
  XNOR2_X1 U774 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G900), .ZN(n729) );
  XNOR2_X1 U776 ( .A(KEYINPUT126), .B(n729), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n730), .A2(G953), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n732), .A2(n731), .ZN(G72) );
  XOR2_X1 U779 ( .A(n733), .B(G119), .Z(G21) );
  XOR2_X1 U780 ( .A(n734), .B(G110), .Z(n735) );
  XNOR2_X1 U781 ( .A(KEYINPUT110), .B(n735), .ZN(G12) );
  XNOR2_X1 U782 ( .A(G122), .B(n736), .ZN(G24) );
  XOR2_X1 U783 ( .A(n737), .B(G131), .Z(G33) );
  XNOR2_X1 U784 ( .A(G137), .B(KEYINPUT127), .ZN(n739) );
  XNOR2_X1 U785 ( .A(n739), .B(n738), .ZN(G39) );
endmodule

