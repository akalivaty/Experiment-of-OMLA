

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749;

  NOR2_X1 U378 ( .A1(n696), .A2(n717), .ZN(n358) );
  AND2_X1 U379 ( .A1(n391), .A2(n390), .ZN(n389) );
  NAND2_X1 U380 ( .A1(n633), .A2(n557), .ZN(n596) );
  XNOR2_X1 U381 ( .A(n422), .B(n526), .ZN(n688) );
  BUF_X1 U382 ( .A(G107), .Z(n357) );
  XNOR2_X1 U383 ( .A(n725), .B(n486), .ZN(n381) );
  XNOR2_X2 U384 ( .A(n417), .B(n367), .ZN(n527) );
  NAND2_X2 U385 ( .A1(n427), .A2(n370), .ZN(n429) );
  XNOR2_X1 U386 ( .A(n358), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U387 ( .A(G953), .ZN(n741) );
  AND2_X2 U388 ( .A1(n718), .A2(n365), .ZN(n428) );
  OR2_X2 U389 ( .A1(n552), .A2(n664), .ZN(n555) );
  XNOR2_X2 U390 ( .A(n514), .B(n513), .ZN(n552) );
  NOR2_X2 U391 ( .A1(n421), .A2(n362), .ZN(n379) );
  AND2_X2 U392 ( .A1(n745), .A2(KEYINPUT44), .ZN(n362) );
  XOR2_X2 U393 ( .A(n541), .B(KEYINPUT100), .Z(n542) );
  XNOR2_X2 U394 ( .A(n470), .B(n469), .ZN(n541) );
  XNOR2_X2 U395 ( .A(n400), .B(KEYINPUT19), .ZN(n387) );
  NAND2_X2 U396 ( .A1(n563), .A2(n652), .ZN(n400) );
  XNOR2_X1 U397 ( .A(n592), .B(KEYINPUT40), .ZN(n747) );
  XOR2_X2 U398 ( .A(G143), .B(G128), .Z(n471) );
  NAND2_X1 U399 ( .A1(n537), .A2(n556), .ZN(n422) );
  INV_X1 U400 ( .A(KEYINPUT16), .ZN(n413) );
  NOR2_X1 U401 ( .A1(n587), .A2(n586), .ZN(n408) );
  XNOR2_X1 U402 ( .A(n594), .B(KEYINPUT42), .ZN(n749) );
  XNOR2_X1 U403 ( .A(n414), .B(KEYINPUT41), .ZN(n686) );
  BUF_X1 U404 ( .A(n527), .Z(n538) );
  INV_X1 U405 ( .A(n635), .ZN(n633) );
  XNOR2_X1 U406 ( .A(KEYINPUT104), .B(n544), .ZN(n635) );
  XNOR2_X1 U407 ( .A(n692), .B(n693), .ZN(n694) );
  XNOR2_X1 U408 ( .A(n383), .B(n384), .ZN(n380) );
  XNOR2_X1 U409 ( .A(n439), .B(n437), .ZN(n384) );
  XNOR2_X1 U410 ( .A(n734), .B(n424), .ZN(n486) );
  XNOR2_X1 U411 ( .A(n480), .B(n413), .ZN(n382) );
  XNOR2_X1 U412 ( .A(n471), .B(n441), .ZN(n734) );
  XNOR2_X1 U413 ( .A(n440), .B(KEYINPUT3), .ZN(n412) );
  AND2_X1 U414 ( .A1(n430), .A2(n429), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n486), .B(n485), .ZN(n498) );
  XNOR2_X1 U416 ( .A(n733), .B(G146), .ZN(n485) );
  XOR2_X1 U417 ( .A(G137), .B(KEYINPUT69), .Z(n499) );
  XNOR2_X1 U418 ( .A(n724), .B(KEYINPUT75), .ZN(n492) );
  NAND2_X1 U419 ( .A1(n403), .A2(n516), .ZN(n402) );
  INV_X1 U420 ( .A(n556), .ZN(n403) );
  XNOR2_X1 U421 ( .A(n410), .B(G469), .ZN(n576) );
  OR2_X1 U422 ( .A1(n698), .A2(G902), .ZN(n410) );
  OR2_X1 U423 ( .A1(n612), .A2(G902), .ZN(n404) );
  XNOR2_X1 U424 ( .A(G137), .B(G116), .ZN(n487) );
  XOR2_X1 U425 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n488) );
  XNOR2_X1 U426 ( .A(G119), .B(G113), .ZN(n411) );
  INV_X1 U427 ( .A(KEYINPUT4), .ZN(n441) );
  XOR2_X1 U428 ( .A(G146), .B(G125), .Z(n454) );
  NOR2_X1 U429 ( .A1(n555), .A2(n567), .ZN(n575) );
  NAND2_X1 U430 ( .A1(n653), .A2(n652), .ZN(n656) );
  XNOR2_X1 U431 ( .A(n600), .B(KEYINPUT38), .ZN(n653) );
  NAND2_X1 U432 ( .A1(n393), .A2(n392), .ZN(n391) );
  NOR2_X1 U433 ( .A1(n688), .A2(n368), .ZN(n392) );
  XNOR2_X1 U434 ( .A(n576), .B(n409), .ZN(n666) );
  INV_X1 U435 ( .A(KEYINPUT1), .ZN(n409) );
  XNOR2_X1 U436 ( .A(n501), .B(n500), .ZN(n735) );
  XNOR2_X1 U437 ( .A(n497), .B(n498), .ZN(n698) );
  INV_X1 U438 ( .A(n402), .ZN(n397) );
  XNOR2_X1 U439 ( .A(n564), .B(n423), .ZN(n556) );
  NAND2_X1 U440 ( .A1(n426), .A2(n425), .ZN(n386) );
  AND2_X1 U441 ( .A1(n483), .A2(n525), .ZN(n425) );
  INV_X1 U442 ( .A(n527), .ZN(n426) );
  BUF_X1 U443 ( .A(n359), .Z(n713) );
  NOR2_X1 U444 ( .A1(G952), .A2(n741), .ZN(n717) );
  XNOR2_X1 U445 ( .A(KEYINPUT46), .B(KEYINPUT86), .ZN(n415) );
  NAND2_X1 U446 ( .A1(n747), .A2(n749), .ZN(n416) );
  XOR2_X1 U447 ( .A(G902), .B(KEYINPUT15), .Z(n611) );
  XNOR2_X1 U448 ( .A(G131), .B(G134), .ZN(n484) );
  AND2_X1 U449 ( .A1(G227), .A2(n741), .ZN(n432) );
  INV_X1 U450 ( .A(KEYINPUT64), .ZN(n418) );
  OR2_X1 U451 ( .A1(G237), .A2(G902), .ZN(n444) );
  NAND2_X1 U452 ( .A1(n387), .A2(n450), .ZN(n417) );
  NOR2_X1 U453 ( .A1(n449), .A2(n431), .ZN(n450) );
  XNOR2_X1 U454 ( .A(n489), .B(n364), .ZN(n371) );
  NAND2_X1 U455 ( .A1(n436), .A2(n435), .ZN(n724) );
  INV_X1 U456 ( .A(G122), .ZN(n419) );
  XOR2_X1 U457 ( .A(KEYINPUT8), .B(n477), .Z(n507) );
  NAND2_X1 U458 ( .A1(G234), .A2(n741), .ZN(n477) );
  XNOR2_X1 U459 ( .A(n455), .B(G140), .ZN(n501) );
  XNOR2_X1 U460 ( .A(G113), .B(G143), .ZN(n458) );
  XOR2_X1 U461 ( .A(G104), .B(G122), .Z(n459) );
  XNOR2_X1 U462 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n461) );
  XNOR2_X1 U463 ( .A(KEYINPUT97), .B(KEYINPUT11), .ZN(n460) );
  XNOR2_X1 U464 ( .A(KEYINPUT74), .B(KEYINPUT17), .ZN(n437) );
  XNOR2_X1 U465 ( .A(KEYINPUT68), .B(G101), .ZN(n424) );
  XNOR2_X1 U466 ( .A(n438), .B(n492), .ZN(n383) );
  XNOR2_X1 U467 ( .A(n454), .B(KEYINPUT18), .ZN(n438) );
  OR2_X1 U468 ( .A1(n656), .A2(n655), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n531), .B(n530), .ZN(n551) );
  NAND2_X1 U470 ( .A1(n389), .A2(n361), .ZN(n531) );
  XNOR2_X1 U471 ( .A(n376), .B(n375), .ZN(n577) );
  INV_X1 U472 ( .A(KEYINPUT28), .ZN(n375) );
  NOR2_X1 U473 ( .A1(n571), .A2(n570), .ZN(n589) );
  BUF_X1 U474 ( .A(n563), .Z(n588) );
  XNOR2_X1 U475 ( .A(n512), .B(KEYINPUT25), .ZN(n513) );
  NAND2_X1 U476 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U477 ( .A(n717), .ZN(n373) );
  XNOR2_X1 U478 ( .A(n701), .B(n702), .ZN(n374) );
  AND2_X1 U479 ( .A1(n610), .A2(n748), .ZN(n360) );
  AND2_X1 U480 ( .A1(n388), .A2(n572), .ZN(n361) );
  XOR2_X1 U481 ( .A(n416), .B(n415), .Z(n363) );
  NAND2_X1 U482 ( .A1(n491), .A2(G210), .ZN(n364) );
  AND2_X1 U483 ( .A1(n748), .A2(n611), .ZN(n365) );
  XOR2_X1 U484 ( .A(G472), .B(KEYINPUT77), .Z(n366) );
  XOR2_X1 U485 ( .A(KEYINPUT89), .B(KEYINPUT0), .Z(n367) );
  XNOR2_X1 U486 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n368) );
  XOR2_X1 U487 ( .A(n595), .B(KEYINPUT71), .Z(n369) );
  XOR2_X1 U488 ( .A(KEYINPUT67), .B(n608), .Z(n370) );
  NAND2_X1 U489 ( .A1(n428), .A2(n610), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n371), .B(n490), .ZN(n405) );
  XNOR2_X1 U491 ( .A(n372), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U492 ( .A1(n708), .A2(n717), .ZN(n372) );
  AND2_X1 U493 ( .A1(n374), .A2(n373), .ZN(G54) );
  NAND2_X1 U494 ( .A1(n746), .A2(n626), .ZN(n522) );
  OR2_X2 U495 ( .A1(n394), .A2(n398), .ZN(n746) );
  NAND2_X1 U496 ( .A1(n575), .A2(n564), .ZN(n376) );
  NAND2_X1 U497 ( .A1(n518), .A2(n517), .ZN(n385) );
  AND2_X2 U498 ( .A1(n430), .A2(n429), .ZN(n703) );
  XNOR2_X2 U499 ( .A(n377), .B(KEYINPUT45), .ZN(n718) );
  NAND2_X1 U500 ( .A1(n379), .A2(n378), .ZN(n377) );
  XNOR2_X1 U501 ( .A(n524), .B(n418), .ZN(n378) );
  XNOR2_X2 U502 ( .A(n381), .B(n380), .ZN(n692) );
  XNOR2_X2 U503 ( .A(n382), .B(n490), .ZN(n725) );
  XNOR2_X2 U504 ( .A(n412), .B(n411), .ZN(n490) );
  NAND2_X1 U505 ( .A1(n385), .A2(n399), .ZN(n398) );
  XNOR2_X2 U506 ( .A(n386), .B(KEYINPUT22), .ZN(n518) );
  NAND2_X1 U507 ( .A1(n593), .A2(n387), .ZN(n579) );
  NAND2_X1 U508 ( .A1(n688), .A2(n368), .ZN(n388) );
  NAND2_X1 U509 ( .A1(n535), .A2(n368), .ZN(n390) );
  INV_X1 U510 ( .A(n535), .ZN(n393) );
  XNOR2_X2 U511 ( .A(n538), .B(KEYINPUT92), .ZN(n535) );
  NOR2_X1 U512 ( .A1(n518), .A2(n395), .ZN(n394) );
  INV_X1 U513 ( .A(n517), .ZN(n396) );
  NAND2_X1 U514 ( .A1(n402), .A2(n517), .ZN(n399) );
  NOR2_X1 U515 ( .A1(n558), .A2(n400), .ZN(n561) );
  NAND2_X1 U516 ( .A1(n580), .A2(n401), .ZN(n581) );
  NAND2_X1 U517 ( .A1(n401), .A2(n627), .ZN(n628) );
  NAND2_X1 U518 ( .A1(n401), .A2(n633), .ZN(n634) );
  NAND2_X1 U519 ( .A1(n583), .A2(n401), .ZN(n584) );
  XNOR2_X2 U520 ( .A(n579), .B(KEYINPUT81), .ZN(n401) );
  NOR2_X1 U521 ( .A1(n518), .A2(n556), .ZN(n546) );
  XNOR2_X2 U522 ( .A(n404), .B(n366), .ZN(n564) );
  XNOR2_X1 U523 ( .A(n405), .B(n498), .ZN(n612) );
  XNOR2_X1 U524 ( .A(n406), .B(n369), .ZN(n602) );
  NAND2_X1 U525 ( .A1(n407), .A2(n363), .ZN(n406) );
  XNOR2_X1 U526 ( .A(n408), .B(KEYINPUT72), .ZN(n407) );
  NOR2_X1 U527 ( .A1(n666), .A2(n667), .ZN(n537) );
  NOR2_X1 U528 ( .A1(n551), .A2(KEYINPUT44), .ZN(n532) );
  INV_X1 U529 ( .A(n649), .ZN(n430) );
  XNOR2_X2 U530 ( .A(n420), .B(n419), .ZN(n480) );
  XNOR2_X2 U531 ( .A(G116), .B(G107), .ZN(n420) );
  NAND2_X1 U532 ( .A1(n550), .A2(n549), .ZN(n421) );
  INV_X1 U533 ( .A(KEYINPUT6), .ZN(n423) );
  NOR2_X2 U534 ( .A1(n717), .A2(n615), .ZN(n617) );
  AND2_X1 U535 ( .A1(G953), .A2(G898), .ZN(n431) );
  XNOR2_X1 U536 ( .A(n499), .B(n432), .ZN(n493) );
  INV_X1 U537 ( .A(KEYINPUT13), .ZN(n468) );
  XNOR2_X1 U538 ( .A(n559), .B(KEYINPUT36), .ZN(n560) );
  XNOR2_X1 U539 ( .A(n468), .B(G475), .ZN(n469) );
  XNOR2_X1 U540 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U541 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U542 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U543 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U544 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U545 ( .A(KEYINPUT63), .B(KEYINPUT111), .ZN(n616) );
  INV_X1 U546 ( .A(G104), .ZN(n433) );
  NAND2_X1 U547 ( .A1(G110), .A2(n433), .ZN(n436) );
  INV_X1 U548 ( .A(G110), .ZN(n434) );
  NAND2_X1 U549 ( .A1(n434), .A2(G104), .ZN(n435) );
  AND2_X1 U550 ( .A1(G224), .A2(n741), .ZN(n439) );
  XNOR2_X2 U551 ( .A(KEYINPUT91), .B(KEYINPUT73), .ZN(n440) );
  NOR2_X2 U552 ( .A1(n692), .A2(n611), .ZN(n443) );
  NAND2_X1 U553 ( .A1(G210), .A2(n444), .ZN(n442) );
  XNOR2_X2 U554 ( .A(n443), .B(n442), .ZN(n563) );
  NAND2_X1 U555 ( .A1(G214), .A2(n444), .ZN(n652) );
  NAND2_X1 U556 ( .A1(G234), .A2(G237), .ZN(n445) );
  XNOR2_X1 U557 ( .A(n445), .B(KEYINPUT14), .ZN(n680) );
  OR2_X1 U558 ( .A1(n741), .A2(G902), .ZN(n446) );
  NAND2_X1 U559 ( .A1(n680), .A2(n446), .ZN(n448) );
  NOR2_X1 U560 ( .A1(G953), .A2(G952), .ZN(n447) );
  NOR2_X1 U561 ( .A1(n448), .A2(n447), .ZN(n554) );
  INV_X1 U562 ( .A(n554), .ZN(n449) );
  INV_X1 U563 ( .A(n611), .ZN(n451) );
  NAND2_X1 U564 ( .A1(n451), .A2(G234), .ZN(n452) );
  XNOR2_X1 U565 ( .A(n452), .B(KEYINPUT20), .ZN(n511) );
  NAND2_X1 U566 ( .A1(n511), .A2(G221), .ZN(n453) );
  XNOR2_X1 U567 ( .A(KEYINPUT21), .B(n453), .ZN(n664) );
  XOR2_X1 U568 ( .A(KEYINPUT94), .B(n664), .Z(n525) );
  XNOR2_X1 U569 ( .A(n454), .B(KEYINPUT10), .ZN(n455) );
  XOR2_X1 U570 ( .A(G131), .B(KEYINPUT12), .Z(n457) );
  NOR2_X1 U571 ( .A1(G953), .A2(G237), .ZN(n491) );
  NAND2_X1 U572 ( .A1(G214), .A2(n491), .ZN(n456) );
  XNOR2_X1 U573 ( .A(n457), .B(n456), .ZN(n466) );
  XNOR2_X1 U574 ( .A(n459), .B(n458), .ZN(n464) );
  INV_X1 U575 ( .A(n460), .ZN(n462) );
  XNOR2_X1 U576 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U577 ( .A(n464), .B(n463), .Z(n465) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U579 ( .A(n501), .B(n467), .ZN(n705) );
  NOR2_X1 U580 ( .A1(n705), .A2(G902), .ZN(n470) );
  XNOR2_X1 U581 ( .A(n471), .B(KEYINPUT9), .ZN(n472) );
  XNOR2_X1 U582 ( .A(n472), .B(KEYINPUT7), .ZN(n476) );
  XOR2_X1 U583 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n474) );
  XNOR2_X1 U584 ( .A(G134), .B(KEYINPUT101), .ZN(n473) );
  XNOR2_X1 U585 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U586 ( .A(n476), .B(n475), .Z(n479) );
  NAND2_X1 U587 ( .A1(G217), .A2(n507), .ZN(n478) );
  XNOR2_X1 U588 ( .A(n479), .B(n478), .ZN(n481) );
  XNOR2_X1 U589 ( .A(n480), .B(n481), .ZN(n709) );
  NOR2_X1 U590 ( .A1(n709), .A2(G902), .ZN(n482) );
  XNOR2_X1 U591 ( .A(n482), .B(G478), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n541), .A2(n543), .ZN(n655) );
  INV_X1 U593 ( .A(n655), .ZN(n483) );
  XNOR2_X1 U594 ( .A(n484), .B(KEYINPUT70), .ZN(n733) );
  XNOR2_X1 U595 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U596 ( .A(n357), .B(G140), .ZN(n496) );
  XNOR2_X1 U597 ( .A(n492), .B(KEYINPUT74), .ZN(n494) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U599 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U600 ( .A(n499), .ZN(n500) );
  XNOR2_X1 U601 ( .A(G128), .B(G110), .ZN(n502) );
  XNOR2_X1 U602 ( .A(n502), .B(KEYINPUT79), .ZN(n506) );
  XOR2_X1 U603 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n504) );
  XNOR2_X1 U604 ( .A(G119), .B(KEYINPUT24), .ZN(n503) );
  XNOR2_X1 U605 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U606 ( .A(n506), .B(n505), .Z(n509) );
  NAND2_X1 U607 ( .A1(G221), .A2(n507), .ZN(n508) );
  XNOR2_X1 U608 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n735), .B(n510), .ZN(n715) );
  NOR2_X1 U610 ( .A1(n715), .A2(G902), .ZN(n514) );
  NAND2_X1 U611 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U612 ( .A(KEYINPUT105), .B(n552), .ZN(n663) );
  INV_X1 U613 ( .A(n663), .ZN(n515) );
  NOR2_X1 U614 ( .A1(n666), .A2(n515), .ZN(n516) );
  XOR2_X1 U615 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n517) );
  INV_X1 U616 ( .A(n666), .ZN(n597) );
  NOR2_X1 U617 ( .A1(n518), .A2(n597), .ZN(n520) );
  NOR2_X1 U618 ( .A1(n564), .A2(n552), .ZN(n519) );
  NAND2_X1 U619 ( .A1(n520), .A2(n519), .ZN(n626) );
  INV_X1 U620 ( .A(KEYINPUT88), .ZN(n521) );
  XNOR2_X1 U621 ( .A(n522), .B(n521), .ZN(n533) );
  INV_X1 U622 ( .A(KEYINPUT44), .ZN(n523) );
  NOR2_X1 U623 ( .A1(n533), .A2(n523), .ZN(n524) );
  XOR2_X1 U624 ( .A(KEYINPUT90), .B(KEYINPUT33), .Z(n526) );
  NAND2_X1 U625 ( .A1(n525), .A2(n552), .ZN(n667) );
  NOR2_X1 U626 ( .A1(n541), .A2(n543), .ZN(n572) );
  XOR2_X1 U627 ( .A(KEYINPUT35), .B(KEYINPUT84), .Z(n529) );
  INV_X1 U628 ( .A(KEYINPUT80), .ZN(n528) );
  NAND2_X1 U629 ( .A1(n533), .A2(n532), .ZN(n550) );
  INV_X1 U630 ( .A(n576), .ZN(n534) );
  NOR2_X1 U631 ( .A1(n534), .A2(n667), .ZN(n568) );
  NOR2_X1 U632 ( .A1(n535), .A2(n564), .ZN(n536) );
  NAND2_X1 U633 ( .A1(n568), .A2(n536), .ZN(n622) );
  NAND2_X1 U634 ( .A1(n564), .A2(n537), .ZN(n674) );
  NOR2_X1 U635 ( .A1(n538), .A2(n674), .ZN(n540) );
  XNOR2_X1 U636 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n539) );
  XNOR2_X1 U637 ( .A(n540), .B(n539), .ZN(n639) );
  NAND2_X1 U638 ( .A1(n622), .A2(n639), .ZN(n545) );
  NOR2_X1 U639 ( .A1(n543), .A2(n542), .ZN(n627) );
  NAND2_X1 U640 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X2 U641 ( .A1(n627), .A2(n633), .ZN(n657) );
  INV_X1 U642 ( .A(n657), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n545), .A2(n574), .ZN(n548) );
  NOR2_X1 U644 ( .A1(n663), .A2(n597), .ZN(n547) );
  NAND2_X1 U645 ( .A1(n546), .A2(n547), .ZN(n618) );
  AND2_X1 U646 ( .A1(n548), .A2(n618), .ZN(n549) );
  BUF_X2 U647 ( .A(n551), .Z(n745) );
  NAND2_X1 U648 ( .A1(G953), .A2(G900), .ZN(n553) );
  NAND2_X1 U649 ( .A1(n554), .A2(n553), .ZN(n567) );
  AND2_X1 U650 ( .A1(n575), .A2(n556), .ZN(n557) );
  XNOR2_X1 U651 ( .A(KEYINPUT108), .B(n596), .ZN(n558) );
  INV_X1 U652 ( .A(KEYINPUT109), .ZN(n559) );
  NAND2_X1 U653 ( .A1(n562), .A2(n597), .ZN(n642) );
  NAND2_X1 U654 ( .A1(n652), .A2(n564), .ZN(n565) );
  XNOR2_X1 U655 ( .A(n565), .B(KEYINPUT30), .ZN(n566) );
  XNOR2_X1 U656 ( .A(n566), .B(KEYINPUT106), .ZN(n571) );
  INV_X1 U657 ( .A(n567), .ZN(n569) );
  NAND2_X1 U658 ( .A1(n569), .A2(n568), .ZN(n570) );
  AND2_X1 U659 ( .A1(n589), .A2(n572), .ZN(n573) );
  NAND2_X1 U660 ( .A1(n588), .A2(n573), .ZN(n632) );
  NAND2_X1 U661 ( .A1(n642), .A2(n632), .ZN(n587) );
  AND2_X1 U662 ( .A1(n574), .A2(KEYINPUT78), .ZN(n580) );
  NAND2_X1 U663 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U664 ( .A(n578), .B(KEYINPUT107), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n581), .A2(KEYINPUT47), .ZN(n585) );
  XNOR2_X1 U666 ( .A(KEYINPUT78), .B(n657), .ZN(n582) );
  NOR2_X1 U667 ( .A1(KEYINPUT47), .A2(n582), .ZN(n583) );
  NAND2_X1 U668 ( .A1(n585), .A2(n584), .ZN(n586) );
  INV_X1 U669 ( .A(n588), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n589), .A2(n653), .ZN(n591) );
  XOR2_X1 U671 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n590) );
  XNOR2_X1 U672 ( .A(n591), .B(n590), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n603), .A2(n633), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n593), .A2(n686), .ZN(n594) );
  XNOR2_X1 U675 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n595) );
  NOR2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n598), .A2(n652), .ZN(n599) );
  XNOR2_X1 U678 ( .A(n599), .B(KEYINPUT43), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n646) );
  NAND2_X1 U680 ( .A1(n602), .A2(n646), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n627), .A2(n603), .ZN(n604) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT110), .ZN(n748) );
  NAND2_X1 U683 ( .A1(n748), .A2(KEYINPUT2), .ZN(n605) );
  XNOR2_X1 U684 ( .A(KEYINPUT82), .B(n605), .ZN(n606) );
  NOR2_X1 U685 ( .A1(n609), .A2(n606), .ZN(n607) );
  AND2_X1 U686 ( .A1(n718), .A2(n607), .ZN(n649) );
  NAND2_X1 U687 ( .A1(n611), .A2(KEYINPUT2), .ZN(n608) );
  INV_X1 U688 ( .A(n609), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n703), .A2(G472), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n612), .B(KEYINPUT62), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n617), .B(n616), .ZN(G57) );
  XNOR2_X1 U692 ( .A(G101), .B(n618), .ZN(G3) );
  NOR2_X1 U693 ( .A1(n635), .A2(n622), .ZN(n619) );
  XOR2_X1 U694 ( .A(G104), .B(n619), .Z(G6) );
  XOR2_X1 U695 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n621) );
  XNOR2_X1 U696 ( .A(n357), .B(KEYINPUT26), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n621), .B(n620), .ZN(n624) );
  INV_X1 U698 ( .A(n627), .ZN(n638) );
  NOR2_X1 U699 ( .A1(n638), .A2(n622), .ZN(n623) );
  XOR2_X1 U700 ( .A(n624), .B(n623), .Z(G9) );
  XOR2_X1 U701 ( .A(G110), .B(KEYINPUT113), .Z(n625) );
  XNOR2_X1 U702 ( .A(n626), .B(n625), .ZN(G12) );
  XOR2_X1 U703 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n629) );
  XNOR2_X1 U704 ( .A(n629), .B(n628), .ZN(n631) );
  XOR2_X1 U705 ( .A(G128), .B(KEYINPUT114), .Z(n630) );
  XNOR2_X1 U706 ( .A(n631), .B(n630), .ZN(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(n632), .ZN(G45) );
  XNOR2_X1 U708 ( .A(n634), .B(G146), .ZN(G48) );
  NOR2_X1 U709 ( .A1(n635), .A2(n639), .ZN(n636) );
  XOR2_X1 U710 ( .A(KEYINPUT116), .B(n636), .Z(n637) );
  XNOR2_X1 U711 ( .A(G113), .B(n637), .ZN(G15) );
  NOR2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n641) );
  XNOR2_X1 U713 ( .A(G116), .B(KEYINPUT117), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G18) );
  BUF_X1 U715 ( .A(n642), .Z(n644) );
  XOR2_X1 U716 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n643) );
  XNOR2_X1 U717 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U718 ( .A(G125), .B(n645), .ZN(G27) );
  XNOR2_X1 U719 ( .A(G140), .B(n646), .ZN(G42) );
  NOR2_X1 U720 ( .A1(KEYINPUT2), .A2(n360), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT83), .ZN(n651) );
  NOR2_X1 U722 ( .A1(n718), .A2(KEYINPUT2), .ZN(n648) );
  NOR2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n685) );
  NOR2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(KEYINPUT120), .ZN(n661) );
  NOR2_X1 U730 ( .A1(n688), .A2(n661), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT121), .ZN(n678) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U733 ( .A(KEYINPUT49), .B(n665), .Z(n672) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(KEYINPUT50), .ZN(n669) );
  XNOR2_X1 U736 ( .A(KEYINPUT119), .B(n669), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n564), .A2(n670), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(n675), .Z(n676) );
  NAND2_X1 U741 ( .A1(n676), .A2(n686), .ZN(n677) );
  NAND2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U743 ( .A(KEYINPUT52), .B(n679), .Z(n682) );
  NAND2_X1 U744 ( .A1(G952), .A2(n680), .ZN(n681) );
  NOR2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U746 ( .A1(G953), .A2(n683), .ZN(n684) );
  NAND2_X1 U747 ( .A1(n685), .A2(n684), .ZN(n690) );
  INV_X1 U748 ( .A(n686), .ZN(n687) );
  NOR2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U751 ( .A(KEYINPUT53), .B(n691), .ZN(G75) );
  NAND2_X1 U752 ( .A1(n703), .A2(G210), .ZN(n695) );
  XOR2_X1 U753 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n693) );
  XNOR2_X1 U754 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U755 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n698), .B(KEYINPUT57), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U758 ( .A1(n713), .A2(G469), .ZN(n701) );
  NAND2_X1 U759 ( .A1(n359), .A2(G475), .ZN(n707) );
  XOR2_X1 U760 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n704) );
  XOR2_X1 U761 ( .A(n709), .B(KEYINPUT123), .Z(n711) );
  NAND2_X1 U762 ( .A1(n713), .A2(G478), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U764 ( .A1(n717), .A2(n712), .ZN(G63) );
  NAND2_X1 U765 ( .A1(G217), .A2(n713), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U768 ( .A1(n718), .A2(n741), .ZN(n723) );
  NAND2_X1 U769 ( .A1(G224), .A2(G953), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n719), .B(KEYINPUT61), .ZN(n720) );
  XNOR2_X1 U771 ( .A(KEYINPUT124), .B(n720), .ZN(n721) );
  NAND2_X1 U772 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n732) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n726), .B(KEYINPUT125), .ZN(n727) );
  XNOR2_X1 U776 ( .A(n727), .B(G101), .ZN(n729) );
  NOR2_X1 U777 ( .A1(n741), .A2(G898), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U779 ( .A(KEYINPUT126), .B(n730), .ZN(n731) );
  XNOR2_X1 U780 ( .A(n732), .B(n731), .ZN(G69) );
  XNOR2_X1 U781 ( .A(n734), .B(n733), .ZN(n736) );
  XNOR2_X1 U782 ( .A(n736), .B(n735), .ZN(n740) );
  XNOR2_X1 U783 ( .A(n740), .B(KEYINPUT127), .ZN(n737) );
  XNOR2_X1 U784 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U785 ( .A1(G900), .A2(n738), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n739), .A2(G953), .ZN(n744) );
  XNOR2_X1 U787 ( .A(n740), .B(n360), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n744), .A2(n743), .ZN(G72) );
  XOR2_X1 U790 ( .A(n745), .B(G122), .Z(G24) );
  XNOR2_X1 U791 ( .A(G119), .B(n746), .ZN(G21) );
  XNOR2_X1 U792 ( .A(n747), .B(G131), .ZN(G33) );
  XNOR2_X1 U793 ( .A(G134), .B(n748), .ZN(G36) );
  XNOR2_X1 U794 ( .A(n749), .B(G137), .ZN(G39) );
endmodule

