//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946;
  INV_X1    g000(.A(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G141gat), .B(G148gat), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  XOR2_X1   g011(.A(G127gat), .B(G134gat), .Z(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G141gat), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT78), .B(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n204), .A2(KEYINPUT79), .A3(new_n205), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n228));
  AND4_X1   g027(.A1(KEYINPUT80), .A2(new_n223), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n220), .A2(new_n222), .B1(KEYINPUT2), .B2(new_n205), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT80), .B1(new_n230), .B2(new_n227), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n210), .B(new_n214), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT84), .B1(new_n232), .B2(KEYINPUT4), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(KEYINPUT4), .B2(new_n232), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n230), .A2(KEYINPUT80), .A3(new_n227), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n209), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n239), .A2(KEYINPUT84), .A3(new_n240), .A4(new_n214), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n214), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n239), .B2(new_n243), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n210), .B1(new_n229), .B2(new_n231), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR4_X1   g052(.A1(new_n242), .A2(new_n251), .A3(KEYINPUT5), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n248), .A2(new_n250), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n214), .B1(new_n239), .B2(new_n243), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT82), .B1(new_n232), .B2(KEYINPUT4), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n232), .A2(KEYINPUT4), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n232), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT83), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT5), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n245), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n232), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n266), .B2(new_n253), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n257), .A2(new_n262), .A3(KEYINPUT83), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n254), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n272));
  XNOR2_X1  g071(.A(G1gat), .B(G29gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT0), .ZN(new_n274));
  XNOR2_X1  g073(.A(G57gat), .B(G85gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  NOR3_X1   g075(.A1(new_n271), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n270), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n278), .A2(new_n263), .A3(new_n268), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT89), .B1(new_n279), .B2(new_n254), .ZN(new_n280));
  INV_X1    g079(.A(new_n276), .ZN(new_n281));
  INV_X1    g080(.A(new_n263), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n270), .A3(new_n267), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT89), .ZN(new_n284));
  INV_X1    g083(.A(new_n254), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT6), .B1(new_n271), .B2(new_n276), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n277), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT25), .B1(new_n294), .B2(KEYINPUT66), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n296), .B(KEYINPUT64), .Z(new_n297));
  AOI21_X1  g096(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n298), .A2(KEYINPUT65), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n297), .B(new_n301), .C1(KEYINPUT65), .C2(new_n298), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n295), .B(new_n302), .C1(KEYINPUT66), .C2(new_n294), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n293), .B(KEYINPUT67), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n292), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT25), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n290), .A2(KEYINPUT70), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n311), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(KEYINPUT26), .B2(new_n311), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT27), .B(G183gat), .Z(new_n314));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n314), .A2(new_n315), .A3(G190gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  AOI21_X1  g117(.A(G190gat), .B1(new_n318), .B2(KEYINPUT27), .ZN(new_n319));
  OR3_X1    g118(.A1(new_n299), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT28), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI221_X1 g120(.A(new_n313), .B1(new_n299), .B2(new_n300), .C1(new_n316), .C2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n310), .A3(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n323), .A2(G226gat), .A3(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n323), .A2(new_n325), .B1(G226gat), .B2(G233gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT74), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT74), .B1(new_n328), .B2(new_n329), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G211gat), .B(G218gat), .Z(new_n334));
  OR3_X1    g133(.A1(new_n333), .A2(KEYINPUT75), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n333), .B2(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OR3_X1    g137(.A1(new_n324), .A2(new_n326), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n324), .B2(new_n326), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G8gat), .B(G36gat), .Z(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT76), .ZN(new_n343));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT30), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n346), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT90), .B1(new_n289), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351));
  INV_X1    g150(.A(new_n349), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n283), .A2(new_n276), .A3(new_n285), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n272), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n283), .A2(new_n285), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n276), .B1(new_n355), .B2(KEYINPUT89), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n356), .B2(new_n286), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n351), .B(new_n352), .C1(new_n357), .C2(new_n277), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n323), .A2(new_n245), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n303), .A2(new_n214), .A3(new_n310), .A4(new_n322), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT34), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT34), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n359), .A2(new_n365), .A3(new_n362), .A4(new_n360), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n362), .B1(new_n359), .B2(new_n360), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT32), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n369), .A2(KEYINPUT33), .ZN(new_n372));
  XOR2_X1   g171(.A(G15gat), .B(G43gat), .Z(new_n373));
  XNOR2_X1  g172(.A(G71gat), .B(G99gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n377));
  AOI221_X4 g176(.A(new_n377), .B1(KEYINPUT33), .B2(new_n375), .C1(new_n361), .C2(new_n363), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n368), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n375), .B1(new_n369), .B2(KEYINPUT33), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n369), .A2(new_n377), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n384), .A2(new_n378), .A3(new_n367), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(KEYINPUT91), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT91), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n380), .B2(new_n385), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT31), .B(G50gat), .ZN(new_n392));
  INV_X1    g191(.A(G106gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n338), .B1(new_n244), .B2(new_n325), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT86), .B1(new_n337), .B2(KEYINPUT29), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n335), .A2(new_n399), .A3(new_n325), .A4(new_n336), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n243), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n249), .ZN(new_n402));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n403), .B(KEYINPUT85), .Z(new_n407));
  INV_X1    g206(.A(new_n333), .ZN(new_n408));
  INV_X1    g207(.A(new_n334), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n409), .B2(new_n408), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n239), .B1(new_n243), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n407), .B1(new_n396), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(new_n406), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n406), .B1(new_n405), .B2(new_n413), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n415), .A2(G78gat), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G78gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n405), .A2(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n420), .B2(new_n414), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n395), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(G78gat), .B1(new_n415), .B2(new_n416), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n418), .A3(new_n414), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n394), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n391), .A2(KEYINPUT35), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n350), .A2(new_n358), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT71), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n364), .A2(new_n429), .A3(new_n366), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n364), .B2(new_n366), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n430), .A2(new_n431), .B1(new_n384), .B2(new_n378), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n376), .A2(new_n379), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n364), .A2(new_n429), .A3(new_n366), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n439), .A3(new_n386), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n426), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n281), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n271), .A2(new_n276), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n354), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n352), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT35), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n281), .B1(new_n271), .B2(new_n284), .ZN(new_n448));
  INV_X1    g247(.A(new_n286), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n288), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT37), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n339), .A2(new_n451), .A3(new_n340), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n339), .B2(new_n340), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n345), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT38), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n456), .B(new_n345), .C1(new_n452), .C2(new_n453), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n455), .A2(new_n348), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n443), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n426), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n253), .B1(new_n242), .B2(new_n251), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(KEYINPUT39), .C1(new_n253), .C2(new_n266), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n463), .B(new_n253), .C1(new_n242), .C2(new_n251), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(new_n465), .A3(new_n276), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n464), .B2(new_n276), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n468), .A2(KEYINPUT88), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT88), .B1(new_n468), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n287), .B(new_n349), .C1(new_n469), .C2(new_n468), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n459), .B(new_n460), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n380), .B2(new_n385), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT73), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n433), .A2(new_n439), .A3(KEYINPUT36), .A4(new_n386), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT73), .B(new_n475), .C1(new_n380), .C2(new_n385), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n446), .B2(new_n426), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n428), .A2(new_n447), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G43gat), .ZN(new_n485));
  INV_X1    g284(.A(G50gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G43gat), .A2(G50gat), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT94), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT15), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(KEYINPUT94), .A3(new_n488), .ZN(new_n492));
  INV_X1    g291(.A(G29gat), .ZN(new_n493));
  INV_X1    g292(.A(G36gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT14), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT95), .ZN(new_n498));
  NAND2_X1  g297(.A1(G29gat), .A2(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT95), .B1(new_n495), .B2(new_n497), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n491), .B(new_n492), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT96), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT95), .ZN(new_n505));
  INV_X1    g304(.A(new_n495), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT14), .B1(new_n493), .B2(new_n494), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n499), .A3(new_n498), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n509), .A2(KEYINPUT96), .A3(new_n492), .A4(new_n491), .ZN(new_n510));
  OR2_X1    g309(.A1(KEYINPUT97), .A2(KEYINPUT15), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT97), .A2(KEYINPUT15), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n511), .A2(new_n487), .A3(new_n488), .A4(new_n512), .ZN(new_n513));
  AND4_X1   g312(.A1(new_n497), .A2(new_n513), .A3(new_n495), .A4(new_n499), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n491), .A2(new_n492), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n504), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT17), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT8), .ZN(new_n521));
  OR2_X1    g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT102), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT102), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n526), .B2(new_n528), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n524), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n525), .A2(KEYINPUT102), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n535), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(new_n524), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n544), .A3(KEYINPUT103), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT103), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n543), .B1(new_n542), .B2(new_n524), .ZN(new_n547));
  AOI211_X1 g346(.A(new_n535), .B(new_n523), .C1(new_n540), .C2(new_n541), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n502), .A2(new_n503), .B1(new_n514), .B2(new_n515), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT17), .A3(new_n510), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n519), .A2(new_n545), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT41), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n545), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(new_n517), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(KEYINPUT104), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT104), .ZN(new_n559));
  AOI211_X1 g358(.A(new_n559), .B(new_n555), .C1(new_n556), .C2(new_n517), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n552), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G190gat), .B(G218gat), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(new_n554), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT101), .Z(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n562), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n568), .B(new_n552), .C1(new_n558), .C2(new_n560), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n563), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n567), .B1(new_n563), .B2(new_n569), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G57gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G64gat), .ZN(new_n575));
  INV_X1    g374(.A(G64gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G57gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT9), .ZN(new_n579));
  INV_X1    g378(.A(G71gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n418), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G71gat), .B(G78gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n578), .A2(new_n583), .A3(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  XNOR2_X1  g390(.A(G15gat), .B(G22gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT16), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(G1gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(KEYINPUT98), .C1(G1gat), .C2(new_n592), .ZN(new_n595));
  INV_X1    g394(.A(G8gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n588), .B2(new_n587), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n591), .B(new_n598), .Z(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT100), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT99), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n599), .B(new_n606), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n573), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n556), .A2(KEYINPUT10), .A3(new_n585), .A4(new_n586), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT105), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n578), .A2(new_n583), .A3(new_n581), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n583), .B1(new_n581), .B2(new_n578), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n585), .A2(KEYINPUT105), .A3(new_n586), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n614), .B(new_n615), .C1(new_n547), .C2(new_n548), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n536), .A2(new_n544), .A3(new_n587), .A4(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT106), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT106), .ZN(new_n621));
  AOI211_X1 g420(.A(new_n621), .B(KEYINPUT10), .C1(new_n616), .C2(new_n617), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n610), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n616), .A2(new_n626), .A3(new_n617), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n625), .A2(new_n627), .A3(new_n631), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n595), .B(G8gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n517), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n597), .B1(new_n517), .B2(new_n518), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT17), .B1(new_n550), .B2(new_n510), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n636), .B(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT18), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n519), .A2(new_n597), .A3(new_n551), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n644), .A2(KEYINPUT18), .A3(new_n636), .A4(new_n638), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n636), .B(KEYINPUT13), .Z(new_n646));
  INV_X1    g445(.A(new_n638), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n517), .A2(new_n637), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n643), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G113gat), .B(G141gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G169gat), .B(G197gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT93), .B(KEYINPUT12), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n643), .A2(new_n657), .A3(new_n645), .A4(new_n649), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n609), .A2(new_n635), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n484), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n445), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n349), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n669), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(G8gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(G1325gat));
  OR3_X1    g476(.A1(new_n664), .A2(G15gat), .A3(new_n391), .ZN(new_n678));
  INV_X1    g477(.A(new_n481), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n664), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(G1326gat));
  OR3_X1    g480(.A1(new_n664), .A2(KEYINPUT108), .A3(new_n460), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT108), .B1(new_n664), .B2(new_n460), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n428), .A2(new_n447), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n474), .A2(new_n482), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n573), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n608), .A2(new_n662), .A3(new_n635), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n493), .A3(new_n666), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n483), .B2(new_n573), .ZN(new_n697));
  AND4_X1   g496(.A1(new_n666), .A2(new_n695), .A3(new_n697), .A4(new_n690), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n694), .B1(new_n493), .B2(new_n698), .ZN(G1328gat));
  NOR3_X1   g498(.A1(new_n691), .A2(G36gat), .A3(new_n352), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  AND4_X1   g502(.A1(new_n349), .A2(new_n695), .A3(new_n697), .A4(new_n690), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n702), .B(new_n703), .C1(new_n494), .C2(new_n704), .ZN(G1329gat));
  OAI21_X1  g504(.A(new_n485), .B1(new_n691), .B2(new_n391), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n679), .A2(new_n485), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n695), .A2(new_n697), .A3(new_n690), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n710), .B(new_n711), .Z(G1330gat));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n691), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n426), .B1(new_n691), .B2(new_n713), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n486), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n460), .A2(new_n486), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n695), .A2(new_n697), .A3(new_n690), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT48), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n717), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1331gat));
  INV_X1    g523(.A(new_n635), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n609), .A2(new_n725), .A3(new_n661), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n484), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n445), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n574), .ZN(G1332gat));
  NOR2_X1   g528(.A1(new_n727), .A2(new_n352), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n727), .B2(new_n679), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n390), .A2(new_n580), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n727), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1334gat));
  NOR2_X1   g538(.A1(new_n727), .A2(new_n460), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n418), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n608), .A2(new_n661), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n725), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n695), .A2(new_n697), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n445), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n689), .B2(new_n742), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NOR4_X1   g547(.A1(new_n483), .A2(new_n748), .A3(new_n573), .A4(new_n743), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(G85gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n666), .A2(new_n751), .A3(new_n635), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n746), .B1(new_n750), .B2(new_n752), .ZN(G1336gat));
  NAND4_X1  g552(.A1(new_n695), .A2(new_n697), .A3(new_n349), .A4(new_n744), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n352), .A2(G92gat), .A3(new_n725), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n747), .B2(new_n749), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n745), .B2(new_n679), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n391), .A2(G99gat), .A3(new_n725), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT112), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n750), .B2(new_n762), .ZN(G1338gat));
  NOR3_X1   g562(.A1(new_n460), .A2(G106gat), .A3(new_n725), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n747), .B2(new_n749), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n695), .A2(new_n697), .A3(new_n426), .A4(new_n744), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n769), .A3(G106gat), .ZN(new_n770));
  OAI211_X1 g569(.A(KEYINPUT114), .B(new_n764), .C1(new_n747), .C2(new_n749), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT53), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(G106gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(KEYINPUT53), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n774), .B(new_n775), .C1(new_n765), .C2(KEYINPUT53), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(G1339gat));
  NAND4_X1  g576(.A1(new_n573), .A2(new_n608), .A3(new_n725), .A4(new_n662), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n626), .B(new_n610), .C1(new_n620), .C2(new_n622), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n625), .A2(KEYINPUT54), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n623), .A2(new_n782), .A3(new_n624), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n781), .A2(KEYINPUT55), .A3(new_n632), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n634), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT115), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n787), .A3(new_n634), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n781), .A2(new_n632), .A3(new_n783), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n636), .B1(new_n644), .B2(new_n638), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n647), .A2(new_n648), .A3(new_n646), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n655), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n660), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n570), .A2(new_n571), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n786), .A2(new_n788), .A3(new_n791), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT116), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n785), .A2(KEYINPUT115), .B1(new_n790), .B2(new_n789), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n788), .A4(new_n796), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n661), .A3(new_n788), .A4(new_n791), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n635), .A2(new_n660), .A3(new_n794), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n798), .B(new_n801), .C1(new_n804), .C2(new_n572), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n779), .B1(new_n805), .B2(new_n607), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n666), .A2(new_n352), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n391), .A2(new_n426), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(G113gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n810), .A2(new_n811), .A3(new_n662), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n798), .A2(new_n801), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n572), .B1(new_n802), .B2(new_n803), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n607), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n778), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n666), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n349), .A3(new_n442), .ZN(new_n818));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n661), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n812), .A2(new_n819), .ZN(G1340gat));
  INV_X1    g619(.A(G120gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n810), .A2(new_n821), .A3(new_n725), .ZN(new_n822));
  AOI21_X1  g621(.A(G120gat), .B1(new_n818), .B2(new_n635), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(G1341gat));
  OAI21_X1  g623(.A(G127gat), .B1(new_n810), .B2(new_n607), .ZN(new_n825));
  INV_X1    g624(.A(G127gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n818), .A2(new_n826), .A3(new_n608), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1342gat));
  INV_X1    g627(.A(new_n817), .ZN(new_n829));
  INV_X1    g628(.A(G134gat), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n349), .A2(new_n573), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n829), .A2(new_n830), .A3(new_n441), .A4(new_n831), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n810), .B2(new_n573), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G1343gat));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n807), .A2(new_n481), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n839), .B(new_n840), .C1(new_n806), .C2(new_n460), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n460), .B1(new_n815), .B2(new_n778), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT117), .B1(new_n842), .B2(KEYINPUT57), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n460), .A2(new_n840), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n791), .A2(new_n661), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n803), .B1(new_n846), .B2(new_n785), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n573), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n798), .A2(new_n848), .A3(new_n801), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n850), .A3(new_n607), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n778), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n849), .B2(new_n607), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n844), .B(new_n845), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n841), .A2(new_n843), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n853), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n778), .A3(new_n851), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n844), .B1(new_n857), .B2(new_n845), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n661), .B(new_n838), .C1(new_n855), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G141gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n481), .A2(new_n460), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n662), .A2(G141gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n808), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n837), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT121), .B(new_n865), .C1(new_n859), .C2(G141gat), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n863), .B(KEYINPUT120), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(G141gat), .B2(new_n859), .ZN(new_n870));
  OAI22_X1  g669(.A1(new_n867), .A2(new_n868), .B1(new_n864), .B2(new_n870), .ZN(G1344gat));
  AND2_X1   g670(.A1(new_n808), .A2(new_n861), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n221), .A3(new_n635), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n838), .B1(new_n855), .B2(new_n858), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n725), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(KEYINPUT59), .A3(new_n221), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  INV_X1    g676(.A(new_n842), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n778), .B(KEYINPUT122), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n608), .B1(new_n848), .B2(new_n797), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n840), .B(new_n426), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n879), .A2(new_n635), .A3(new_n838), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n873), .B1(new_n876), .B2(new_n884), .ZN(G1345gat));
  NOR3_X1   g684(.A1(new_n874), .A2(new_n202), .A3(new_n607), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n872), .A2(new_n608), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(KEYINPUT123), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(G155gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(KEYINPUT123), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1346gat));
  OAI211_X1 g690(.A(new_n572), .B(new_n838), .C1(new_n855), .C2(new_n858), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G162gat), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n829), .A2(new_n203), .A3(new_n831), .A4(new_n861), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(KEYINPUT124), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n666), .A2(new_n352), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n816), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(new_n441), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n661), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n809), .ZN(new_n904));
  INV_X1    g703(.A(G169gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(new_n662), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n906), .ZN(G1348gat));
  INV_X1    g706(.A(G176gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n902), .A2(new_n908), .A3(new_n635), .ZN(new_n909));
  OAI21_X1  g708(.A(G176gat), .B1(new_n904), .B2(new_n725), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1349gat));
  NOR2_X1   g710(.A1(new_n607), .A2(new_n314), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n901), .A2(new_n809), .A3(new_n608), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n902), .A2(new_n912), .B1(new_n913), .B2(G183gat), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g714(.A1(new_n902), .A2(new_n300), .A3(new_n572), .ZN(new_n916));
  OAI21_X1  g715(.A(G190gat), .B1(new_n904), .B2(new_n573), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n917), .A2(KEYINPUT61), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(KEYINPUT61), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n922), .B(new_n916), .C1(new_n918), .C2(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1351gat));
  AND3_X1   g723(.A1(new_n842), .A2(new_n679), .A3(new_n900), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n662), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n879), .A2(new_n679), .A3(new_n882), .A4(new_n900), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n661), .A2(G197gat), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n927), .A2(G197gat), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(G1352gat));
  NOR3_X1   g730(.A1(new_n926), .A2(G204gat), .A3(new_n725), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  OAI21_X1  g732(.A(G204gat), .B1(new_n928), .B2(new_n725), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1353gat));
  OAI21_X1  g734(.A(G211gat), .B1(new_n928), .B2(new_n607), .ZN(new_n936));
  NOR2_X1   g735(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI221_X1 g737(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .C1(new_n928), .C2(new_n607), .ZN(new_n939));
  NAND2_X1  g738(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n607), .A2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n926), .B2(new_n942), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n928), .B2(new_n573), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n573), .A2(G218gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n926), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


