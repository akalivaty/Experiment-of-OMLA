

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576;

  XNOR2_X1 U320 ( .A(KEYINPUT48), .B(n379), .ZN(n509) );
  NOR2_X1 U321 ( .A1(n574), .A2(n468), .ZN(n354) );
  NOR2_X1 U322 ( .A1(n542), .A2(n371), .ZN(n372) );
  NOR2_X2 U323 ( .A1(n512), .A2(n288), .ZN(n545) );
  XNOR2_X1 U324 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U325 ( .A(n390), .B(n305), .Z(n503) );
  XOR2_X1 U326 ( .A(KEYINPUT55), .B(n436), .Z(n288) );
  XOR2_X1 U327 ( .A(n369), .B(G127GAT), .Z(n289) );
  INV_X1 U328 ( .A(G106GAT), .ZN(n364) );
  XNOR2_X1 U329 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U330 ( .A(n347), .B(G71GAT), .ZN(n348) );
  XNOR2_X1 U331 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U332 ( .A(n565), .B(KEYINPUT41), .Z(n544) );
  XOR2_X1 U333 ( .A(n353), .B(n352), .Z(n570) );
  XOR2_X1 U334 ( .A(KEYINPUT28), .B(n448), .Z(n515) );
  XNOR2_X1 U335 ( .A(n437), .B(G190GAT), .ZN(n438) );
  XNOR2_X1 U336 ( .A(n439), .B(n438), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT19), .B(KEYINPUT79), .Z(n291) );
  XNOR2_X1 U338 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U340 ( .A(n292), .B(G183GAT), .Z(n294) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G176GAT), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n390) );
  XOR2_X1 U343 ( .A(G120GAT), .B(G71GAT), .Z(n363) );
  XOR2_X1 U344 ( .A(G99GAT), .B(G190GAT), .Z(n296) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G15GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U347 ( .A(n363), .B(n297), .Z(n299) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n302) );
  XOR2_X1 U350 ( .A(G127GAT), .B(KEYINPUT0), .Z(n301) );
  XNOR2_X1 U351 ( .A(G113GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n415) );
  XOR2_X1 U353 ( .A(n302), .B(n415), .Z(n304) );
  XNOR2_X1 U354 ( .A(KEYINPUT20), .B(KEYINPUT80), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n305) );
  INV_X1 U356 ( .A(n503), .ZN(n512) );
  XOR2_X1 U357 ( .A(G141GAT), .B(G197GAT), .Z(n307) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(G113GAT), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U360 ( .A(KEYINPUT66), .B(n308), .Z(n310) );
  NAND2_X1 U361 ( .A1(G229GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U363 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U366 ( .A(n314), .B(n313), .Z(n323) );
  XNOR2_X1 U367 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n315), .B(G29GAT), .ZN(n316) );
  XOR2_X1 U369 ( .A(n316), .B(KEYINPUT8), .Z(n318) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G50GAT), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n327) );
  XOR2_X1 U372 ( .A(G22GAT), .B(G15GAT), .Z(n320) );
  XNOR2_X1 U373 ( .A(KEYINPUT68), .B(G1GAT), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U375 ( .A(G8GAT), .B(n321), .ZN(n352) );
  XOR2_X1 U376 ( .A(n327), .B(n352), .Z(n322) );
  XOR2_X1 U377 ( .A(n323), .B(n322), .Z(n482) );
  XOR2_X1 U378 ( .A(KEYINPUT70), .B(n482), .Z(n542) );
  XOR2_X1 U379 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n325) );
  XNOR2_X1 U380 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n336) );
  XNOR2_X1 U383 ( .A(G99GAT), .B(G92GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n328), .B(G85GAT), .ZN(n360) );
  XOR2_X1 U385 ( .A(G162GAT), .B(G106GAT), .Z(n424) );
  XNOR2_X1 U386 ( .A(n360), .B(n424), .ZN(n330) );
  AND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(n331), .B(KEYINPUT65), .Z(n334) );
  XNOR2_X1 U390 ( .A(G190GAT), .B(G218GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n332), .B(KEYINPUT72), .ZN(n380) );
  XNOR2_X1 U392 ( .A(n380), .B(KEYINPUT10), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n539) );
  XNOR2_X1 U395 ( .A(KEYINPUT73), .B(n539), .ZN(n527) );
  XNOR2_X1 U396 ( .A(KEYINPUT36), .B(n527), .ZN(n574) );
  XOR2_X1 U397 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n338) );
  XNOR2_X1 U398 ( .A(KEYINPUT12), .B(KEYINPUT78), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n351) );
  XNOR2_X1 U400 ( .A(G64GAT), .B(G57GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(KEYINPUT13), .B(n339), .ZN(n369) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n289), .B(n340), .ZN(n349) );
  XOR2_X1 U404 ( .A(G155GAT), .B(G78GAT), .Z(n342) );
  XNOR2_X1 U405 ( .A(G183GAT), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U407 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n344) );
  XNOR2_X1 U408 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U410 ( .A(n346), .B(n345), .Z(n347) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n353) );
  INV_X1 U412 ( .A(n570), .ZN(n468) );
  XNOR2_X1 U413 ( .A(KEYINPUT45), .B(n354), .ZN(n370) );
  XOR2_X1 U414 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n356) );
  NAND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U417 ( .A(n357), .B(KEYINPUT33), .Z(n362) );
  XOR2_X1 U418 ( .A(G78GAT), .B(G148GAT), .Z(n359) );
  XNOR2_X1 U419 ( .A(KEYINPUT71), .B(G204GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n430) );
  XNOR2_X1 U421 ( .A(n430), .B(n360), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n367) );
  XNOR2_X1 U423 ( .A(G176GAT), .B(n363), .ZN(n365) );
  XOR2_X1 U424 ( .A(n369), .B(n368), .Z(n458) );
  NAND2_X1 U425 ( .A1(n370), .A2(n458), .ZN(n371) );
  XNOR2_X1 U426 ( .A(KEYINPUT107), .B(n372), .ZN(n378) );
  INV_X1 U427 ( .A(n482), .ZN(n562) );
  INV_X1 U428 ( .A(n458), .ZN(n565) );
  NAND2_X1 U429 ( .A1(n562), .A2(n544), .ZN(n373) );
  XNOR2_X1 U430 ( .A(KEYINPUT46), .B(n373), .ZN(n374) );
  XOR2_X1 U431 ( .A(KEYINPUT106), .B(n570), .Z(n551) );
  NAND2_X1 U432 ( .A1(n374), .A2(n551), .ZN(n375) );
  NOR2_X1 U433 ( .A1(n375), .A2(n539), .ZN(n376) );
  XNOR2_X1 U434 ( .A(KEYINPUT47), .B(n376), .ZN(n377) );
  NAND2_X1 U435 ( .A1(n378), .A2(n377), .ZN(n379) );
  XOR2_X1 U436 ( .A(G92GAT), .B(KEYINPUT92), .Z(n382) );
  XNOR2_X1 U437 ( .A(G36GAT), .B(n380), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U439 ( .A(KEYINPUT91), .B(G64GAT), .Z(n384) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U442 ( .A(n386), .B(n385), .Z(n388) );
  XNOR2_X1 U443 ( .A(G8GAT), .B(G204GAT), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n395) );
  XOR2_X1 U446 ( .A(KEYINPUT84), .B(G211GAT), .Z(n392) );
  XNOR2_X1 U447 ( .A(G197GAT), .B(KEYINPUT82), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U449 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n393) );
  XOR2_X1 U450 ( .A(n394), .B(n393), .Z(n429) );
  XOR2_X1 U451 ( .A(n395), .B(n429), .Z(n500) );
  NAND2_X1 U452 ( .A1(n509), .A2(n500), .ZN(n397) );
  XOR2_X1 U453 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n418) );
  XOR2_X1 U455 ( .A(G85GAT), .B(G162GAT), .Z(n399) );
  XNOR2_X1 U456 ( .A(G29GAT), .B(G120GAT), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U458 ( .A(KEYINPUT89), .B(G57GAT), .Z(n401) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(G148GAT), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U461 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n405) );
  NAND2_X1 U463 ( .A1(G225GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U465 ( .A(KEYINPUT1), .B(n406), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U467 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n410) );
  XNOR2_X1 U468 ( .A(KEYINPUT90), .B(KEYINPUT6), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U470 ( .A(n412), .B(n411), .Z(n417) );
  XOR2_X1 U471 ( .A(G155GAT), .B(KEYINPUT2), .Z(n414) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n427) );
  XNOR2_X1 U474 ( .A(n415), .B(n427), .ZN(n416) );
  XOR2_X1 U475 ( .A(n417), .B(n416), .Z(n442) );
  INV_X1 U476 ( .A(n442), .ZN(n496) );
  NOR2_X2 U477 ( .A1(n418), .A2(n496), .ZN(n559) );
  XOR2_X1 U478 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n420) );
  XNOR2_X1 U479 ( .A(KEYINPUT85), .B(KEYINPUT23), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n420), .B(n419), .ZN(n435) );
  XOR2_X1 U481 ( .A(KEYINPUT22), .B(G218GAT), .Z(n422) );
  XNOR2_X1 U482 ( .A(G50GAT), .B(G22GAT), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U484 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U487 ( .A(n428), .B(n427), .Z(n433) );
  INV_X1 U488 ( .A(n429), .ZN(n431) );
  XOR2_X1 U489 ( .A(n431), .B(n430), .Z(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n448) );
  NAND2_X1 U492 ( .A1(n559), .A2(n448), .ZN(n436) );
  INV_X1 U493 ( .A(n545), .ZN(n550) );
  NOR2_X1 U494 ( .A1(n550), .A2(n527), .ZN(n439) );
  XNOR2_X1 U495 ( .A(KEYINPUT119), .B(KEYINPUT58), .ZN(n437) );
  NAND2_X1 U496 ( .A1(n570), .A2(n527), .ZN(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT16), .B(n440), .Z(n457) );
  XOR2_X1 U498 ( .A(n512), .B(KEYINPUT81), .Z(n443) );
  XNOR2_X1 U499 ( .A(KEYINPUT27), .B(KEYINPUT93), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n441), .B(n500), .ZN(n450) );
  NOR2_X1 U501 ( .A1(n442), .A2(n450), .ZN(n510) );
  NAND2_X1 U502 ( .A1(n443), .A2(n510), .ZN(n444) );
  NOR2_X1 U503 ( .A1(n515), .A2(n444), .ZN(n445) );
  XOR2_X1 U504 ( .A(KEYINPUT94), .B(n445), .Z(n456) );
  NAND2_X1 U505 ( .A1(n503), .A2(n500), .ZN(n446) );
  NAND2_X1 U506 ( .A1(n448), .A2(n446), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n447), .B(KEYINPUT25), .ZN(n452) );
  NOR2_X1 U508 ( .A1(n503), .A2(n448), .ZN(n449) );
  XOR2_X1 U509 ( .A(KEYINPUT26), .B(n449), .Z(n558) );
  NOR2_X1 U510 ( .A1(n450), .A2(n558), .ZN(n451) );
  NOR2_X1 U511 ( .A1(n452), .A2(n451), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n496), .A2(n453), .ZN(n454) );
  XNOR2_X1 U513 ( .A(KEYINPUT95), .B(n454), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n456), .A2(n455), .ZN(n467) );
  NAND2_X1 U515 ( .A1(n457), .A2(n467), .ZN(n483) );
  NAND2_X1 U516 ( .A1(n458), .A2(n542), .ZN(n471) );
  NOR2_X1 U517 ( .A1(n483), .A2(n471), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT96), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n465), .A2(n496), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT34), .ZN(n461) );
  XNOR2_X1 U521 ( .A(G1GAT), .B(n461), .ZN(G1324GAT) );
  NAND2_X1 U522 ( .A1(n465), .A2(n500), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n462), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U524 ( .A(G15GAT), .B(KEYINPUT35), .Z(n464) );
  NAND2_X1 U525 ( .A1(n503), .A2(n465), .ZN(n463) );
  XNOR2_X1 U526 ( .A(n464), .B(n463), .ZN(G1326GAT) );
  NAND2_X1 U527 ( .A1(n465), .A2(n515), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U529 ( .A(KEYINPUT97), .B(KEYINPUT39), .Z(n474) );
  NAND2_X1 U530 ( .A1(n468), .A2(n467), .ZN(n469) );
  NOR2_X1 U531 ( .A1(n574), .A2(n469), .ZN(n470) );
  XNOR2_X1 U532 ( .A(KEYINPUT37), .B(n470), .ZN(n495) );
  NOR2_X1 U533 ( .A1(n471), .A2(n495), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n472), .B(KEYINPUT38), .ZN(n480) );
  NAND2_X1 U535 ( .A1(n496), .A2(n480), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U537 ( .A(G29GAT), .B(n475), .Z(G1328GAT) );
  NAND2_X1 U538 ( .A1(n480), .A2(n500), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT40), .B(KEYINPUT98), .Z(n478) );
  NAND2_X1 U541 ( .A1(n503), .A2(n480), .ZN(n477) );
  XNOR2_X1 U542 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U543 ( .A(G43GAT), .B(n479), .Z(G1330GAT) );
  NAND2_X1 U544 ( .A1(n480), .A2(n515), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n481), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT99), .B(KEYINPUT42), .Z(n485) );
  NAND2_X1 U547 ( .A1(n482), .A2(n544), .ZN(n494) );
  NOR2_X1 U548 ( .A1(n483), .A2(n494), .ZN(n490) );
  NAND2_X1 U549 ( .A1(n490), .A2(n496), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U551 ( .A(G57GAT), .B(n486), .ZN(G1332GAT) );
  NAND2_X1 U552 ( .A1(n500), .A2(n490), .ZN(n487) );
  XNOR2_X1 U553 ( .A(n487), .B(KEYINPUT100), .ZN(n488) );
  XNOR2_X1 U554 ( .A(G64GAT), .B(n488), .ZN(G1333GAT) );
  NAND2_X1 U555 ( .A1(n490), .A2(n503), .ZN(n489) );
  XNOR2_X1 U556 ( .A(n489), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT43), .B(KEYINPUT101), .Z(n492) );
  NAND2_X1 U558 ( .A1(n490), .A2(n515), .ZN(n491) );
  XNOR2_X1 U559 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U560 ( .A(G78GAT), .B(n493), .Z(G1335GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n498) );
  NOR2_X1 U562 ( .A1(n495), .A2(n494), .ZN(n505) );
  NAND2_X1 U563 ( .A1(n505), .A2(n496), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U565 ( .A(G85GAT), .B(n499), .ZN(G1336GAT) );
  NAND2_X1 U566 ( .A1(n500), .A2(n505), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n501), .B(KEYINPUT104), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G92GAT), .B(n502), .ZN(G1337GAT) );
  NAND2_X1 U569 ( .A1(n505), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n507) );
  NAND2_X1 U572 ( .A1(n505), .A2(n515), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G106GAT), .B(n508), .ZN(G1339GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(KEYINPUT108), .ZN(n531) );
  NOR2_X1 U577 ( .A1(n531), .A2(n512), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT109), .ZN(n514) );
  NOR2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n542), .A2(n523), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT110), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G113GAT), .B(n517), .ZN(G1340GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n519) );
  NAND2_X1 U584 ( .A1(n523), .A2(n544), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(G120GAT), .B(n520), .Z(G1341GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n522) );
  XNOR2_X1 U588 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n525) );
  INV_X1 U590 ( .A(n523), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n551), .A2(n526), .ZN(n524) );
  XOR2_X1 U592 ( .A(n525), .B(n524), .Z(G1342GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U594 ( .A(KEYINPUT51), .B(KEYINPUT114), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G134GAT), .B(n530), .ZN(G1343GAT) );
  NOR2_X1 U597 ( .A1(n531), .A2(n558), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n562), .A2(n540), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G141GAT), .B(n532), .ZN(G1344GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT53), .Z(n534) );
  NAND2_X1 U601 ( .A1(n540), .A2(n544), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U603 ( .A(G148GAT), .B(KEYINPUT52), .Z(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1345GAT) );
  NAND2_X1 U605 ( .A1(n540), .A2(n570), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n537), .B(KEYINPUT116), .ZN(n538) );
  XNOR2_X1 U607 ( .A(G155GAT), .B(n538), .ZN(G1346GAT) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n541), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U610 ( .A1(n542), .A2(n545), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n543), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U612 ( .A(G176GAT), .B(KEYINPUT118), .ZN(n549) );
  XOR2_X1 U613 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n547) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1349GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(G183GAT), .B(n552), .Z(G1350GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT121), .B(KEYINPUT123), .Z(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(n555), .B(KEYINPUT124), .Z(n557) );
  XNOR2_X1 U623 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n564) );
  INV_X1 U625 ( .A(n558), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT120), .B(n561), .ZN(n573) );
  INV_X1 U628 ( .A(n573), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n569), .A2(n562), .ZN(n563) );
  XOR2_X1 U630 ( .A(n564), .B(n563), .Z(G1352GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n567) );
  NAND2_X1 U632 ( .A1(n569), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G204GAT), .B(n568), .Z(G1353GAT) );
  XNOR2_X1 U635 ( .A(G211GAT), .B(KEYINPUT126), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1354GAT) );
  NOR2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT62), .B(n575), .Z(n576) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(n576), .ZN(G1355GAT) );
endmodule

