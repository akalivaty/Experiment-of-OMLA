//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n461), .B1(new_n477), .B2(new_n478), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n461), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n481), .A2(new_n486), .ZN(G162));
  AND2_X1   g062(.A1(KEYINPUT69), .A2(G114), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT69), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n482), .A2(G126), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n461), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n477), .B2(new_n478), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n493), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT70), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT70), .A2(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(KEYINPUT6), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT71), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n505), .A2(new_n512), .A3(KEYINPUT6), .A4(new_n506), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n504), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n511), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G88), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT70), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT70), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n516), .A2(new_n517), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT72), .Z(new_n528));
  OAI21_X1  g103(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n515), .A2(new_n520), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  XOR2_X1   g106(.A(KEYINPUT73), .B(G89), .Z(new_n532));
  NAND2_X1  g107(.A1(new_n519), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n509), .B1(new_n523), .B2(KEYINPUT6), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n535));
  NOR4_X1   g110(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT71), .A4(new_n535), .ZN(new_n536));
  OAI211_X1 g111(.A(G51), .B(G543), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n533), .A2(new_n537), .A3(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n519), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n514), .A2(G52), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n523), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  XOR2_X1   g124(.A(KEYINPUT74), .B(G43), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n514), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n519), .A2(G81), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n523), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT76), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  OAI211_X1 g137(.A(G53), .B(G543), .C1(new_n534), .C2(new_n536), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n514), .A2(new_n565), .A3(G53), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n516), .B2(new_n517), .ZN(new_n569));
  AND2_X1   g144(.A1(G78), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g148(.A(KEYINPUT77), .B(G651), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n573), .A2(new_n574), .B1(new_n519), .B2(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n567), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G74), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n508), .B1(new_n518), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n514), .B2(G49), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n519), .A2(KEYINPUT78), .A3(G87), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT78), .B1(new_n519), .B2(G87), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(G288));
  OAI211_X1 g157(.A(G86), .B(new_n525), .C1(new_n534), .C2(new_n536), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n518), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n514), .A2(G48), .B1(new_n524), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n519), .A2(G85), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(G543), .B1(new_n534), .B2(new_n536), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT80), .B(G47), .Z(new_n594));
  OAI221_X1 g169(.A(new_n591), .B1(new_n523), .B2(new_n592), .C1(new_n593), .C2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n519), .A2(G92), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT10), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n508), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n514), .A2(KEYINPUT81), .ZN(new_n601));
  OAI21_X1  g176(.A(G54), .B1(new_n514), .B2(KEYINPUT81), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n596), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n567), .A2(new_n575), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  OAI21_X1  g187(.A(KEYINPUT82), .B1(new_n555), .B2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n604), .A2(new_n611), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  MUX2_X1   g190(.A(KEYINPUT82), .B(new_n613), .S(new_n615), .Z(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n494), .A2(new_n466), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT84), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT13), .Z(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n479), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n482), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n461), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(new_n624), .A3(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT87), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT86), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(new_n637), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  AND2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(G14), .B1(new_n646), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(G401));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2096), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n665), .A2(new_n668), .A3(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT90), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(KEYINPUT104), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(G23), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G288), .B2(G16), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT33), .B(G1976), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(G22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT94), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G303), .B2(G16), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT95), .B(G1971), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n688), .A2(new_n689), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n690), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n686), .B1(new_n585), .B2(new_n589), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n686), .A2(G6), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n700), .A2(new_n701), .A3(new_n699), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT32), .B(G1981), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n697), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n706), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n703), .B2(new_n704), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n685), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n690), .A2(new_n695), .A3(new_n696), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n701), .B1(G305), .B2(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(new_n698), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(new_n706), .A3(new_n702), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n711), .A2(new_n709), .A3(new_n685), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n479), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n482), .A2(G119), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n461), .A2(G107), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT35), .B(G1991), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT91), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n721), .B(new_n723), .Z(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n686), .A2(G24), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G290), .B2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT36), .B1(new_n710), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n711), .A2(new_n714), .ZN(new_n732));
  INV_X1    g307(.A(new_n709), .ZN(new_n733));
  OAI21_X1  g308(.A(KEYINPUT34), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n734), .A2(new_n735), .A3(new_n715), .A4(new_n729), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n555), .A2(G16), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G16), .B2(G19), .ZN(new_n739));
  INV_X1    g314(.A(G1341), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n686), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n686), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G1966), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G32), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT26), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n750), .A2(new_n751), .B1(G105), .B2(new_n466), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n479), .A2(G141), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n482), .A2(G129), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n747), .B1(new_n756), .B2(new_n746), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G160), .A2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G34), .Z(new_n762));
  OAI21_X1  g337(.A(new_n760), .B1(G29), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n757), .A2(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n746), .A2(G27), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G164), .B2(new_n746), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G2078), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n765), .B(new_n768), .C1(new_n757), .C2(new_n759), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT31), .B(G11), .Z(new_n770));
  INV_X1    g345(.A(G28), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(KEYINPUT30), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT102), .Z(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n771), .B2(KEYINPUT30), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(new_n746), .B2(new_n629), .C1(new_n767), .C2(G2078), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n479), .A2(G139), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT97), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n494), .A2(G127), .ZN(new_n780));
  INV_X1    g355(.A(G115), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n465), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n783));
  NAND2_X1  g358(.A1(G103), .A2(G2104), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G2105), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n782), .A2(G2105), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n779), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n746), .A2(G33), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(G29), .B1(new_n481), .B2(new_n486), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n746), .A2(G35), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(KEYINPUT29), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT29), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n796), .A2(new_n800), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G2090), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n745), .A2(new_n777), .A3(new_n795), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G171), .A2(G16), .ZN(new_n805));
  OR2_X1    g380(.A1(G5), .A2(G16), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1961), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n479), .A2(G140), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n482), .A2(G128), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n461), .A2(G116), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n813), .A2(G29), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n746), .A2(G26), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT28), .Z(new_n816));
  OAI21_X1  g391(.A(KEYINPUT96), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G2067), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n814), .A2(KEYINPUT96), .A3(new_n816), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n820), .ZN(new_n822));
  AOI21_X1  g397(.A(G2067), .B1(new_n822), .B2(new_n817), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n763), .A2(new_n764), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT100), .Z(new_n826));
  AOI22_X1  g401(.A1(new_n739), .A2(new_n740), .B1(new_n743), .B2(G1966), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n808), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n804), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G2090), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n799), .A2(new_n830), .A3(new_n801), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(KEYINPUT101), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n686), .A2(G4), .ZN(new_n835));
  INV_X1    g410(.A(new_n604), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(G16), .ZN(new_n837));
  INV_X1    g412(.A(G1348), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n746), .B1(new_n789), .B2(new_n790), .ZN(new_n840));
  INV_X1    g415(.A(new_n794), .ZN(new_n841));
  OAI211_X1 g416(.A(KEYINPUT101), .B(G2072), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n834), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n837), .A2(new_n838), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n686), .A2(G20), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT23), .Z(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G299), .B2(G16), .ZN(new_n849));
  INV_X1    g424(.A(G1956), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n845), .A2(new_n846), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n829), .A2(new_n844), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n684), .B1(new_n737), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g430(.A(KEYINPUT104), .B(new_n853), .C1(new_n731), .C2(new_n736), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(G311));
  NAND2_X1  g432(.A1(new_n737), .A2(new_n854), .ZN(G150));
  NAND2_X1  g433(.A1(new_n514), .A2(G55), .ZN(new_n859));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  INV_X1    g435(.A(G67), .ZN(new_n861));
  OAI211_X1 g436(.A(KEYINPUT105), .B(new_n860), .C1(new_n518), .C2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n861), .B1(new_n516), .B2(new_n517), .ZN(new_n864));
  INV_X1    g439(.A(new_n860), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n524), .A3(new_n866), .ZN(new_n867));
  OAI211_X1 g442(.A(G93), .B(new_n525), .C1(new_n534), .C2(new_n536), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n859), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n604), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(KEYINPUT106), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n859), .A2(new_n867), .A3(new_n875), .A4(new_n868), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n555), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n555), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n873), .B(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n883));
  INV_X1    g458(.A(G860), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n882), .B2(KEYINPUT39), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n871), .B1(new_n883), .B2(new_n885), .ZN(G145));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n629), .B(G160), .Z(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(G162), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n813), .B(new_n502), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n756), .ZN(new_n891));
  INV_X1    g466(.A(new_n788), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n482), .A2(G130), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n461), .A2(G118), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(G142), .B2(new_n479), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n720), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n621), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n891), .A2(new_n790), .A3(new_n789), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n893), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n893), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n889), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(new_n889), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n903), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n903), .A2(new_n906), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n887), .B(new_n904), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  AND3_X1   g485(.A1(new_n874), .A2(new_n555), .A3(new_n876), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n555), .B1(new_n874), .B2(new_n876), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n614), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT10), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n597), .B(new_n915), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n601), .A2(new_n602), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n608), .A2(new_n916), .A3(new_n917), .A4(new_n600), .ZN(new_n918));
  OAI21_X1  g493(.A(G299), .B1(new_n598), .B2(new_n603), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n923), .A3(new_n919), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n918), .B2(new_n919), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n922), .B1(new_n927), .B2(new_n914), .ZN(new_n928));
  NOR2_X1   g503(.A1(KEYINPUT108), .A2(KEYINPUT42), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI221_X1 g505(.A(new_n922), .B1(KEYINPUT108), .B2(KEYINPUT42), .C1(new_n927), .C2(new_n914), .ZN(new_n931));
  XNOR2_X1  g506(.A(G305), .B(G290), .ZN(new_n932));
  XNOR2_X1  g507(.A(G288), .B(G303), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(KEYINPUT108), .B2(KEYINPUT42), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n930), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n930), .B2(new_n931), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G868), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n869), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(G295));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n940), .ZN(G331));
  AND2_X1   g517(.A1(G301), .A2(G286), .ZN(new_n943));
  NOR2_X1   g518(.A1(G301), .A2(G286), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n880), .A3(new_n879), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n911), .B2(new_n912), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n921), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n881), .B2(new_n945), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n945), .B(new_n950), .C1(new_n911), .C2(new_n912), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n947), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n920), .A2(KEYINPUT41), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n924), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n949), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n957), .B2(new_n934), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n920), .B1(new_n913), .B2(new_n946), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n948), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n948), .A2(KEYINPUT109), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n961), .A2(new_n952), .B1(new_n913), .B2(new_n946), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n962), .B2(new_n927), .ZN(new_n963));
  INV_X1    g538(.A(new_n934), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT43), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n960), .B(new_n934), .C1(new_n962), .C2(new_n927), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n887), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n955), .A2(new_n969), .A3(new_n924), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n947), .A2(new_n948), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n925), .A2(KEYINPUT110), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n959), .B1(new_n951), .B2(new_n953), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n934), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n968), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT44), .B1(new_n966), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n958), .B2(new_n965), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n968), .A2(new_n975), .A3(KEYINPUT43), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n982), .ZN(G397));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n984));
  INV_X1    g559(.A(G1981), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n583), .A2(new_n584), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT79), .B1(new_n519), .B2(G86), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n985), .B(new_n589), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(G288), .A2(G1976), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT116), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n588), .A2(new_n524), .ZN(new_n991));
  INV_X1    g566(.A(G48), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n593), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n583), .ZN(new_n994));
  OAI21_X1  g569(.A(G1981), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n988), .A2(KEYINPUT49), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT49), .B1(new_n988), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n988), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n493), .B2(new_n501), .ZN(new_n1001));
  INV_X1    g576(.A(G40), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n468), .A2(new_n473), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  INV_X1    g580(.A(G125), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n476), .A2(new_n465), .ZN(new_n1007));
  NAND2_X1  g582(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n472), .ZN(new_n1010));
  OAI21_X1  g585(.A(G2105), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1011), .A2(G40), .A3(new_n464), .A4(new_n467), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n495), .A2(G2105), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n462), .B2(new_n463), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1015), .A2(KEYINPUT4), .B1(new_n494), .B2(new_n496), .ZN(new_n1016));
  OAI211_X1 g591(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n1017));
  OR2_X1    g592(.A1(KEYINPUT69), .A2(G114), .ZN(new_n1018));
  NAND2_X1  g593(.A1(KEYINPUT69), .A2(G114), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n461), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1017), .B1(new_n1020), .B2(new_n491), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1013), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1012), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1001), .A2(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1023), .A2(new_n830), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1012), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT45), .B(new_n1013), .C1(new_n1016), .C2(new_n1021), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1971), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1005), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(G166), .B2(new_n1000), .ZN(new_n1033));
  NAND3_X1  g608(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1971), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1003), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1029), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1023), .A2(new_n830), .A3(new_n1025), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT115), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1031), .A2(new_n1035), .A3(new_n1041), .A4(G8), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1004), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n996), .A2(new_n997), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G288), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  OAI211_X1 g623(.A(G1976), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1004), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1004), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1045), .A2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n999), .A2(new_n1004), .B1(new_n1043), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1035), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT117), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT117), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1029), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1001), .A2(KEYINPUT118), .A3(KEYINPUT45), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1028), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1966), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1062), .A2(new_n764), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1068), .A2(new_n1000), .A3(G286), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1054), .A2(new_n1042), .A3(new_n1060), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT63), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1073));
  INV_X1    g648(.A(new_n997), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n988), .A2(new_n995), .A3(KEYINPUT49), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1004), .A3(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1042), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1023), .A2(new_n764), .A3(new_n1025), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1080), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1031), .A2(G8), .A3(new_n1041), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1056), .B2(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n984), .B(new_n1055), .C1(new_n1072), .C2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1070), .A2(new_n1071), .B1(new_n1077), .B2(new_n1083), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n999), .A2(new_n1004), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1054), .A2(new_n1043), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT119), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G286), .A2(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT125), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n1093));
  NAND3_X1  g668(.A1(G286), .A2(new_n1093), .A3(G8), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1080), .B2(G8), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT51), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G2078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1028), .A2(new_n1101), .A3(new_n1029), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  INV_X1    g678(.A(G1961), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1102), .A2(new_n1103), .B1(new_n1061), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(G2078), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1028), .A2(new_n1064), .A3(new_n1065), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G301), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1106), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1037), .A2(new_n1038), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1111), .B2(new_n1109), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1108), .A2(new_n1112), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1095), .A2(KEYINPUT126), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1117), .A2(KEYINPUT51), .B1(new_n1068), .B2(new_n1097), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1100), .B(new_n1116), .C1(new_n1096), .C2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1054), .A2(new_n1042), .A3(new_n1060), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1028), .A2(new_n1029), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(G1956), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n567), .A2(new_n575), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n567), .B2(new_n575), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1124), .A2(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1061), .A2(new_n850), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1126), .ZN(new_n1131));
  NAND2_X1  g706(.A1(G299), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n567), .A2(new_n575), .A3(new_n1126), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1130), .A2(new_n1132), .A3(new_n1123), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1129), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  OAI221_X1 g712(.A(KEYINPUT124), .B1(new_n1127), .B2(new_n1128), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(G2067), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1061), .B2(new_n838), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n836), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(KEYINPUT60), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  AOI21_X1  g720(.A(G1348), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(new_n1141), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1147), .A3(new_n604), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1132), .A2(new_n1150), .A3(new_n1133), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1149), .A2(new_n1151), .B1(new_n1130), .B2(new_n1123), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1134), .A2(KEYINPUT61), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1143), .B(new_n1148), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1155));
  INV_X1    g730(.A(G1996), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n1029), .A4(new_n1003), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT58), .B(G1341), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1140), .A2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1157), .A2(KEYINPUT123), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT123), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n555), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(KEYINPUT59), .B(new_n555), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1139), .A2(new_n1154), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1134), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n836), .A2(new_n1142), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1169), .A2(KEYINPUT121), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(new_n1152), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(KEYINPUT121), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1121), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1100), .B1(new_n1118), .B2(new_n1096), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1108), .A2(G171), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1120), .A2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1100), .B(KEYINPUT62), .C1(new_n1096), .C2(new_n1118), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1085), .A2(new_n1090), .A3(new_n1174), .A4(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1022), .A2(new_n1003), .A3(new_n1027), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT112), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n813), .B(new_n819), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1156), .B2(new_n756), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1183), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1156), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1187), .B1(new_n755), .B2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT113), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n720), .A2(new_n723), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n720), .A2(new_n723), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1184), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OR3_X1    g769(.A1(G290), .A2(G1986), .A3(new_n1183), .ZN(new_n1195));
  NAND3_X1  g770(.A1(G290), .A2(new_n1188), .A3(G1986), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT111), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1191), .A2(new_n1194), .A3(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT114), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1182), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1184), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n813), .A2(G2067), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g780(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1195), .B(new_n1206), .Z(new_n1207));
  AND3_X1   g782(.A1(new_n1191), .A2(new_n1194), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1202), .B1(new_n756), .B2(new_n1185), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1189), .B(KEYINPUT46), .Z(new_n1210));
  NOR2_X1   g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT47), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1205), .A2(new_n1208), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1201), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g789(.A1(new_n459), .A2(G227), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1216), .B1(new_n648), .B2(new_n649), .ZN(new_n1217));
  NOR2_X1   g791(.A1(G229), .A2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g792(.A(new_n909), .B(new_n1218), .C1(new_n980), .C2(new_n981), .ZN(G225));
  INV_X1    g793(.A(G225), .ZN(G308));
endmodule


