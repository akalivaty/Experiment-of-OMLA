//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n460), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n467), .B2(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n462), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n470), .B2(new_n471), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n465), .A2(KEYINPUT67), .A3(new_n466), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n474), .A2(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g059(.A(KEYINPUT69), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(G136), .B2(new_n467), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n476), .A2(new_n477), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  OAI211_X1 g076(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n500), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n501), .B1(new_n500), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n515), .B1(KEYINPUT5), .B2(new_n512), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(G543), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G166));
  AND2_X1   g101(.A1(new_n516), .A2(new_n520), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n520), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n528), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n518), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n529), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n516), .A2(G90), .A3(new_n520), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n537), .B(KEYINPUT73), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G171));
  AOI22_X1  g122(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n518), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT74), .B(G43), .Z(new_n551));
  OAI22_X1  g126(.A1(new_n521), .A2(new_n550), .B1(new_n524), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n529), .A2(new_n560), .A3(G53), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n524), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n527), .A2(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n518), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  NAND3_X1  g148(.A1(new_n520), .A2(G49), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT75), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n520), .A2(new_n576), .A3(G49), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n516), .A2(G87), .A3(new_n520), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n521), .A2(new_n582), .B1(new_n583), .B2(new_n524), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n516), .A2(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n518), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n513), .A2(new_n515), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n521), .A2(new_n598), .B1(new_n599), .B2(new_n524), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n597), .A2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(new_n527), .A2(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n593), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G868), .B2(G171), .ZN(G284));
  XOR2_X1   g186(.A(G284), .B(KEYINPUT76), .Z(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n569), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(G868), .B2(new_n569), .ZN(G280));
  INV_X1    g190(.A(new_n609), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(G111), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G2105), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G135), .B2(new_n467), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n486), .B2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n476), .A2(new_n477), .A3(new_n461), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT13), .B(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT80), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT79), .ZN(new_n645));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n643), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n656), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n659), .B2(new_n655), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2096), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(KEYINPUT83), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT20), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT84), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n689), .A2(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  OR2_X1    g271(.A1(G95), .A2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT85), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G131), .B2(new_n467), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n487), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n696), .B1(new_n703), .B2(new_n695), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT86), .Z(new_n706));
  XOR2_X1   g281(.A(new_n704), .B(new_n706), .Z(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G24), .ZN(new_n710));
  INV_X1    g285(.A(G290), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT87), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n709), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT33), .B(G1976), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n717), .B(new_n718), .Z(new_n719));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n709), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G166), .B2(new_n709), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G6), .A2(G16), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n588), .B2(G16), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT32), .B(G1981), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n721), .A2(new_n722), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n714), .B1(new_n708), .B2(new_n713), .C1(new_n731), .C2(KEYINPUT34), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT89), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT36), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n695), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n695), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT29), .Z(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT97), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n695), .A2(G33), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n476), .A2(new_n477), .A3(G127), .ZN(new_n744));
  INV_X1    g319(.A(G115), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n460), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n469), .B1(new_n746), .B2(KEYINPUT90), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT90), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n749));
  NAND2_X1  g324(.A1(G103), .A2(G2104), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G2105), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n469), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n467), .A2(G139), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n743), .B1(new_n754), .B2(new_n695), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G2072), .Z(new_n756));
  NOR2_X1   g331(.A1(G4), .A2(G16), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n616), .B2(G16), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n739), .A2(new_n740), .B1(G1348), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n709), .A2(G19), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n554), .B2(new_n709), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1341), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n695), .A2(G27), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT96), .Z(new_n765));
  INV_X1    g340(.A(G164), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G29), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  AND4_X1   g343(.A1(new_n742), .A2(new_n756), .A3(new_n759), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G5), .A2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT94), .Z(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G171), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  INV_X1    g348(.A(G1961), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n709), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n709), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT93), .B(G1966), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n767), .A2(new_n763), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n630), .A2(G29), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n695), .A2(G32), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n461), .A2(G105), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT26), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n784), .B(new_n786), .C1(G141), .C2(new_n467), .ZN(new_n787));
  INV_X1    g362(.A(G129), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n486), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n782), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n780), .A2(new_n781), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n695), .A2(G26), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT28), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n487), .A2(G128), .ZN(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n797));
  INV_X1    g372(.A(G116), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G2105), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G140), .B2(new_n467), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(G28), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n695), .B1(new_n804), .B2(G28), .ZN(new_n806));
  AND2_X1   g381(.A1(KEYINPUT31), .A2(G11), .ZN(new_n807));
  NOR2_X1   g382(.A1(KEYINPUT31), .A2(G11), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n790), .B2(new_n791), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G2084), .ZN(new_n812));
  AND2_X1   g387(.A1(KEYINPUT24), .A2(G34), .ZN(new_n813));
  NOR2_X1   g388(.A1(KEYINPUT24), .A2(G34), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n695), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT91), .Z(new_n816));
  INV_X1    g391(.A(G160), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n695), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n811), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n709), .A2(G20), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT23), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n569), .B2(new_n709), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1956), .ZN(new_n823));
  INV_X1    g398(.A(new_n758), .ZN(new_n824));
  INV_X1    g399(.A(G1348), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n818), .A2(new_n812), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT92), .ZN(new_n828));
  AND4_X1   g403(.A1(new_n793), .A2(new_n819), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n769), .A2(new_n775), .A3(new_n776), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n736), .A2(new_n830), .ZN(G311));
  INV_X1    g406(.A(G311), .ZN(G150));
  AOI22_X1  g407(.A1(new_n527), .A2(G93), .B1(G55), .B2(new_n529), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n516), .A2(G67), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G651), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT98), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n553), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT38), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n616), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n838), .A2(new_n845), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  INV_X1    g425(.A(G37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n500), .A2(new_n507), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n789), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n801), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n754), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n702), .B(new_n633), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n487), .A2(G130), .ZN(new_n860));
  AOI211_X1 g435(.A(new_n859), .B(new_n860), .C1(G142), .C2(new_n467), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n856), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(new_n862), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n630), .B(KEYINPUT99), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n817), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n493), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n863), .A2(new_n869), .A3(new_n864), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n855), .A2(new_n869), .A3(new_n862), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n867), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n851), .B(new_n868), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g449(.A(G868), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n609), .A2(new_n569), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT101), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n616), .A2(G299), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT102), .B1(new_n616), .B2(G299), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n876), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(KEYINPUT41), .B2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n840), .B(new_n619), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(G166), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n588), .B(G288), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(new_n887), .B2(new_n893), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n875), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n838), .A2(G868), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n897), .A2(new_n898), .ZN(G331));
  NAND2_X1  g474(.A1(G331), .A2(KEYINPUT104), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n897), .A2(KEYINPUT104), .A3(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(G295));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  XNOR2_X1  g478(.A(G171), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G168), .ZN(new_n905));
  XNOR2_X1  g480(.A(G171), .B(KEYINPUT105), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G286), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n840), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n840), .A2(new_n905), .A3(new_n907), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n884), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n840), .A2(new_n905), .A3(new_n907), .A4(KEYINPUT106), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n905), .A2(new_n907), .ZN(new_n917));
  INV_X1    g492(.A(new_n840), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n917), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n913), .B(new_n914), .C1(new_n916), .C2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n890), .B(new_n911), .C1(new_n920), .C2(new_n880), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n851), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n908), .B(new_n915), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n913), .A2(new_n914), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n879), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n890), .B1(new_n925), .B2(new_n911), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n890), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n880), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n929), .B2(new_n883), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n923), .B2(new_n924), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n910), .A2(new_n908), .A3(new_n880), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n851), .A4(new_n921), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n922), .B2(new_n926), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n851), .A3(new_n921), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  MUX2_X1   g515(.A(new_n937), .B(new_n940), .S(KEYINPUT44), .Z(G397));
  AOI21_X1  g516(.A(new_n506), .B1(new_n499), .B2(new_n497), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  XNOR2_X1  g518(.A(KEYINPUT108), .B(G1384), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n478), .A2(new_n479), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(G2105), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n467), .A2(new_n463), .A3(G137), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n948), .A2(new_n949), .B1(G101), .B2(new_n461), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(G40), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n852), .A2(KEYINPUT70), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n942), .A2(new_n501), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n952), .B1(new_n955), .B2(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n725), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n508), .B2(new_n509), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n942), .A2(G1384), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n951), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n740), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G8), .ZN(new_n966));
  NOR2_X1   g541(.A1(G166), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT55), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(G8), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(G160), .A2(new_n962), .A3(G40), .ZN(new_n970));
  INV_X1    g545(.A(G1976), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n578), .A2(G1976), .A3(new_n579), .A4(new_n580), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n970), .A2(new_n972), .A3(G8), .A4(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT110), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n527), .A2(G86), .B1(G48), .B2(new_n529), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n585), .A2(new_n586), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G651), .ZN(new_n978));
  INV_X1    g553(.A(G1981), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n852), .A2(new_n958), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n951), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n966), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n981), .A3(KEYINPUT49), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n970), .A2(G8), .A3(new_n973), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT52), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n969), .A2(new_n975), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n970), .A2(G8), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(new_n971), .A3(new_n716), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(new_n980), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n975), .A2(new_n992), .A3(KEYINPUT111), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT49), .B1(new_n980), .B2(new_n981), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n994), .A2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1001), .A2(new_n988), .B1(KEYINPUT52), .B2(new_n990), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n987), .A2(KEYINPUT110), .A3(new_n973), .A4(new_n972), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n974), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n999), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n998), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n961), .B1(new_n852), .B2(new_n958), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(new_n951), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n961), .B(new_n958), .C1(new_n508), .C2(new_n509), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n740), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n966), .B1(new_n957), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n969), .B1(new_n968), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT45), .B1(new_n852), .B2(new_n958), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(new_n951), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n958), .C1(new_n508), .C2(new_n509), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1966), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(KEYINPUT112), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n960), .A2(new_n812), .A3(new_n963), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT112), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1016), .B1(new_n1026), .B2(G286), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n1023), .A3(new_n1022), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(KEYINPUT113), .A3(G8), .A4(G168), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT63), .B1(new_n1015), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n968), .ZN(new_n1035));
  INV_X1    g610(.A(new_n965), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n966), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n975), .A2(new_n992), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(KEYINPUT63), .A3(new_n1038), .A4(new_n969), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1032), .B2(new_n1027), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n997), .B1(new_n1034), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n960), .A2(new_n963), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n825), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(G2067), .B2(new_n970), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(KEYINPUT60), .B2(new_n616), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(G1341), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n986), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n944), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(G160), .A3(G40), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n943), .B2(new_n959), .ZN(new_n1057));
  INV_X1    g632(.A(G1996), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1053), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT117), .B1(new_n1059), .B2(new_n553), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1053), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n952), .B(new_n1058), .C1(new_n955), .C2(KEYINPUT45), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n554), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1067));
  INV_X1    g642(.A(G1956), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT114), .B(KEYINPUT57), .C1(new_n566), .C2(new_n568), .ZN(new_n1070));
  INV_X1    g645(.A(new_n568), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n563), .A2(new_n561), .B1(new_n527), .B2(G91), .ZN(new_n1072));
  OR2_X1    g647(.A1(KEYINPUT114), .A2(KEYINPUT57), .ZN(new_n1073));
  NAND2_X1  g648(.A1(KEYINPUT114), .A2(KEYINPUT57), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT115), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n952), .B(new_n1079), .C1(new_n955), .C2(KEYINPUT45), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1069), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1069), .B2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT61), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1080), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1956), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1076), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1069), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1050), .A2(new_n1066), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1060), .A2(KEYINPUT59), .A3(new_n1065), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1049), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1064), .B1(new_n1063), .B2(new_n554), .ZN(new_n1094));
  AOI211_X1 g669(.A(KEYINPUT117), .B(new_n553), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1050), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AND4_X1   g671(.A1(new_n1049), .A2(new_n1093), .A3(new_n1091), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1048), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1086), .B1(new_n1045), .B2(new_n609), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1088), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT124), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT111), .B1(new_n975), .B2(new_n992), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1002), .A2(new_n1006), .A3(new_n999), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1013), .A2(new_n968), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n969), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1057), .A2(new_n763), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1042), .A2(new_n774), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1018), .A2(new_n1019), .A3(KEYINPUT53), .A4(new_n763), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1112), .A2(KEYINPUT121), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT121), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1111), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n545), .A2(new_n1118), .A3(new_n546), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1112), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1042), .A2(KEYINPUT122), .A3(new_n774), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1123), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n474), .A2(KEYINPUT123), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1110), .A2(G2078), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1126), .A2(G40), .A3(new_n947), .A4(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT45), .B1(new_n852), .B2(new_n1054), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n474), .A2(KEYINPUT123), .ZN(new_n1130));
  NOR4_X1   g705(.A1(new_n1128), .A2(new_n945), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1116), .A2(new_n1121), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1102), .A2(new_n1108), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G168), .A2(new_n966), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1136), .B2(KEYINPUT119), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1026), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(G8), .B(new_n1138), .C1(new_n1031), .C2(G286), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1024), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1136), .B1(new_n1143), .B2(new_n1030), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1142), .A2(KEYINPUT120), .A3(new_n1145), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1134), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1041), .B1(new_n1101), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1148), .A2(new_n1152), .A3(new_n1149), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT120), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n1147), .B(new_n1144), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT62), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1116), .A2(G171), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1102), .A2(new_n1108), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1153), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT125), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1153), .A2(new_n1156), .A3(new_n1161), .A4(new_n1158), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1151), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n951), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1129), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n711), .A2(new_n708), .ZN(new_n1167));
  NOR2_X1   g742(.A1(G290), .A2(G1986), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT109), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n801), .A2(G2067), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n801), .A2(G2067), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n789), .B(new_n1058), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n702), .B(new_n705), .Z(new_n1176));
  OAI21_X1  g751(.A(new_n1166), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1163), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1168), .A2(new_n1166), .A3(KEYINPUT48), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1168), .A2(new_n1166), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT48), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1177), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1173), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1166), .B1(new_n1185), .B2(new_n789), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT46), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1166), .B2(new_n1058), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1165), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT47), .Z(new_n1191));
  NAND2_X1  g766(.A1(new_n703), .A2(new_n705), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1171), .B1(new_n1175), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g768(.A(new_n1184), .B(new_n1191), .C1(new_n1166), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1179), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1179), .A2(KEYINPUT126), .A3(new_n1194), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  OR3_X1    g775(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1202), .B1(new_n689), .B2(new_n693), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1203), .A2(new_n873), .ZN(new_n1204));
  INV_X1    g778(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1201), .B1(new_n937), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g780(.A(KEYINPUT127), .B(new_n1204), .C1(new_n927), .C2(new_n936), .ZN(new_n1207));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n1207), .ZN(G308));
  NAND2_X1  g782(.A1(new_n937), .A2(new_n1205), .ZN(G225));
endmodule


