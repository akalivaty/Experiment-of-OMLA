//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n963, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202));
  AOI21_X1  g001(.A(G190gat), .B1(new_n202), .B2(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT27), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(KEYINPUT28), .A3(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT70), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n203), .A2(KEYINPUT70), .A3(KEYINPUT28), .A4(new_n205), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n202), .B2(G183gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n204), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n203), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n214), .A2(KEYINPUT69), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT69), .B1(new_n214), .B2(new_n215), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT71), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n220), .B(new_n210), .C1(new_n216), .C2(new_n217), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(KEYINPUT26), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n226), .B1(new_n231), .B2(KEYINPUT26), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n221), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT72), .ZN(new_n237));
  INV_X1    g036(.A(G113gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(G120gat), .ZN(new_n240));
  INV_X1    g039(.A(G120gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT73), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n239), .A2(new_n242), .A3(new_n245), .A4(new_n240), .ZN(new_n246));
  INV_X1    g045(.A(G134gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G127gat), .ZN(new_n248));
  INV_X1    g047(.A(G127gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G134gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n244), .A2(new_n246), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n240), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n238), .A2(G120gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n248), .A2(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT23), .ZN(new_n261));
  INV_X1    g060(.A(new_n224), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n265), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT23), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT65), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT23), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n227), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G183gat), .B(G190gat), .Z(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT24), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n233), .A2(KEYINPUT24), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n267), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n272), .A2(new_n224), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n225), .B2(new_n268), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n227), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n280), .A2(new_n284), .A3(new_n276), .A4(new_n277), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n273), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n236), .A2(new_n260), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n260), .B1(new_n236), .B2(new_n287), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G227gat), .ZN(new_n291));
  INV_X1    g090(.A(G233gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT34), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT34), .ZN(new_n295));
  INV_X1    g094(.A(new_n293), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n295), .B(new_n296), .C1(new_n288), .C2(new_n289), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT33), .B1(new_n290), .B2(new_n293), .ZN(new_n298));
  XNOR2_X1  g097(.A(G15gat), .B(G43gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT74), .ZN(new_n300));
  INV_X1    g099(.A(G71gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(G99gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n294), .B(new_n297), .C1(new_n298), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n236), .A2(new_n287), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n252), .B1(new_n243), .B2(KEYINPUT73), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n306), .A2(new_n246), .B1(new_n257), .B2(new_n258), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n267), .A2(new_n278), .B1(new_n285), .B2(new_n273), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n234), .B1(new_n218), .B2(KEYINPUT71), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n221), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n260), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n312), .A3(new_n293), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT33), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n303), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(new_n312), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n295), .B1(new_n316), .B2(new_n296), .ZN(new_n317));
  INV_X1    g116(.A(new_n297), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(KEYINPUT32), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT85), .B(G22gat), .Z(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G197gat), .B(G204gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327));
  INV_X1    g126(.A(G211gat), .ZN(new_n328));
  INV_X1    g127(.A(G218gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT84), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n330), .ZN(new_n333));
  INV_X1    g132(.A(new_n325), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n325), .A2(new_n326), .A3(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n331), .B(new_n332), .C1(new_n337), .C2(KEYINPUT84), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT2), .ZN(new_n342));
  INV_X1    g141(.A(G141gat), .ZN(new_n343));
  INV_X1    g142(.A(G148gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OR2_X1    g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n341), .ZN(new_n350));
  AND2_X1   g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT80), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  AND2_X1   g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n355), .A2(new_n358), .A3(new_n349), .A4(new_n342), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT81), .B1(new_n360), .B2(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(new_n359), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n339), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n361), .B1(new_n366), .B2(new_n337), .ZN(new_n367));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n368), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT3), .B1(new_n337), .B2(new_n332), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(new_n363), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n362), .A2(new_n365), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n332), .ZN(new_n374));
  INV_X1    g173(.A(new_n337), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n324), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  OAI221_X1 g176(.A(new_n370), .B1(new_n363), .B2(new_n371), .C1(new_n366), .C2(new_n337), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n374), .A2(new_n375), .B1(new_n360), .B2(new_n340), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n378), .B(new_n323), .C1(new_n379), .C2(new_n370), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT31), .B(G50gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT86), .B1(new_n369), .B2(new_n376), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n378), .B(new_n388), .C1(new_n379), .C2(new_n370), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n387), .A2(G22gat), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n376), .B1(new_n368), .B2(new_n367), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT87), .A3(new_n323), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n380), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n394), .A3(new_n384), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n386), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n321), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n304), .A2(new_n319), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n322), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT76), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n311), .B2(KEYINPUT29), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT77), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(new_n305), .B2(new_n401), .ZN(new_n405));
  AOI211_X1 g204(.A(KEYINPUT77), .B(new_n402), .C1(new_n236), .C2(new_n287), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n375), .B(new_n403), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G64gat), .B(G92gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n401), .B1(new_n305), .B2(new_n332), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n402), .B1(new_n236), .B2(new_n287), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n337), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n407), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n407), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT78), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G1gat), .B(G29gat), .Z(new_n419));
  XNOR2_X1  g218(.A(G57gat), .B(G85gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n254), .A2(new_n363), .A3(new_n259), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT82), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n307), .A2(new_n427), .A3(new_n363), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n260), .A2(new_n360), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n424), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n426), .A2(new_n428), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n364), .B1(new_n363), .B2(new_n339), .ZN(new_n437));
  AOI211_X1 g236(.A(KEYINPUT81), .B(KEYINPUT3), .C1(new_n354), .C2(new_n359), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n260), .B(new_n436), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n307), .A2(KEYINPUT4), .A3(new_n363), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n435), .A2(new_n439), .A3(new_n440), .A4(new_n431), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n433), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n307), .B1(KEYINPUT3), .B2(new_n360), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n432), .B1(new_n373), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n428), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT4), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n434), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n424), .A4(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n423), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(new_n448), .A3(new_n423), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n451), .B(new_n423), .C1(new_n442), .C2(new_n448), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n407), .A2(new_n411), .A3(new_n414), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n305), .A2(new_n401), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n375), .B1(new_n403), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT77), .B1(new_n311), .B2(new_n402), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n305), .A2(new_n404), .A3(new_n401), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n305), .A2(new_n332), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n461), .A2(new_n462), .B1(new_n463), .B2(new_n402), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n460), .B1(new_n464), .B2(new_n375), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n457), .B(new_n458), .C1(new_n465), .C2(new_n416), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n465), .B2(new_n411), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n418), .A2(new_n456), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT35), .B1(new_n399), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n304), .A2(new_n397), .A3(new_n319), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n397), .B1(new_n304), .B2(new_n319), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n456), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n407), .A2(new_n414), .ZN(new_n476));
  INV_X1    g275(.A(new_n416), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n411), .B1(new_n407), .B2(new_n414), .ZN(new_n479));
  INV_X1    g278(.A(new_n467), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n478), .B(new_n457), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n473), .A2(new_n475), .A3(new_n396), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n470), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(KEYINPUT40), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n446), .A2(new_n447), .A3(new_n439), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n432), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n423), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT39), .B1(new_n430), .B2(new_n432), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n487), .B2(new_n432), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n486), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n492), .ZN(new_n494));
  INV_X1    g293(.A(new_n486), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n423), .A3(new_n495), .A4(new_n489), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n493), .A2(new_n496), .A3(new_n450), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n396), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n411), .A2(KEYINPUT37), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n457), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n407), .A2(KEYINPUT37), .A3(new_n414), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n504), .B2(KEYINPUT38), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n452), .A2(new_n451), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(new_n449), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n507), .A2(new_n479), .A3(new_n454), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n337), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n413), .B1(new_n463), .B2(new_n402), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n375), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT38), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n502), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT38), .ZN(new_n518));
  AOI211_X1 g317(.A(KEYINPUT89), .B(new_n518), .C1(new_n502), .C2(new_n503), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n499), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n384), .B1(new_n377), .B2(new_n380), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n384), .B1(new_n380), .B2(new_n393), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT87), .B1(new_n391), .B2(new_n323), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n387), .A2(G22gat), .A3(new_n389), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n469), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(KEYINPUT75), .B(KEYINPUT36), .C1(new_n471), .C2(new_n472), .ZN(new_n529));
  NAND2_X1  g328(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n530));
  OR2_X1    g329(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n322), .A2(new_n530), .A3(new_n531), .A4(new_n398), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n484), .B1(new_n521), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n484), .B(KEYINPUT90), .C1(new_n521), .C2(new_n533), .ZN(new_n537));
  INV_X1    g336(.A(G43gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G50gat), .ZN(new_n539));
  INV_X1    g338(.A(G50gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G43gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n541), .A3(KEYINPUT15), .ZN(new_n542));
  NOR2_X1   g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT14), .Z(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT91), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n544), .A2(KEYINPUT91), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(KEYINPUT92), .B(G50gat), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n538), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n550), .A2(KEYINPUT93), .B1(G43gat), .B2(new_n540), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n552), .A3(new_n538), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT15), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G29gat), .A2(G36gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n544), .A2(new_n542), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n548), .B(KEYINPUT17), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558));
  INV_X1    g357(.A(G1gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT16), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G8gat), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n561), .B(new_n562), .C1(G1gat), .C2(new_n558), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n558), .A2(new_n560), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n561), .B(KEYINPUT94), .C1(G1gat), .C2(new_n558), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n566), .A2(KEYINPUT95), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT95), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n563), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n554), .A2(new_n556), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n547), .ZN(new_n575));
  OAI211_X1 g374(.A(KEYINPUT96), .B(new_n563), .C1(new_n568), .C2(new_n569), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n557), .A2(new_n572), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n570), .B1(new_n547), .B2(new_n574), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OR3_X1    g381(.A1(new_n570), .A2(new_n547), .A3(new_n574), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n579), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n578), .B(KEYINPUT13), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n577), .A2(KEYINPUT18), .A3(new_n578), .A4(new_n579), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G197gat), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT11), .B(G169gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT12), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n580), .A2(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n595));
  INV_X1    g394(.A(new_n593), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n587), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n536), .A2(new_n537), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT97), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n536), .A2(new_n601), .A3(new_n537), .A4(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G57gat), .B(G64gat), .Z(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  INV_X1    g404(.A(G78gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n301), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G71gat), .B(G78gat), .Z(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n613));
  AND2_X1   g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT20), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n570), .B1(KEYINPUT21), .B2(new_n612), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT99), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n618), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G190gat), .B(G218gat), .Z(new_n629));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n630));
  NAND2_X1  g429(.A1(G85gat), .A2(G92gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT7), .ZN(new_n632));
  XOR2_X1   g431(.A(G99gat), .B(G106gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(G85gat), .A2(G92gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(G99gat), .A2(G106gat), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(KEYINPUT8), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n632), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n634), .B1(new_n632), .B2(new_n637), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n557), .A2(new_n575), .A3(new_n630), .A4(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n574), .B2(new_n547), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644));
  NAND3_X1  g443(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n643), .B2(new_n645), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n557), .A2(new_n575), .A3(new_n641), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(KEYINPUT100), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n629), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n647), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n629), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n649), .A2(KEYINPUT100), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .A4(new_n642), .ZN(new_n657));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n651), .B2(new_n657), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G230gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n292), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n612), .A2(new_n640), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT10), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n610), .A2(new_n611), .ZN(new_n672));
  OAI22_X1  g471(.A1(new_n672), .A2(new_n668), .B1(new_n638), .B2(new_n639), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n612), .A2(new_n640), .A3(KEYINPUT10), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n667), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n673), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n667), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n677), .A2(new_n679), .A3(new_n683), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n628), .A2(new_n665), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n603), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n456), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(new_n559), .ZN(G1324gat));
  XNOR2_X1  g492(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G8gat), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n603), .A2(new_n481), .A3(new_n690), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT103), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(KEYINPUT103), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G8gat), .B1(new_n691), .B2(new_n482), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(G1325gat));
  AND2_X1   g501(.A1(new_n529), .A2(new_n532), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n691), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n473), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n691), .B2(new_n706), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n396), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(new_n628), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n664), .A3(new_n688), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT105), .Z(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n600), .B2(new_n602), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n456), .A2(G29gat), .ZN(new_n717));
  OR3_X1    g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n527), .B1(new_n481), .B2(new_n497), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n518), .B1(new_n502), .B2(new_n503), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n515), .B(new_n508), .C1(new_n720), .C2(new_n500), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n721), .B2(new_n519), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n469), .A2(KEYINPUT106), .A3(new_n527), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n528), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n703), .A2(new_n722), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n470), .A2(new_n483), .A3(KEYINPUT107), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT107), .B1(new_n470), .B2(new_n483), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n664), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n665), .A2(new_n731), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n536), .A2(new_n537), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n598), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n628), .A2(new_n735), .A3(new_n687), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n456), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n716), .B1(new_n715), .B2(new_n717), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n718), .A2(new_n738), .A3(new_n739), .ZN(G1328gat));
  NOR2_X1   g539(.A1(new_n482), .A2(G36gat), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n742), .B(new_n713), .C1(new_n600), .C2(new_n602), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n536), .A2(new_n537), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n745), .A2(new_n733), .B1(new_n731), .B2(new_n730), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n481), .A3(new_n736), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n743), .A2(new_n744), .B1(new_n747), .B2(G36gat), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT108), .B1(new_n743), .B2(new_n744), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n750), .B(KEYINPUT46), .C1(new_n715), .C2(new_n742), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(G1329gat));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n754));
  INV_X1    g553(.A(new_n703), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n732), .A2(new_n755), .A3(new_n734), .A4(new_n736), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(G43gat), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n705), .A2(G43gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n714), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n753), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n713), .ZN(new_n761));
  AND4_X1   g560(.A1(KEYINPUT110), .A2(new_n603), .A3(new_n761), .A4(new_n758), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT110), .B1(new_n714), .B2(new_n758), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n756), .A2(new_n765), .A3(G43gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n757), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n760), .B1(new_n764), .B2(new_n767), .ZN(G1330gat));
  OAI21_X1  g567(.A(new_n549), .B1(new_n737), .B2(new_n396), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n396), .A2(new_n549), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n715), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n769), .B(KEYINPUT48), .C1(new_n715), .C2(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1331gat));
  NOR4_X1   g574(.A1(new_n711), .A2(new_n598), .A3(new_n664), .A4(new_n688), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n729), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n474), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g579(.A1(new_n777), .A2(new_n482), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  NOR3_X1   g584(.A1(new_n777), .A2(G71gat), .A3(new_n705), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n778), .A2(new_n755), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(G71gat), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g588(.A1(new_n777), .A2(new_n396), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(new_n606), .ZN(G1335gat));
  NOR3_X1   g590(.A1(new_n628), .A2(new_n598), .A3(new_n688), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n732), .A2(new_n734), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n456), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n628), .A2(new_n598), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n729), .A2(new_n664), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n729), .A2(KEYINPUT51), .A3(new_n664), .A4(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n456), .A2(new_n688), .A3(G85gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT111), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n794), .A2(new_n805), .A3(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1336gat));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  OAI21_X1  g607(.A(G92gat), .B1(new_n793), .B2(new_n482), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n482), .A2(G92gat), .A3(new_n688), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n800), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n810), .B1(new_n800), .B2(new_n811), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n808), .B(new_n809), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n811), .B(KEYINPUT112), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n808), .B2(new_n817), .ZN(G1337gat));
  OAI21_X1  g617(.A(G99gat), .B1(new_n793), .B2(new_n703), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n688), .A2(G99gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n473), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1338gat));
  OAI21_X1  g621(.A(KEYINPUT115), .B1(new_n793), .B2(new_n396), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n746), .A2(new_n824), .A3(new_n527), .A4(new_n792), .ZN(new_n825));
  XNOR2_X1  g624(.A(KEYINPUT114), .B(G106gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n396), .A2(G106gat), .A3(new_n688), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT53), .B1(new_n800), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n826), .B1(new_n793), .B2(new_n396), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n800), .A2(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n835), .ZN(G1339gat));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n838), .A2(new_n839), .B1(new_n584), .B2(new_n585), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n592), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n597), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n674), .A2(new_n667), .A3(new_n675), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n677), .A2(KEYINPUT54), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n683), .B1(new_n676), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(KEYINPUT55), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT116), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n846), .A2(new_n851), .A3(KEYINPUT55), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n686), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n846), .A2(new_n848), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n844), .A2(new_n664), .A3(new_n853), .A4(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n597), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n596), .B1(new_n595), .B2(new_n587), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n853), .B(new_n857), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n842), .A2(new_n597), .A3(new_n687), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n837), .B(new_n858), .C1(new_n863), .C2(new_n664), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n664), .B1(new_n861), .B2(new_n862), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n651), .A2(new_n657), .ZN(new_n866));
  INV_X1    g665(.A(new_n660), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n868), .A2(new_n853), .A3(new_n661), .A4(new_n857), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n843), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT118), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n864), .A2(new_n711), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n690), .A2(new_n735), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n399), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n874), .A2(new_n474), .A3(new_n482), .A4(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n238), .A3(new_n735), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n874), .A2(new_n474), .A3(new_n875), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT119), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n456), .B1(new_n872), .B2(new_n873), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n875), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n482), .A3(new_n598), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n877), .B1(new_n884), .B2(new_n238), .ZN(G1340gat));
  NOR3_X1   g684(.A1(new_n876), .A2(new_n241), .A3(new_n688), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n883), .A2(new_n482), .A3(new_n687), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n241), .ZN(G1341gat));
  NOR3_X1   g687(.A1(new_n876), .A2(new_n249), .A3(new_n711), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n481), .B(new_n711), .C1(new_n879), .C2(new_n882), .ZN(new_n890));
  AOI21_X1  g689(.A(G127gat), .B1(new_n890), .B2(KEYINPUT120), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n883), .A2(new_n482), .A3(new_n628), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n889), .B1(new_n891), .B2(new_n894), .ZN(G1342gat));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n664), .A2(new_n482), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT121), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n247), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n897), .B1(new_n883), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT122), .B(new_n900), .C1(new_n879), .C2(new_n882), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n896), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n878), .A2(KEYINPUT119), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n881), .B1(new_n880), .B2(new_n875), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n883), .A2(new_n897), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(KEYINPUT56), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G134gat), .B1(new_n876), .B2(new_n665), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(G1343gat));
  NOR3_X1   g711(.A1(new_n755), .A2(new_n456), .A3(new_n481), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n874), .B2(new_n527), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n527), .A2(KEYINPUT57), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n711), .B1(new_n865), .B2(new_n870), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n873), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G141gat), .B1(new_n918), .B2(new_n735), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n880), .A2(new_n527), .A3(new_n703), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n920), .A2(new_n343), .A3(new_n482), .A4(new_n598), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT58), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT58), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n919), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1344gat));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n915), .B1(new_n872), .B2(new_n873), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT123), .B(new_n858), .C1(new_n863), .C2(new_n664), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n865), .B2(new_n870), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n930), .A2(new_n711), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n396), .B1(new_n933), .B2(new_n873), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n934), .B2(KEYINPUT57), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n687), .A3(new_n913), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n927), .B1(new_n936), .B2(G148gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n927), .A2(G148gat), .ZN(new_n938));
  INV_X1    g737(.A(new_n918), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n687), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n482), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n687), .A2(new_n344), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n937), .A2(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1345gat));
  NOR2_X1   g742(.A1(new_n941), .A2(new_n711), .ZN(new_n944));
  AOI21_X1  g743(.A(G155gat), .B1(new_n944), .B2(KEYINPUT124), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n941), .B2(new_n711), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n628), .A2(G155gat), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT125), .Z(new_n949));
  AOI22_X1  g748(.A1(new_n945), .A2(new_n947), .B1(new_n939), .B2(new_n949), .ZN(G1346gat));
  OAI21_X1  g749(.A(G162gat), .B1(new_n918), .B2(new_n665), .ZN(new_n951));
  INV_X1    g750(.A(G162gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n920), .A2(new_n952), .A3(new_n899), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n951), .A2(KEYINPUT126), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1347gat));
  NOR2_X1   g757(.A1(new_n482), .A2(new_n474), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n874), .A2(new_n875), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n598), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n687), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g763(.A1(new_n960), .A2(new_n202), .A3(new_n628), .ZN(new_n965));
  XNOR2_X1  g764(.A(KEYINPUT60), .B(G183gat), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n965), .B(new_n966), .ZN(G1350gat));
  NOR2_X1   g766(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n968), .B1(new_n960), .B2(new_n664), .ZN(new_n969));
  NAND2_X1  g768(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n969), .B(new_n970), .Z(G1351gat));
  AND2_X1   g770(.A1(new_n703), .A2(new_n959), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n874), .A2(new_n527), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n598), .ZN(new_n974));
  INV_X1    g773(.A(new_n935), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n972), .B(KEYINPUT127), .Z(new_n976));
  NOR2_X1   g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n598), .A2(G197gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  INV_X1    g778(.A(G204gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n973), .A2(new_n980), .A3(new_n687), .ZN(new_n981));
  XOR2_X1   g780(.A(new_n981), .B(KEYINPUT62), .Z(new_n982));
  NAND2_X1  g781(.A1(new_n935), .A2(new_n687), .ZN(new_n983));
  OAI21_X1  g782(.A(G204gat), .B1(new_n983), .B2(new_n976), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1353gat));
  NAND3_X1  g784(.A1(new_n973), .A2(new_n328), .A3(new_n628), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n935), .A2(new_n628), .A3(new_n972), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(G1354gat));
  AOI21_X1  g789(.A(G218gat), .B1(new_n973), .B2(new_n664), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n665), .A2(new_n329), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n991), .B1(new_n977), .B2(new_n992), .ZN(G1355gat));
endmodule


