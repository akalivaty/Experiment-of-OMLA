//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT65), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n212), .B(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT66), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n221), .B(new_n222), .C1(new_n217), .C2(new_n218), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT67), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n211), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  INV_X1    g0029(.A(G58), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n235), .A2(new_n209), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n229), .B(new_n237), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n226), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT68), .ZN(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XOR2_X1   g0053(.A(G107), .B(G116), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  NAND2_X1  g0056(.A1(new_n202), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n209), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n209), .A2(G33), .ZN(new_n261));
  OR3_X1    g0061(.A1(new_n230), .A2(KEYINPUT70), .A3(KEYINPUT71), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(KEYINPUT70), .B2(new_n230), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n230), .A2(KEYINPUT71), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n262), .A2(new_n264), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n257), .B1(new_n258), .B2(new_n260), .C1(new_n261), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n270), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n235), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT72), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(new_n209), .B2(G1), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n208), .A2(KEYINPUT72), .A3(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n269), .A2(new_n271), .A3(new_n235), .A4(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G50), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n279), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n282), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n273), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n259), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n290), .A2(G223), .B1(new_n293), .B2(G77), .ZN(new_n294));
  INV_X1    g0094(.A(G222), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n289), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n286), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(new_n235), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(G274), .B1(new_n299), .B2(new_n235), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n235), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n303), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n304), .B1(new_n309), .B2(G226), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n285), .B1(G169), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n312), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(G190), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  INV_X1    g0117(.A(new_n285), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n316), .B1(new_n317), .B2(new_n312), .C1(new_n318), .C2(KEYINPUT9), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT9), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n285), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n320), .B(new_n321), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n323), .B(KEYINPUT73), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT10), .B1(new_n328), .B2(new_n319), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n315), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G159), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n260), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT70), .B(G58), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n232), .B1(new_n334), .B2(new_n231), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n333), .B1(new_n335), .B2(G20), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n288), .A2(new_n209), .A3(new_n289), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n289), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT77), .B1(new_n341), .B2(G68), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  AOI211_X1 g0143(.A(new_n343), .B(new_n231), .C1(new_n339), .C2(new_n340), .ZN(new_n344));
  OAI211_X1 g0144(.A(KEYINPUT16), .B(new_n336), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n269), .A2(new_n235), .A3(new_n271), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT7), .B1(new_n293), .B2(new_n209), .ZN(new_n347));
  INV_X1    g0147(.A(new_n340), .ZN(new_n348));
  OAI21_X1  g0148(.A(G68), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n336), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n308), .A2(new_n241), .B1(new_n302), .B2(new_n303), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G223), .A2(G1698), .ZN(new_n357));
  INV_X1    g0157(.A(G226), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(G1698), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(new_n296), .B1(G33), .B2(G87), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n300), .B1(new_n360), .B2(KEYINPUT78), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G87), .ZN(new_n362));
  OR2_X1    g0162(.A1(G223), .A2(G1698), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n362), .B1(new_n365), .B2(new_n293), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT78), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n354), .B(new_n356), .C1(new_n361), .C2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n307), .B1(new_n366), .B2(new_n367), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n355), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n369), .B1(G200), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n266), .A2(new_n278), .ZN(new_n374));
  INV_X1    g0174(.A(new_n280), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n374), .A2(new_n375), .B1(new_n283), .B2(new_n266), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n353), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT79), .A2(KEYINPUT17), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n353), .A2(new_n376), .ZN(new_n380));
  INV_X1    g0180(.A(G169), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n370), .A2(new_n371), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n356), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n314), .B(new_n355), .C1(new_n370), .C2(new_n371), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT18), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n380), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n376), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n345), .B2(new_n352), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n383), .A2(new_n384), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT18), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g0191(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n373), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n379), .A2(new_n387), .A3(new_n391), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G20), .A2(G77), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT8), .B(G58), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n396), .B1(new_n397), .B2(new_n261), .C1(new_n260), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n272), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n375), .A2(G77), .A3(new_n277), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(G77), .C2(new_n279), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n290), .A2(G238), .B1(new_n293), .B2(G107), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n296), .A2(G232), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(G1698), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n300), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n304), .B1(new_n309), .B2(G244), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n402), .B1(new_n408), .B2(G190), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n317), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n314), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n407), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n381), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n402), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n395), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G97), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n416), .B1(new_n297), .B2(new_n358), .C1(new_n286), .C2(new_n404), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n300), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n419));
  AOI21_X1  g0219(.A(new_n304), .B1(new_n309), .B2(G238), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n419), .B1(new_n418), .B2(new_n420), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(G169), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n418), .A2(new_n420), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n427), .A2(KEYINPUT75), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT13), .B1(new_n427), .B2(KEYINPUT75), .ZN(new_n429));
  OAI211_X1 g0229(.A(G179), .B(new_n421), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G169), .B1(new_n422), .B2(new_n423), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n278), .A2(new_n280), .A3(new_n231), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT76), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n260), .A2(new_n281), .B1(new_n209), .B2(G68), .ZN(new_n436));
  INV_X1    g0236(.A(G77), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n261), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n272), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT11), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n440), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n283), .A2(new_n231), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT12), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n433), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n424), .A2(G200), .ZN(new_n449));
  OAI211_X1 g0249(.A(G190), .B(new_n421), .C1(new_n428), .C2(new_n429), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(new_n446), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n331), .A2(new_n415), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(G41), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n208), .B(G45), .C1(new_n458), .C2(KEYINPUT5), .ZN(new_n461));
  OAI211_X1 g0261(.A(G257), .B(new_n307), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n457), .A2(KEYINPUT84), .A3(new_n459), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT84), .B1(new_n457), .B2(new_n459), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G274), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n305), .B2(new_n306), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT82), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n456), .A2(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT82), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n467), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n462), .B1(new_n465), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n461), .A2(new_n468), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n471), .A2(KEYINPUT82), .A3(new_n472), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n467), .C1(new_n464), .C2(new_n463), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n462), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT4), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1698), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(G244), .C1(new_n292), .C2(new_n291), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n296), .A2(KEYINPUT80), .A3(G244), .A4(new_n485), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G244), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n288), .B2(new_n289), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT4), .B1(new_n492), .B2(new_n286), .ZN(new_n493));
  OAI211_X1 g0293(.A(G250), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n494));
  INV_X1    g0294(.A(G283), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n259), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n490), .A2(new_n499), .A3(KEYINPUT81), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n290), .B2(G250), .ZN(new_n501));
  OAI211_X1 g0301(.A(G244), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n484), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n501), .A2(new_n488), .A3(new_n503), .A4(new_n489), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT81), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n500), .A2(new_n506), .A3(new_n300), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n483), .A2(new_n507), .A3(new_n314), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n260), .A2(new_n437), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n510));
  XOR2_X1   g0310(.A(G97), .B(G107), .Z(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n512), .B2(G20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n341), .A2(G107), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n346), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n259), .A2(G1), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n280), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n204), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n279), .A2(G97), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n307), .B1(new_n504), .B2(new_n505), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n476), .A2(new_n482), .B1(new_n523), .B2(new_n500), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n508), .B(new_n522), .C1(G169), .C2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n483), .A2(new_n507), .A3(G190), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n521), .C1(new_n317), .C2(new_n524), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT86), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT86), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n471), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT87), .B1(new_n302), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT87), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n467), .A2(new_n535), .A3(new_n471), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n491), .A2(G1698), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(G238), .B2(G1698), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n540), .B2(new_n293), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n300), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n307), .A2(new_n533), .A3(G250), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n537), .A2(new_n542), .A3(new_n544), .A4(G190), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT89), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n541), .B2(new_n300), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(KEYINPUT89), .A3(G190), .A4(new_n537), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT90), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT19), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n209), .B1(new_n416), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(G87), .B2(new_n206), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n209), .B(G68), .C1(new_n291), .C2(new_n292), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n553), .B1(new_n261), .B2(new_n204), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n272), .B1(new_n283), .B2(new_n397), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT88), .B1(new_n517), .B2(G87), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT88), .ZN(new_n561));
  INV_X1    g0361(.A(G87), .ZN(new_n562));
  NOR4_X1   g0362(.A1(new_n280), .A2(new_n561), .A3(new_n562), .A4(new_n516), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n559), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n317), .B1(new_n548), .B2(new_n537), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n547), .A2(KEYINPUT90), .A3(new_n549), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n552), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n548), .A2(new_n537), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n381), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n559), .B1(new_n397), .B2(new_n518), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n571), .C1(G179), .C2(new_n569), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT91), .B1(new_n532), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT86), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT86), .B1(new_n525), .B2(new_n527), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT91), .B(new_n574), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(G20), .B1(G33), .B2(G283), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n259), .A2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(G116), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n581), .A2(new_n582), .B1(G20), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n272), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n586), .A2(KEYINPUT92), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(KEYINPUT92), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n516), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n346), .A2(G116), .A3(new_n279), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n283), .A2(new_n583), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n272), .A2(new_n584), .A3(KEYINPUT92), .A4(new_n586), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n589), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n595));
  OAI211_X1 g0395(.A(G257), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n288), .A2(G303), .A3(new_n289), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n300), .ZN(new_n599));
  OAI211_X1 g0399(.A(G270), .B(new_n307), .C1(new_n460), .C2(new_n461), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n480), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n601), .A2(KEYINPUT21), .A3(G169), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n314), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n594), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G264), .B(new_n307), .C1(new_n460), .C2(new_n461), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n606));
  OAI211_X1 g0406(.A(G250), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G33), .A2(G294), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n300), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n480), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n381), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n480), .A2(new_n314), .A3(new_n610), .A4(new_n605), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n209), .B(G87), .C1(new_n291), .C2(new_n292), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT22), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT22), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n296), .A2(new_n616), .A3(new_n209), .A4(G87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT23), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n209), .B2(G107), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT24), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT24), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n618), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n346), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n517), .A2(G107), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n279), .A2(G107), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT25), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n612), .B(new_n613), .C1(new_n630), .C2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n594), .A2(new_n601), .A3(G169), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n636), .A2(KEYINPUT93), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT93), .B1(new_n636), .B2(new_n637), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n604), .B(new_n635), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  AOI211_X1 g0440(.A(KEYINPUT24), .B(new_n624), .C1(new_n615), .C2(new_n617), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n628), .B1(new_n618), .B2(new_n625), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n272), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n634), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n611), .A2(G200), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n480), .A2(new_n610), .A3(G190), .A4(new_n605), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n643), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n601), .A2(G200), .ZN(new_n648));
  INV_X1    g0448(.A(new_n594), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n648), .B(new_n649), .C1(new_n354), .C2(new_n601), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NOR4_X1   g0451(.A1(new_n454), .A2(new_n580), .A3(new_n640), .A4(new_n651), .ZN(G372));
  INV_X1    g0452(.A(new_n414), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n433), .A2(new_n447), .B1(new_n451), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n379), .A2(new_n393), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n391), .B(new_n387), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n327), .A2(new_n329), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n315), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n573), .B2(new_n525), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n566), .A2(new_n550), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n660), .A2(new_n572), .A3(new_n647), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n640), .A2(new_n661), .A3(new_n525), .A4(new_n527), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n572), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n483), .A2(new_n507), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n521), .B1(new_n665), .B2(new_n381), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n664), .A2(new_n666), .A3(new_n667), .A4(new_n508), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n659), .A2(new_n662), .A3(new_n572), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n658), .B1(new_n454), .B2(new_n670), .ZN(G369));
  OR2_X1    g0471(.A1(new_n638), .A2(new_n639), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n604), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n649), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n673), .B(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n650), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n635), .A2(new_n679), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n679), .B1(new_n630), .B2(new_n634), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n647), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n686), .B1(new_n635), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n679), .B1(new_n672), .B2(new_n604), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n689), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n686), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT94), .ZN(G399));
  INV_X1    g0496(.A(new_n227), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n233), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n640), .A2(new_n651), .A3(new_n679), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n575), .B2(new_n579), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n569), .A2(new_n601), .A3(new_n314), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT97), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n665), .A2(new_n611), .ZN(new_n709));
  AND4_X1   g0509(.A1(new_n537), .A2(new_n548), .A3(new_n605), .A4(new_n610), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n483), .A2(new_n507), .A3(new_n710), .A4(new_n603), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT96), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n708), .A2(new_n709), .B1(new_n712), .B2(KEYINPUT30), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n712), .A2(KEYINPUT30), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n680), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n704), .B1(new_n706), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  INV_X1    g0521(.A(new_n525), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n574), .A2(new_n667), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT26), .B1(new_n525), .B2(new_n663), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n572), .B(KEYINPUT98), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n662), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n721), .B1(new_n728), .B2(new_n680), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n669), .A2(new_n680), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n720), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n703), .B1(new_n732), .B2(G1), .ZN(G364));
  INV_X1    g0533(.A(KEYINPUT99), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n684), .B(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n209), .A2(G13), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n208), .B1(new_n737), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n698), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n736), .B(new_n741), .C1(G330), .C2(new_n683), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n227), .A2(new_n296), .ZN(new_n743));
  INV_X1    g0543(.A(G355), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n744), .B1(G116), .B2(new_n227), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n252), .A2(G45), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n697), .A2(new_n296), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n470), .B2(new_n234), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n745), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n235), .B1(G20), .B2(new_n381), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n740), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n209), .A2(new_n314), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT100), .Z(new_n759));
  NOR2_X1   g0559(.A1(G190), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n209), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n760), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT101), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n762), .A2(G311), .B1(G329), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n296), .B1(new_n768), .B2(G303), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n354), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n759), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n766), .B(new_n769), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n758), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n354), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n771), .A2(new_n314), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n775), .A2(G326), .B1(new_n777), .B2(G294), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n774), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(G317), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n763), .A2(new_n354), .A3(G200), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n778), .B(new_n783), .C1(new_n495), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n767), .A2(new_n562), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n296), .B1(new_n784), .B2(new_n205), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(G50), .C2(new_n775), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n788), .B1(new_n437), .B2(new_n761), .C1(new_n334), .C2(new_n772), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n764), .A2(new_n332), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  INV_X1    g0591(.A(new_n779), .ZN(new_n792));
  INV_X1    g0592(.A(new_n777), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n791), .B1(new_n231), .B2(new_n792), .C1(new_n204), .C2(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n773), .A2(new_n785), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n757), .B1(new_n754), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT102), .Z(new_n797));
  INV_X1    g0597(.A(new_n753), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n683), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n742), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  INV_X1    g0601(.A(new_n720), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT108), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n414), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n402), .A2(new_n679), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(new_n410), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n653), .A2(new_n679), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n730), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n804), .A2(new_n410), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n669), .A2(new_n680), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n802), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n740), .B1(new_n802), .B2(new_n812), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n754), .A2(new_n751), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT103), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n740), .B1(new_n817), .B2(G77), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G137), .A2(new_n775), .B1(new_n779), .B2(G150), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT106), .Z(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n772), .C1(new_n332), .C2(new_n761), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT34), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n793), .A2(new_n334), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n296), .B1(new_n767), .B2(new_n281), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n784), .A2(new_n231), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  INV_X1    g0628(.A(new_n765), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n823), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n775), .ZN(new_n831));
  INV_X1    g0631(.A(G303), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n832), .B1(new_n784), .B2(new_n562), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n583), .A2(new_n761), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n833), .B(new_n835), .C1(G283), .C2(new_n779), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n772), .A2(new_n837), .B1(new_n204), .B2(new_n793), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT105), .Z(new_n839));
  OAI21_X1  g0639(.A(new_n293), .B1(new_n767), .B2(new_n205), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT104), .Z(new_n841));
  NAND3_X1  g0641(.A1(new_n836), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n830), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n818), .B1(new_n843), .B2(new_n754), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT107), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n808), .A2(new_n751), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n814), .A2(new_n815), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  OR2_X1    g0648(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(G116), .A3(new_n236), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT36), .Z(new_n852));
  OAI211_X1 g0652(.A(new_n234), .B(G77), .C1(new_n231), .C2(new_n334), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n281), .A2(G68), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n208), .B(G13), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n448), .A2(new_n679), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT110), .ZN(new_n858));
  INV_X1    g0658(.A(new_n336), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n349), .A2(new_n343), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n341), .A2(KEYINPUT77), .A3(G68), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(KEYINPUT16), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n345), .A2(new_n272), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n376), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n677), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n394), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n865), .A2(new_n866), .B1(new_n389), .B2(new_n373), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n865), .A2(new_n385), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT109), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n380), .A2(new_n385), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT109), .B1(new_n389), .B2(new_n390), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT37), .B1(new_n389), .B2(new_n373), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n380), .A2(new_n866), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n869), .B(KEYINPUT38), .C1(new_n873), .C2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n346), .B1(new_n862), .B2(KEYINPUT16), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n336), .B1(new_n342), .B2(new_n344), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n351), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n388), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n377), .B1(new_n886), .B2(new_n677), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n390), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n879), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n890), .B2(new_n869), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n858), .B(KEYINPUT39), .C1(new_n882), .C2(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(KEYINPUT111), .B(KEYINPUT38), .Z(new_n893));
  OAI21_X1  g0693(.A(new_n377), .B1(new_n389), .B2(new_n390), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n389), .A2(new_n677), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT112), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(new_n879), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n394), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n897), .B1(new_n896), .B2(new_n879), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n893), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(new_n881), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n892), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n871), .A2(new_n872), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n875), .A2(new_n876), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n877), .A2(new_n878), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n907), .A2(KEYINPUT37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n869), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n881), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n858), .B1(new_n913), .B2(KEYINPUT39), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n857), .B1(new_n905), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT113), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n866), .B1(new_n387), .B2(new_n391), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n804), .A2(new_n679), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n811), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n447), .A2(new_n679), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n448), .A2(new_n451), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n451), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n447), .B(new_n679), .C1(new_n922), .C2(new_n433), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n917), .B1(new_n926), .B2(new_n913), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n915), .A2(new_n916), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n916), .B1(new_n915), .B2(new_n927), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n453), .B1(new_n729), .B2(new_n731), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n658), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n931), .B(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n808), .B1(new_n921), .B2(new_n923), .ZN(new_n935));
  INV_X1    g0735(.A(new_n705), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT91), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n936), .B1(new_n939), .B2(new_n578), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n715), .B2(new_n716), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n935), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n913), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n943), .A2(KEYINPUT40), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n896), .A2(new_n879), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT112), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n899), .A3(new_n898), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n882), .B1(new_n948), .B2(new_n893), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT40), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n940), .A2(new_n942), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n454), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n704), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n951), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n934), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n208), .B2(new_n737), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n934), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n856), .B1(new_n957), .B2(new_n958), .ZN(G367));
  OAI221_X1 g0759(.A(new_n755), .B1(new_n227), .B2(new_n397), .C1(new_n748), .C2(new_n247), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n740), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n293), .B1(new_n764), .B2(new_n780), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G107), .B2(new_n777), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n772), .B2(new_n832), .C1(new_n495), .C2(new_n761), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT116), .B1(new_n768), .B2(G116), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT46), .Z(new_n966));
  INV_X1    g0766(.A(new_n784), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n775), .A2(G311), .B1(new_n967), .B2(G97), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n837), .B2(new_n792), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n964), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n793), .A2(new_n231), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G143), .B2(new_n775), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n258), .B2(new_n772), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT117), .Z(new_n974));
  INV_X1    g0774(.A(G137), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n296), .B1(new_n764), .B2(new_n975), .C1(new_n334), .C2(new_n767), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n792), .A2(new_n332), .B1(new_n784), .B2(new_n437), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(new_n762), .C2(G50), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n970), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n961), .B1(new_n980), .B2(new_n754), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n564), .A2(new_n679), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n664), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n572), .A2(new_n982), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT114), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(KEYINPUT114), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n981), .B1(new_n798), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n691), .A2(new_n689), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n693), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT115), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n684), .B(new_n990), .C1(new_n734), .C2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n735), .A2(KEYINPUT115), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(new_n993), .B2(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n732), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n722), .A2(new_n679), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n525), .B(new_n527), .C1(new_n521), .C2(new_n680), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n694), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT45), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n694), .A2(new_n998), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT44), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1000), .A2(new_n690), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n690), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n732), .B1(new_n995), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n698), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n739), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n997), .A2(new_n635), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n679), .B1(new_n1011), .B2(new_n525), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n693), .A2(new_n998), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(KEYINPUT42), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(KEYINPUT42), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1014), .A2(new_n1015), .B1(KEYINPUT43), .B2(new_n987), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n690), .B1(new_n997), .B2(new_n996), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n988), .B1(new_n1010), .B2(new_n1020), .ZN(G387));
  NOR2_X1   g0821(.A1(new_n994), .A2(new_n732), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n995), .A2(new_n698), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(KEYINPUT119), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT119), .B2(new_n1023), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n743), .A2(new_n700), .B1(G107), .B2(new_n227), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n244), .A2(new_n470), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n700), .ZN(new_n1028));
  AOI211_X1 g0828(.A(G45), .B(new_n1028), .C1(G68), .C2(G77), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n398), .A2(G50), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n748), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1026), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n740), .B1(new_n1033), .B2(new_n756), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n767), .A2(new_n437), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n793), .A2(new_n397), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(G159), .C2(new_n775), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n266), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n762), .A2(G68), .B1(new_n1038), .B2(new_n779), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n296), .B1(new_n764), .B2(new_n258), .C1(new_n204), .C2(new_n784), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n772), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(G50), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1037), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n764), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n296), .B1(new_n1044), .B2(G326), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n793), .A2(new_n495), .B1(new_n767), .B2(new_n837), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G311), .A2(new_n779), .B1(new_n775), .B2(G322), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n772), .B2(new_n780), .C1(new_n832), .C2(new_n761), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1045), .B1(new_n583), .B2(new_n784), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1034), .B1(new_n1055), .B2(new_n754), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n689), .B2(new_n798), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT118), .Z(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n994), .B2(new_n739), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1025), .A2(new_n1059), .ZN(G393));
  OAI21_X1  g0860(.A(new_n698), .B1(new_n995), .B2(new_n1006), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1005), .B1(new_n732), .B2(new_n994), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n755), .B1(new_n204), .B2(new_n227), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n747), .B2(new_n255), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n772), .A2(new_n332), .B1(new_n258), .B2(new_n831), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  AOI22_X1  g0867(.A1(new_n779), .A2(G50), .B1(new_n777), .B2(G77), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n231), .B2(new_n767), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n761), .A2(new_n398), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n296), .B1(new_n764), .B2(new_n821), .C1(new_n562), .C2(new_n784), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT120), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT120), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n772), .A2(new_n834), .B1(new_n780), .B2(new_n831), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT121), .B(KEYINPUT52), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n792), .A2(new_n832), .B1(new_n793), .B2(new_n583), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G283), .B2(new_n768), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n293), .B1(new_n764), .B2(new_n770), .C1(new_n205), .C2(new_n784), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n762), .B2(G294), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1073), .A2(new_n1074), .A3(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n741), .B(new_n1065), .C1(new_n1083), .C2(new_n754), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n998), .B2(new_n798), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1006), .B2(new_n738), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1063), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G390));
  INV_X1    g0888(.A(new_n942), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n704), .B1(new_n1089), .B2(new_n706), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n808), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n715), .A2(new_n716), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n715), .B2(KEYINPUT31), .ZN(new_n1093));
  OAI211_X1 g0893(.A(G330), .B(new_n1091), .C1(new_n940), .C2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n921), .A2(new_n923), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n935), .A2(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n919), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n924), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n680), .B(new_n810), .C1(new_n726), .C2(new_n727), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1099), .A2(new_n918), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1096), .A2(new_n1097), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n935), .B(G330), .C1(new_n940), .C2(new_n942), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n857), .B1(new_n919), .B2(new_n924), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n905), .A2(new_n914), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1095), .B1(new_n1099), .B2(new_n918), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1107), .A2(new_n949), .A3(new_n857), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1104), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n857), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n925), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT39), .B1(new_n882), .B2(new_n891), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT110), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1111), .A2(new_n1113), .A3(new_n904), .A4(new_n892), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n949), .A2(new_n857), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n720), .A2(new_n1091), .A3(new_n924), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1090), .A2(new_n453), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n932), .A3(new_n658), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1102), .A2(new_n1109), .A3(new_n1118), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n924), .B1(new_n720), .B2(new_n1091), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n919), .B1(new_n1124), .B2(new_n1104), .ZN(new_n1125));
  OAI21_X1  g0925(.A(G330), .B1(new_n940), .B2(new_n942), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1095), .B1(new_n1126), .B2(new_n808), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1117), .A2(new_n1127), .A3(new_n1100), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1120), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT122), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1129), .A2(new_n1130), .A3(new_n1118), .A4(new_n1109), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n1131), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1103), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1132), .B(new_n698), .C1(new_n1135), .C2(new_n1129), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n739), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n740), .B1(new_n817), .B2(new_n1038), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n792), .A2(new_n205), .B1(new_n831), .B2(new_n495), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n826), .B(new_n1139), .C1(G77), .C2(new_n777), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n296), .B(new_n786), .C1(new_n1041), .C2(G116), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n765), .A2(G294), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n762), .A2(G97), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n767), .A2(KEYINPUT53), .A3(new_n258), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT53), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n768), .B2(G150), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT54), .B(G143), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1145), .B(new_n1147), .C1(new_n762), .C2(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n792), .A2(new_n975), .B1(new_n793), .B2(new_n332), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G128), .B2(new_n775), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1041), .A2(G132), .B1(G125), .B2(new_n765), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n296), .B1(new_n784), .B2(new_n281), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT123), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1144), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1138), .B1(new_n1157), .B2(new_n754), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1113), .A2(new_n904), .A3(new_n892), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n752), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1136), .A2(new_n1137), .A3(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(KEYINPUT124), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n318), .A2(new_n677), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n331), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n331), .A2(new_n1163), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1167), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n929), .B2(new_n930), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n915), .A2(new_n927), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT113), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(new_n928), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n951), .A2(G330), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1171), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1178), .A2(new_n1179), .A3(new_n738), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1170), .A2(new_n751), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n754), .A2(G50), .A3(new_n751), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1041), .A2(G107), .B1(G283), .B2(new_n765), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n293), .A2(new_n458), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n971), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(new_n397), .C2(new_n761), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n784), .A2(new_n334), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n792), .A2(new_n204), .B1(new_n831), .B2(new_n583), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1186), .A2(new_n1035), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G128), .A2(new_n1041), .B1(new_n762), .B2(G137), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n775), .A2(G125), .B1(new_n777), .B2(G150), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n779), .A2(G132), .B1(new_n768), .B2(new_n1149), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n967), .A2(G159), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n1044), .C2(G124), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1184), .B(new_n281), .C1(G33), .C2(G41), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1190), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n741), .B(new_n1182), .C1(new_n1202), .C2(new_n754), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1181), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1162), .B1(new_n1180), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1179), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1171), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n739), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(KEYINPUT124), .A3(new_n1204), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1122), .A2(KEYINPUT122), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1130), .B1(new_n1135), .B2(new_n1129), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1121), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(KEYINPUT125), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT125), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1132), .A2(new_n1216), .A3(new_n1121), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT57), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT57), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1178), .A2(new_n1179), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1216), .B1(new_n1132), .B2(new_n1121), .ZN(new_n1223));
  AOI211_X1 g1023(.A(KEYINPUT125), .B(new_n1120), .C1(new_n1123), .C2(new_n1131), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n698), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1211), .B1(new_n1220), .B2(new_n1226), .ZN(G375));
  NAND2_X1  g1027(.A1(new_n1102), .A2(new_n739), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n740), .B1(new_n817), .B2(G68), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n293), .B(new_n1187), .C1(new_n1041), .C2(G137), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G132), .A2(new_n775), .B1(new_n779), .B2(new_n1149), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G159), .A2(new_n768), .B1(new_n777), .B2(G50), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n762), .A2(G150), .B1(G128), .B2(new_n765), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n767), .A2(new_n204), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1235), .B(new_n1036), .C1(G294), .C2(new_n775), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n293), .B1(new_n784), .B2(new_n437), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n765), .B2(G303), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1236), .B(new_n1238), .C1(new_n495), .C2(new_n772), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n761), .A2(new_n205), .B1(new_n583), .B2(new_n792), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT126), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1234), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1229), .B1(new_n1242), .B2(new_n754), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n924), .B2(new_n752), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1228), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1102), .A2(new_n1121), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1102), .A2(new_n1121), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1009), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1247), .B2(new_n1249), .ZN(G381));
  AOI21_X1  g1050(.A(new_n699), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1219), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1221), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1251), .A2(new_n1253), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1254));
  INV_X1    g1054(.A(G378), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1025), .A2(new_n800), .A3(new_n1059), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G384), .A2(new_n1257), .A3(G390), .A4(G387), .ZN(new_n1258));
  OR3_X1    g1058(.A1(new_n1256), .A2(new_n1258), .A3(G381), .ZN(G407));
  OAI211_X1 g1059(.A(G407), .B(G213), .C1(G343), .C2(new_n1256), .ZN(G409));
  NAND3_X1  g1060(.A1(new_n1247), .A2(KEYINPUT60), .A3(new_n1248), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n698), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1247), .B1(KEYINPUT60), .B2(new_n1248), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1246), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1264), .A2(new_n847), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n847), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G213), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(G343), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(G2897), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1267), .B(new_n1270), .Z(new_n1271));
  OAI211_X1 g1071(.A(G378), .B(new_n1211), .C1(new_n1220), .C2(new_n1226), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1180), .A2(new_n1205), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1252), .B2(new_n1008), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1255), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1269), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1271), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1218), .A2(new_n1009), .A3(new_n1219), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G378), .B1(new_n1279), .B2(new_n1273), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1254), .B2(G378), .ZN(new_n1281));
  OAI21_X1  g1081(.A(KEYINPUT127), .B1(new_n1281), .B2(new_n1269), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  OR2_X1    g1083(.A1(G387), .A2(new_n1087), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G387), .A2(new_n1087), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1257), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1284), .A2(new_n1257), .A3(new_n1287), .A4(new_n1285), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1269), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1267), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1292), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1276), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1283), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1276), .A2(new_n1301), .A3(new_n1295), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1290), .B1(new_n1276), .B2(new_n1271), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1301), .B1(new_n1276), .B2(new_n1295), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1300), .B1(new_n1305), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1108(.A1(G375), .A2(new_n1255), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1272), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1295), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1309), .A2(new_n1272), .A3(new_n1267), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1313), .B(new_n1306), .ZN(G402));
endmodule


