//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n468), .B1(new_n461), .B2(new_n462), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G113), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n461), .A2(new_n462), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n463), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(KEYINPUT69), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n489), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n464), .C1(new_n491), .C2(new_n492), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n478), .A2(new_n500), .A3(G138), .A4(new_n464), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G50), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n511), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(new_n509), .A3(KEYINPUT5), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n505), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n507), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n517), .A2(new_n520), .ZN(G166));
  XNOR2_X1  g096(.A(new_n515), .B(KEYINPUT71), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n506), .A2(G51), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n516), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n523), .A2(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(new_n506), .A2(G52), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n532), .B2(new_n516), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n510), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n513), .B1(KEYINPUT5), .B2(new_n509), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n511), .A2(KEYINPUT70), .A3(G543), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT71), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n534), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n533), .B1(new_n544), .B2(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT72), .ZN(G171));
  AOI22_X1  g121(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n519), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n515), .A2(new_n505), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT73), .B(G43), .Z(new_n550));
  AOI22_X1  g125(.A1(new_n549), .A2(G81), .B1(new_n506), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n506), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n549), .A2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n515), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n519), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n559), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n568), .A2(new_n569), .B1(G91), .B2(new_n549), .ZN(new_n570));
  INV_X1    g145(.A(new_n566), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(KEYINPUT74), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n545), .B(new_n575), .ZN(G301));
  OR2_X1    g151(.A1(new_n523), .A2(new_n529), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND3_X1  g153(.A1(new_n515), .A2(G87), .A3(new_n505), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(G74), .B1(new_n539), .B2(new_n541), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n519), .ZN(G288));
  NAND2_X1  g158(.A1(new_n512), .A2(new_n514), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n584), .A2(G86), .A3(new_n535), .A4(new_n505), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n505), .A2(G48), .A3(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n515), .B2(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n588), .B1(new_n592), .B2(new_n519), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  AOI211_X1 g169(.A(new_n594), .B(new_n510), .C1(new_n512), .C2(new_n514), .ZN(new_n595));
  OAI211_X1 g170(.A(KEYINPUT76), .B(G651), .C1(new_n595), .C2(new_n591), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n587), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n542), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n519), .B1(new_n601), .B2(KEYINPUT77), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(KEYINPUT77), .B2(new_n601), .ZN(new_n603));
  XNOR2_X1  g178(.A(KEYINPUT78), .B(G85), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n549), .A2(new_n604), .B1(G47), .B2(new_n506), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(new_n506), .A2(G54), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT81), .B(G66), .Z(new_n608));
  AOI22_X1  g183(.A1(new_n515), .A2(new_n608), .B1(G79), .B2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n519), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n549), .A2(G92), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(KEYINPUT80), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(KEYINPUT79), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G171), .ZN(new_n621));
  NAND3_X1  g196(.A1(G301), .A2(KEYINPUT79), .A3(G868), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n621), .A2(new_n622), .ZN(G284));
  XNOR2_X1  g198(.A(G284), .B(KEYINPUT82), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n573), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n573), .B2(G868), .ZN(G280));
  AND2_X1   g202(.A1(new_n616), .A2(new_n617), .ZN(new_n628));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND3_X1  g205(.A1(new_n616), .A2(new_n629), .A3(new_n617), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n478), .A2(new_n466), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n463), .A2(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n464), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(G123), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n642), .B1(new_n643), .B2(new_n644), .C1(new_n645), .C2(new_n479), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(G156));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n665), .B1(new_n667), .B2(KEYINPUT84), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(KEYINPUT84), .B2(new_n667), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n666), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n665), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n669), .B(new_n671), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n671), .A2(new_n666), .A3(new_n674), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n674), .A3(new_n670), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n689), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n690), .A2(KEYINPUT20), .A3(new_n689), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n691), .B1(new_n689), .B2(new_n687), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(G35), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n485), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT29), .ZN(new_n706));
  INV_X1    g281(.A(G2090), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT95), .Z(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G19), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n553), .B2(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G1341), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n463), .A2(G140), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n716));
  INV_X1    g291(.A(G116), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(G2105), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n480), .B2(G128), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G29), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT89), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n703), .A2(G26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT90), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G2067), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n709), .A2(new_n712), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G21), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G286), .B2(G16), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT92), .B(G1966), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G1341), .B2(new_n711), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT31), .B(G11), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n646), .A2(new_n703), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT30), .B(G28), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n738), .B(new_n739), .C1(new_n703), .C2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n703), .B1(KEYINPUT24), .B2(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(KEYINPUT24), .B2(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n476), .B2(G29), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n703), .A2(G32), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  INV_X1    g323(.A(G129), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n479), .B2(new_n749), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n463), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(G29), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n741), .B1(new_n742), .B2(new_n745), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n733), .A2(new_n734), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n754), .A2(new_n755), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT91), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n745), .A2(new_n742), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT94), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n707), .B2(new_n706), .ZN(new_n763));
  NOR2_X1   g338(.A1(G27), .A2(G29), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G164), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2078), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n703), .A2(G33), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n491), .A2(new_n492), .ZN(new_n769));
  INV_X1    g344(.A(G127), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G2105), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT25), .ZN(new_n773));
  NAND2_X1  g348(.A1(G103), .A2(G2104), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G2105), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n463), .A2(G139), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n767), .B1(new_n778), .B2(new_n703), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2072), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n766), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n758), .A2(new_n760), .A3(new_n763), .A4(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n729), .A2(new_n737), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n628), .B2(G16), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(G1348), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(G1348), .ZN(new_n787));
  NAND2_X1  g362(.A1(G299), .A2(G16), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n730), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT23), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n788), .A2(G1956), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(G1956), .B1(new_n788), .B2(new_n790), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n786), .B(new_n787), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1961), .Z(new_n797));
  NAND3_X1  g372(.A1(new_n783), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n730), .A2(G24), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n603), .A2(new_n605), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n730), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(G1986), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(G1986), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n463), .A2(G131), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n464), .A2(G107), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(G119), .ZN(new_n809));
  OAI221_X1 g384(.A(new_n806), .B1(new_n807), .B2(new_n808), .C1(new_n809), .C2(new_n479), .ZN(new_n810));
  MUX2_X1   g385(.A(G25), .B(new_n810), .S(G29), .Z(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n804), .A2(new_n805), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n730), .A2(G6), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n597), .B2(new_n730), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G23), .B(G288), .S(G16), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT33), .B(G1976), .Z(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n730), .A2(G22), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G166), .B2(new_n730), .ZN(new_n824));
  INV_X1    g399(.A(G1971), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n820), .A2(new_n821), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n819), .A2(new_n822), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n815), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT87), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n831), .B(new_n833), .Z(new_n834));
  OR2_X1    g409(.A1(new_n832), .A2(KEYINPUT87), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n799), .A2(new_n800), .B1(new_n834), .B2(new_n835), .ZN(G311));
  NAND2_X1  g411(.A1(new_n799), .A2(new_n800), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(G150));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n628), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n519), .ZN(new_n845));
  INV_X1    g420(.A(new_n506), .ZN(new_n846));
  INV_X1    g421(.A(G55), .ZN(new_n847));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n846), .A2(new_n847), .B1(new_n516), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n845), .A2(KEYINPUT97), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT97), .B1(new_n845), .B2(new_n849), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(new_n553), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n553), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n843), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n842), .B(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n856), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n840), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n856), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n843), .A2(new_n857), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT39), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT99), .B(G860), .Z(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n845), .A2(new_n849), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n866), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(G145));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n778), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n753), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n503), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n503), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n720), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n874), .A2(new_n503), .ZN(new_n879));
  INV_X1    g454(.A(new_n720), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n875), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n810), .B(new_n637), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n463), .A2(G142), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT101), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G118), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n885), .A2(new_n886), .B1(new_n888), .B2(G2105), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n480), .A2(G130), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n882), .B(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n878), .A2(new_n881), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n878), .B2(new_n881), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(KEYINPUT103), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n878), .A2(new_n881), .A3(new_n896), .A4(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n646), .B(new_n476), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n485), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n878), .A2(new_n881), .ZN(new_n902));
  INV_X1    g477(.A(new_n892), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n900), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n905), .A3(new_n893), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n908), .A3(KEYINPUT104), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n905), .B1(new_n895), .B2(new_n897), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n907), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n631), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n616), .A2(KEYINPUT105), .A3(new_n629), .A4(new_n617), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n854), .B2(new_n855), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n618), .A2(new_n573), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n616), .A2(new_n567), .A3(new_n572), .A4(new_n617), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n852), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n552), .B1(new_n924), .B2(new_n850), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(new_n853), .A3(new_n917), .A4(new_n918), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n920), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  INV_X1    g503(.A(new_n922), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n617), .A2(new_n616), .B1(new_n567), .B2(new_n572), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n922), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n920), .A2(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(G288), .B(G166), .Z(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G290), .A2(new_n597), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(G290), .A2(new_n597), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n939), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n935), .A3(new_n937), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n942), .A3(KEYINPUT106), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n940), .A2(new_n942), .A3(KEYINPUT106), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n934), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n944), .B(new_n946), .C1(new_n927), .C2(new_n933), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(G868), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n868), .A2(G868), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n619), .B1(new_n948), .B2(new_n949), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT107), .B1(new_n956), .B2(new_n953), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(G295));
  NAND2_X1  g533(.A1(new_n951), .A2(new_n954), .ZN(G331));
  NAND2_X1  g534(.A1(new_n931), .A2(new_n932), .ZN(new_n960));
  NAND2_X1  g535(.A1(G301), .A2(G168), .ZN(new_n961));
  NAND2_X1  g536(.A1(G171), .A2(G286), .ZN(new_n962));
  AND4_X1   g537(.A1(new_n853), .A2(new_n925), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n853), .A2(new_n925), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n962), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n854), .B2(new_n855), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n925), .A2(new_n853), .A3(new_n961), .A4(new_n962), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n923), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n940), .A2(new_n942), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G37), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n965), .A2(new_n971), .A3(new_n969), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n977), .A3(new_n974), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n970), .A2(new_n972), .ZN(new_n981));
  AND4_X1   g556(.A1(new_n977), .A2(new_n981), .A3(new_n907), .A4(new_n974), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n973), .B2(new_n974), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n497), .B2(new_n502), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n467), .A2(new_n475), .A3(G40), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(G1976), .B(new_n581), .C1(new_n582), .C2(new_n519), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(KEYINPUT109), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n992), .A3(G288), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n991), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n584), .A2(G61), .A3(new_n535), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n589), .B(KEYINPUT75), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n519), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(G1981), .B1(new_n1001), .B2(new_n587), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT110), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(G1981), .C1(new_n1001), .C2(new_n587), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(G1981), .B(new_n587), .C1(new_n593), .C2(new_n596), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n998), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1981), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n597), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(KEYINPUT49), .A3(new_n1005), .A4(new_n1003), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1008), .A2(new_n1011), .A3(new_n989), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT114), .B1(new_n997), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1008), .A2(new_n1011), .A3(new_n989), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1014), .B(new_n1015), .C1(new_n996), .C2(new_n995), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n503), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n467), .A2(new_n475), .A3(G40), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1020), .A2(G1384), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n503), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1971), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1019), .A2(KEYINPUT50), .ZN(new_n1027));
  NOR2_X1   g602(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1022), .B1(new_n503), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n707), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n986), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G166), .A2(new_n986), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(KEYINPUT108), .A2(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1034), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1037), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n503), .A2(new_n1028), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1040), .B(new_n988), .C1(new_n1041), .C2(new_n987), .ZN(new_n1042));
  AOI21_X1  g617(.A(G2090), .B1(new_n1042), .B2(KEYINPUT112), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1027), .A2(new_n1044), .A3(new_n1029), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1025), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g623(.A(KEYINPUT113), .B(new_n1025), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1039), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n503), .A2(new_n1023), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n988), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n503), .B2(new_n1018), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n734), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1027), .A2(new_n742), .A3(new_n1029), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n986), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1056), .A2(G168), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1017), .A2(new_n1038), .A3(new_n1050), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT115), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1038), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1042), .A2(KEYINPUT112), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n707), .A3(new_n1045), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1026), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT113), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(G8), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1067), .B2(new_n1039), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n1017), .A4(new_n1057), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1059), .A2(new_n1060), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1057), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1072), .A2(new_n1061), .A3(new_n1060), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n995), .A2(new_n996), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1014), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n997), .A2(new_n1012), .A3(KEYINPUT111), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1071), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1017), .A2(new_n1038), .A3(new_n1050), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1056), .A2(G286), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1054), .A2(G168), .A3(new_n1055), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(G8), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(KEYINPUT120), .A3(KEYINPUT51), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1084), .A2(KEYINPUT120), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(G8), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(KEYINPUT120), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1081), .B(new_n1085), .C1(new_n1086), .C2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1091));
  INV_X1    g666(.A(G2078), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT53), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G171), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT121), .B(G1961), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n467), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n467), .A2(new_n1097), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1092), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1098), .A2(new_n475), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n503), .B2(new_n1023), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1096), .B1(new_n1021), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1094), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1092), .A2(KEYINPUT53), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1052), .A2(new_n1053), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT122), .B1(new_n1106), .B2(new_n1096), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1095), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1042), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1021), .A2(KEYINPUT53), .A3(new_n1092), .A4(new_n1024), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1093), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1104), .B1(G301), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1094), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1093), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n1103), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1115), .B1(new_n1119), .B2(G171), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1114), .A2(new_n1115), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1080), .A2(KEYINPUT124), .A3(new_n1090), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n1123));
  AOI21_X1  g698(.A(G301), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1118), .A2(G301), .A3(new_n1103), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1115), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1120), .A2(new_n1117), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1090), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1017), .A2(new_n1038), .A3(new_n1050), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1123), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(KEYINPUT57), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n570), .A2(new_n571), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(KEYINPUT57), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  INV_X1    g711(.A(G1956), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1091), .A2(new_n1136), .B1(new_n1042), .B2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n987), .A2(new_n988), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(G2067), .ZN(new_n1141));
  INV_X1    g716(.A(G1348), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n1042), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1139), .B1(new_n618), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT117), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1135), .A2(new_n1147), .A3(new_n1138), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(KEYINPUT118), .A3(new_n618), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n618), .B(KEYINPUT118), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1152), .B(new_n1153), .C1(new_n1154), .C2(new_n1151), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1139), .A2(KEYINPUT61), .A3(new_n1145), .ZN(new_n1156));
  INV_X1    g731(.A(G1996), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1091), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT58), .B(G1341), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n1140), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n552), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT59), .Z(new_n1162));
  NAND3_X1  g737(.A1(new_n1155), .A2(new_n1156), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1149), .A2(KEYINPUT61), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1150), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1122), .A2(new_n1130), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1061), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1012), .A2(G1976), .A3(G288), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n989), .B1(new_n1168), .B2(new_n1007), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1129), .B1(KEYINPUT62), .B2(new_n1090), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1090), .A2(KEYINPUT62), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1124), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1079), .A2(new_n1166), .A3(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n720), .B(new_n727), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n753), .B(new_n1157), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n810), .A2(new_n813), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n810), .A2(new_n813), .ZN(new_n1181));
  AND4_X1   g756(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(G1986), .B2(G290), .ZN(new_n1183));
  AND2_X1   g758(.A1(G290), .A2(G1986), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1177), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1176), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1177), .ZN(new_n1187));
  INV_X1    g762(.A(new_n753), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1187), .B1(new_n1188), .B2(new_n1178), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT125), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1177), .A2(new_n1157), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT46), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g768(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT127), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1193), .B(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1197));
  INV_X1    g772(.A(G1986), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n802), .A2(new_n1198), .A3(new_n1177), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1200), .B2(KEYINPUT48), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(KEYINPUT48), .B2(new_n1200), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1203), .A2(new_n1180), .B1(G2067), .B2(new_n720), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1177), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1196), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1186), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g783(.A(G319), .B(new_n681), .C1(new_n662), .C2(new_n663), .ZN(new_n1210));
  NOR2_X1   g784(.A1(G229), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g785(.A(new_n914), .B(new_n1211), .C1(new_n982), .C2(new_n983), .ZN(G225));
  INV_X1    g786(.A(G225), .ZN(G308));
endmodule


