

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(n740), .B(n739), .ZN(n745) );
  INV_X1 U550 ( .A(KEYINPUT29), .ZN(n739) );
  NAND2_X1 U551 ( .A1(n745), .A2(n744), .ZN(n756) );
  NOR2_X1 U552 ( .A1(G651), .A2(G543), .ZN(n638) );
  AND2_X1 U553 ( .A1(n729), .A2(n728), .ZN(n514) );
  OR2_X1 U554 ( .A1(n514), .A2(n734), .ZN(n735) );
  INV_X1 U555 ( .A(KEYINPUT31), .ZN(n752) );
  XNOR2_X1 U556 ( .A(n752), .B(KEYINPUT90), .ZN(n753) );
  XNOR2_X1 U557 ( .A(n754), .B(n753), .ZN(n755) );
  AND2_X1 U558 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X2 U559 ( .A1(n710), .A2(n709), .ZN(n741) );
  NOR2_X1 U560 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n708) );
  INV_X1 U562 ( .A(G651), .ZN(n529) );
  NOR2_X1 U563 ( .A1(G651), .A2(n628), .ZN(n634) );
  XOR2_X1 U564 ( .A(n591), .B(KEYINPUT15), .Z(n994) );
  XNOR2_X1 U565 ( .A(KEYINPUT1), .B(n526), .ZN(n635) );
  XNOR2_X1 U566 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n516) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  XNOR2_X1 U568 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X2 U569 ( .A(KEYINPUT64), .B(n517), .ZN(n873) );
  NAND2_X1 U570 ( .A1(G138), .A2(n873), .ZN(n519) );
  INV_X1 U571 ( .A(G2105), .ZN(n520) );
  AND2_X1 U572 ( .A1(n520), .A2(G2104), .ZN(n872) );
  NAND2_X1 U573 ( .A1(n872), .A2(G102), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n519), .A2(n518), .ZN(n524) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n876) );
  NAND2_X1 U576 ( .A1(G114), .A2(n876), .ZN(n522) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n520), .ZN(n877) );
  NAND2_X1 U578 ( .A1(G126), .A2(n877), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n524), .A2(n523), .ZN(G164) );
  NAND2_X1 U581 ( .A1(G85), .A2(n638), .ZN(n528) );
  NOR2_X1 U582 ( .A1(G543), .A2(n529), .ZN(n525) );
  XOR2_X1 U583 ( .A(KEYINPUT66), .B(n525), .Z(n526) );
  NAND2_X1 U584 ( .A1(G60), .A2(n635), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n628) );
  NOR2_X1 U587 ( .A1(n628), .A2(n529), .ZN(n631) );
  NAND2_X1 U588 ( .A1(G72), .A2(n631), .ZN(n531) );
  NAND2_X1 U589 ( .A1(G47), .A2(n634), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n531), .A2(n530), .ZN(n532) );
  OR2_X1 U591 ( .A1(n533), .A2(n532), .ZN(G290) );
  XNOR2_X1 U592 ( .A(G2454), .B(G2443), .ZN(n543) );
  XOR2_X1 U593 ( .A(KEYINPUT98), .B(G2430), .Z(n535) );
  XNOR2_X1 U594 ( .A(G2446), .B(KEYINPUT99), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n535), .B(n534), .ZN(n539) );
  XOR2_X1 U596 ( .A(G2451), .B(G2427), .Z(n537) );
  INV_X1 U597 ( .A(G1341), .ZN(n1004) );
  XOR2_X1 U598 ( .A(G1348), .B(n1004), .Z(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U600 ( .A(n539), .B(n538), .Z(n541) );
  XNOR2_X1 U601 ( .A(G2435), .B(G2438), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n543), .B(n542), .ZN(n544) );
  AND2_X1 U604 ( .A1(n544), .A2(G14), .ZN(G401) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U606 ( .A1(n876), .A2(G111), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G135), .A2(n873), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n877), .A2(G123), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT18), .B(n547), .Z(n548) );
  NOR2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n872), .A2(G99), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n915) );
  XNOR2_X1 U614 ( .A(G2096), .B(n915), .ZN(n552) );
  OR2_X1 U615 ( .A1(G2100), .A2(n552), .ZN(G156) );
  NAND2_X1 U616 ( .A1(n638), .A2(G89), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U618 ( .A1(G76), .A2(n631), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n556), .B(KEYINPUT5), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n634), .A2(G51), .ZN(n558) );
  NAND2_X1 U622 ( .A1(G63), .A2(n635), .ZN(n557) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n559), .Z(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n563) );
  XOR2_X1 U629 ( .A(n563), .B(KEYINPUT10), .Z(n906) );
  NAND2_X1 U630 ( .A1(n906), .A2(G567), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U632 ( .A1(G43), .A2(n634), .ZN(n575) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n566) );
  NAND2_X1 U634 ( .A1(G56), .A2(n635), .ZN(n565) );
  XNOR2_X1 U635 ( .A(n566), .B(n565), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n638), .A2(G81), .ZN(n567) );
  XNOR2_X1 U637 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U638 ( .A1(G68), .A2(n631), .ZN(n568) );
  NAND2_X1 U639 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U640 ( .A(KEYINPUT13), .B(n570), .Z(n571) );
  NOR2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U642 ( .A(KEYINPUT71), .B(n573), .Z(n574) );
  AND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n1005) );
  NAND2_X1 U644 ( .A1(n1005), .A2(G860), .ZN(G153) );
  NAND2_X1 U645 ( .A1(n634), .A2(G52), .ZN(n576) );
  XNOR2_X1 U646 ( .A(KEYINPUT67), .B(n576), .ZN(n582) );
  NAND2_X1 U647 ( .A1(G90), .A2(n638), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G77), .A2(n631), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U650 ( .A(KEYINPUT68), .B(n579), .Z(n580) );
  XNOR2_X1 U651 ( .A(KEYINPUT9), .B(n580), .ZN(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G64), .A2(n635), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U656 ( .A1(n634), .A2(G54), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G66), .A2(n635), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G92), .A2(n638), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G79), .A2(n631), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U663 ( .A(n994), .ZN(n733) );
  INV_X1 U664 ( .A(G868), .ZN(n605) );
  NAND2_X1 U665 ( .A1(n733), .A2(n605), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G91), .A2(n638), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G78), .A2(n631), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n634), .A2(G53), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G65), .A2(n635), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n728) );
  INV_X1 U674 ( .A(n728), .ZN(G299) );
  NOR2_X1 U675 ( .A1(G286), .A2(n605), .ZN(n601) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U677 ( .A1(n601), .A2(n600), .ZN(G297) );
  INV_X1 U678 ( .A(G860), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n603), .A2(n994), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U682 ( .A1(n1005), .A2(n605), .ZN(n606) );
  XOR2_X1 U683 ( .A(KEYINPUT72), .B(n606), .Z(n609) );
  NAND2_X1 U684 ( .A1(G868), .A2(n994), .ZN(n607) );
  NOR2_X1 U685 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U687 ( .A1(n634), .A2(G55), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G67), .A2(n635), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G93), .A2(n638), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G80), .A2(n631), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n648) );
  NAND2_X1 U694 ( .A1(n994), .A2(G559), .ZN(n653) );
  XOR2_X1 U695 ( .A(n1005), .B(n653), .Z(n616) );
  NOR2_X1 U696 ( .A1(G860), .A2(n616), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n648), .B(n617), .ZN(G145) );
  NAND2_X1 U698 ( .A1(G88), .A2(n638), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G75), .A2(n631), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n634), .A2(G50), .ZN(n621) );
  NAND2_X1 U702 ( .A1(G62), .A2(n635), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n623), .A2(n622), .ZN(G166) );
  NAND2_X1 U705 ( .A1(G49), .A2(n634), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U708 ( .A(KEYINPUT73), .B(n626), .Z(n627) );
  NOR2_X1 U709 ( .A1(n635), .A2(n627), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(G288) );
  XOR2_X1 U712 ( .A(KEYINPUT2), .B(KEYINPUT75), .Z(n633) );
  NAND2_X1 U713 ( .A1(G73), .A2(n631), .ZN(n632) );
  XNOR2_X1 U714 ( .A(n633), .B(n632), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n634), .A2(G48), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G61), .A2(n635), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n638), .A2(G86), .ZN(n639) );
  XOR2_X1 U719 ( .A(KEYINPUT74), .B(n639), .Z(n640) );
  NOR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(G305) );
  NOR2_X1 U722 ( .A1(G868), .A2(n648), .ZN(n644) );
  XNOR2_X1 U723 ( .A(n644), .B(KEYINPUT77), .ZN(n656) );
  XNOR2_X1 U724 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n646) );
  XOR2_X1 U725 ( .A(G288), .B(G299), .Z(n645) );
  XNOR2_X1 U726 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n648), .B(n647), .ZN(n650) );
  XNOR2_X1 U728 ( .A(G305), .B(n1005), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U730 ( .A(G166), .B(n651), .Z(n652) );
  XNOR2_X1 U731 ( .A(G290), .B(n652), .ZN(n894) );
  XNOR2_X1 U732 ( .A(n894), .B(n653), .ZN(n654) );
  NAND2_X1 U733 ( .A1(G868), .A2(n654), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n656), .A2(n655), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n658), .ZN(n659) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n660), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U740 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U741 ( .A(KEYINPUT78), .B(G44), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n661), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U743 ( .A1(G108), .A2(G120), .ZN(n662) );
  NOR2_X1 U744 ( .A1(G237), .A2(n662), .ZN(n663) );
  NAND2_X1 U745 ( .A1(G69), .A2(n663), .ZN(n826) );
  NAND2_X1 U746 ( .A1(n826), .A2(G567), .ZN(n670) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(KEYINPUT79), .Z(n665) );
  NAND2_X1 U748 ( .A1(G132), .A2(G82), .ZN(n664) );
  XNOR2_X1 U749 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U750 ( .A1(n666), .A2(G218), .ZN(n667) );
  NAND2_X1 U751 ( .A1(G96), .A2(n667), .ZN(n668) );
  XNOR2_X1 U752 ( .A(KEYINPUT80), .B(n668), .ZN(n827) );
  NAND2_X1 U753 ( .A1(n827), .A2(G2106), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n670), .A2(n669), .ZN(n905) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n671) );
  NOR2_X1 U756 ( .A1(n905), .A2(n671), .ZN(n825) );
  NAND2_X1 U757 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U758 ( .A1(G137), .A2(n873), .ZN(n674) );
  NAND2_X1 U759 ( .A1(G101), .A2(n872), .ZN(n672) );
  XOR2_X1 U760 ( .A(KEYINPUT23), .B(n672), .Z(n673) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n678) );
  NAND2_X1 U762 ( .A1(G113), .A2(n876), .ZN(n676) );
  NAND2_X1 U763 ( .A1(G125), .A2(n877), .ZN(n675) );
  NAND2_X1 U764 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U765 ( .A1(n678), .A2(n677), .ZN(G160) );
  INV_X1 U766 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U767 ( .A(KEYINPUT81), .B(G166), .ZN(G303) );
  NAND2_X1 U768 ( .A1(G117), .A2(n876), .ZN(n680) );
  NAND2_X1 U769 ( .A1(G129), .A2(n877), .ZN(n679) );
  NAND2_X1 U770 ( .A1(n680), .A2(n679), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n872), .A2(G105), .ZN(n681) );
  XOR2_X1 U772 ( .A(KEYINPUT38), .B(n681), .Z(n682) );
  NOR2_X1 U773 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U774 ( .A(n684), .B(KEYINPUT84), .ZN(n686) );
  NAND2_X1 U775 ( .A1(G141), .A2(n873), .ZN(n685) );
  NAND2_X1 U776 ( .A1(n686), .A2(n685), .ZN(n890) );
  NAND2_X1 U777 ( .A1(G1996), .A2(n890), .ZN(n687) );
  XOR2_X1 U778 ( .A(KEYINPUT85), .B(n687), .Z(n695) );
  NAND2_X1 U779 ( .A1(n876), .A2(G107), .ZN(n689) );
  NAND2_X1 U780 ( .A1(G131), .A2(n873), .ZN(n688) );
  NAND2_X1 U781 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U782 ( .A1(G95), .A2(n872), .ZN(n691) );
  NAND2_X1 U783 ( .A1(G119), .A2(n877), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n869) );
  NAND2_X1 U786 ( .A1(G1991), .A2(n869), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n918) );
  NAND2_X1 U788 ( .A1(G160), .A2(G40), .ZN(n709) );
  NOR2_X1 U789 ( .A1(n708), .A2(n709), .ZN(n817) );
  NAND2_X1 U790 ( .A1(n918), .A2(n817), .ZN(n696) );
  XOR2_X1 U791 ( .A(KEYINPUT86), .B(n696), .Z(n809) );
  NAND2_X1 U792 ( .A1(n872), .A2(G104), .ZN(n698) );
  NAND2_X1 U793 ( .A1(G140), .A2(n873), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U795 ( .A(KEYINPUT34), .B(n699), .ZN(n705) );
  NAND2_X1 U796 ( .A1(G116), .A2(n876), .ZN(n701) );
  NAND2_X1 U797 ( .A1(G128), .A2(n877), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U799 ( .A(KEYINPUT35), .B(n702), .Z(n703) );
  XNOR2_X1 U800 ( .A(KEYINPUT82), .B(n703), .ZN(n704) );
  NOR2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U802 ( .A(n706), .B(KEYINPUT36), .Z(n707) );
  XNOR2_X1 U803 ( .A(KEYINPUT83), .B(n707), .ZN(n891) );
  XNOR2_X1 U804 ( .A(KEYINPUT37), .B(G2067), .ZN(n814) );
  NOR2_X1 U805 ( .A1(n891), .A2(n814), .ZN(n912) );
  NAND2_X1 U806 ( .A1(n817), .A2(n912), .ZN(n812) );
  XOR2_X1 U807 ( .A(G1981), .B(G305), .Z(n986) );
  INV_X1 U808 ( .A(n708), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n741), .A2(G2072), .ZN(n711) );
  XNOR2_X1 U810 ( .A(n711), .B(KEYINPUT27), .ZN(n713) );
  INV_X1 U811 ( .A(G1956), .ZN(n836) );
  NOR2_X1 U812 ( .A1(n836), .A2(n741), .ZN(n712) );
  NOR2_X1 U813 ( .A1(n713), .A2(n712), .ZN(n729) );
  NOR2_X1 U814 ( .A1(n729), .A2(n728), .ZN(n714) );
  XOR2_X1 U815 ( .A(n714), .B(KEYINPUT28), .Z(n738) );
  XNOR2_X1 U816 ( .A(G1996), .B(KEYINPUT88), .ZN(n938) );
  NAND2_X1 U817 ( .A1(n938), .A2(n741), .ZN(n716) );
  XOR2_X1 U818 ( .A(KEYINPUT26), .B(KEYINPUT89), .Z(n721) );
  INV_X1 U819 ( .A(n721), .ZN(n715) );
  NAND2_X1 U820 ( .A1(n716), .A2(n715), .ZN(n720) );
  INV_X1 U821 ( .A(n741), .ZN(n757) );
  NAND2_X1 U822 ( .A1(G1348), .A2(n733), .ZN(n717) );
  NAND2_X1 U823 ( .A1(n1004), .A2(n717), .ZN(n718) );
  NAND2_X1 U824 ( .A1(n757), .A2(n718), .ZN(n719) );
  NAND2_X1 U825 ( .A1(n720), .A2(n719), .ZN(n727) );
  NAND2_X1 U826 ( .A1(n721), .A2(n938), .ZN(n723) );
  NAND2_X1 U827 ( .A1(G2067), .A2(n733), .ZN(n722) );
  NAND2_X1 U828 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U829 ( .A1(n724), .A2(n741), .ZN(n725) );
  NAND2_X1 U830 ( .A1(n725), .A2(n1005), .ZN(n726) );
  NOR2_X1 U831 ( .A1(n727), .A2(n726), .ZN(n736) );
  NAND2_X1 U832 ( .A1(G1348), .A2(n757), .ZN(n731) );
  NAND2_X1 U833 ( .A1(G2067), .A2(n741), .ZN(n730) );
  NAND2_X1 U834 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U835 ( .A1(n733), .A2(n732), .ZN(n734) );
  OR2_X1 U836 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U837 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U838 ( .A(G1961), .B(KEYINPUT87), .ZN(n962) );
  NAND2_X1 U839 ( .A1(n757), .A2(n962), .ZN(n743) );
  XNOR2_X1 U840 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NAND2_X1 U841 ( .A1(n741), .A2(n943), .ZN(n742) );
  NAND2_X1 U842 ( .A1(n743), .A2(n742), .ZN(n746) );
  NAND2_X1 U843 ( .A1(n746), .A2(G171), .ZN(n744) );
  NOR2_X1 U844 ( .A1(G171), .A2(n746), .ZN(n751) );
  NAND2_X1 U845 ( .A1(G8), .A2(n757), .ZN(n796) );
  NOR2_X1 U846 ( .A1(G1966), .A2(n796), .ZN(n771) );
  NOR2_X1 U847 ( .A1(G2084), .A2(n757), .ZN(n768) );
  NOR2_X1 U848 ( .A1(n771), .A2(n768), .ZN(n747) );
  NAND2_X1 U849 ( .A1(G8), .A2(n747), .ZN(n748) );
  XNOR2_X1 U850 ( .A(KEYINPUT30), .B(n748), .ZN(n749) );
  NOR2_X1 U851 ( .A1(G168), .A2(n749), .ZN(n750) );
  NOR2_X1 U852 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U853 ( .A1(n756), .A2(n755), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n769), .A2(G286), .ZN(n766) );
  INV_X1 U855 ( .A(G8), .ZN(n764) );
  NOR2_X1 U856 ( .A1(G1971), .A2(n796), .ZN(n759) );
  NOR2_X1 U857 ( .A1(G2090), .A2(n757), .ZN(n758) );
  NOR2_X1 U858 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U859 ( .A(KEYINPUT91), .B(n760), .Z(n761) );
  NAND2_X1 U860 ( .A1(n761), .A2(G303), .ZN(n762) );
  XNOR2_X1 U861 ( .A(n762), .B(KEYINPUT92), .ZN(n763) );
  OR2_X1 U862 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U863 ( .A(n767), .B(KEYINPUT32), .ZN(n775) );
  NAND2_X1 U864 ( .A1(G8), .A2(n768), .ZN(n773) );
  INV_X1 U865 ( .A(n769), .ZN(n770) );
  NOR2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n794) );
  NOR2_X1 U869 ( .A1(G1976), .A2(G288), .ZN(n783) );
  NOR2_X1 U870 ( .A1(G1971), .A2(G303), .ZN(n776) );
  NOR2_X1 U871 ( .A1(n783), .A2(n776), .ZN(n998) );
  NAND2_X1 U872 ( .A1(n794), .A2(n998), .ZN(n778) );
  AND2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  NOR2_X1 U874 ( .A1(n1000), .A2(n796), .ZN(n777) );
  NAND2_X1 U875 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U876 ( .A1(KEYINPUT93), .A2(n779), .ZN(n780) );
  NOR2_X1 U877 ( .A1(KEYINPUT33), .A2(n780), .ZN(n788) );
  INV_X1 U878 ( .A(KEYINPUT93), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n783), .A2(KEYINPUT33), .ZN(n781) );
  NAND2_X1 U880 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U881 ( .A1(n783), .A2(KEYINPUT93), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U883 ( .A1(n796), .A2(n786), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n986), .A2(n789), .ZN(n801) );
  NOR2_X1 U885 ( .A1(G1981), .A2(G305), .ZN(n790) );
  XOR2_X1 U886 ( .A(n790), .B(KEYINPUT24), .Z(n791) );
  NOR2_X1 U887 ( .A1(n796), .A2(n791), .ZN(n799) );
  NOR2_X1 U888 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U889 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U892 ( .A(KEYINPUT94), .B(n797), .Z(n798) );
  NOR2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n812), .A2(n802), .ZN(n803) );
  NOR2_X1 U896 ( .A1(n809), .A2(n803), .ZN(n805) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U898 ( .A1(n990), .A2(n817), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n820) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n890), .ZN(n909) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n869), .ZN(n914) );
  NOR2_X1 U903 ( .A1(n806), .A2(n914), .ZN(n807) );
  XOR2_X1 U904 ( .A(KEYINPUT95), .B(n807), .Z(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n909), .A2(n810), .ZN(n811) );
  XNOR2_X1 U907 ( .A(KEYINPUT39), .B(n811), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n814), .A2(n891), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(KEYINPUT96), .ZN(n925) );
  NAND2_X1 U911 ( .A1(n816), .A2(n925), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n822) );
  XOR2_X1 U914 ( .A(KEYINPUT97), .B(KEYINPUT40), .Z(n821) );
  XNOR2_X1 U915 ( .A(n822), .B(n821), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n906), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U918 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U922 ( .A(G132), .ZN(G219) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G82), .ZN(G220) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XOR2_X1 U930 ( .A(G2100), .B(G2096), .Z(n829) );
  XNOR2_X1 U931 ( .A(KEYINPUT42), .B(G2678), .ZN(n828) );
  XNOR2_X1 U932 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U933 ( .A(KEYINPUT43), .B(G2090), .Z(n831) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U935 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U936 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U937 ( .A(G2084), .B(G2078), .ZN(n834) );
  XNOR2_X1 U938 ( .A(n835), .B(n834), .ZN(G227) );
  XNOR2_X1 U939 ( .A(n836), .B(G1961), .ZN(n838) );
  XNOR2_X1 U940 ( .A(G1976), .B(G1971), .ZN(n837) );
  XNOR2_X1 U941 ( .A(n838), .B(n837), .ZN(n848) );
  XOR2_X1 U942 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n840) );
  XNOR2_X1 U943 ( .A(G1991), .B(KEYINPUT41), .ZN(n839) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U945 ( .A(G1966), .B(G1981), .Z(n842) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1986), .ZN(n841) );
  XNOR2_X1 U947 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U948 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U949 ( .A(KEYINPUT100), .B(G2474), .ZN(n845) );
  XNOR2_X1 U950 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U952 ( .A1(n872), .A2(G100), .ZN(n849) );
  XOR2_X1 U953 ( .A(KEYINPUT103), .B(n849), .Z(n851) );
  NAND2_X1 U954 ( .A1(n876), .A2(G112), .ZN(n850) );
  NAND2_X1 U955 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U956 ( .A(KEYINPUT104), .B(n852), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G124), .A2(n877), .ZN(n853) );
  XNOR2_X1 U958 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U959 ( .A1(G136), .A2(n873), .ZN(n854) );
  NAND2_X1 U960 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U961 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U962 ( .A1(G118), .A2(n876), .ZN(n859) );
  NAND2_X1 U963 ( .A1(G130), .A2(n877), .ZN(n858) );
  NAND2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n872), .A2(G106), .ZN(n861) );
  NAND2_X1 U966 ( .A1(G142), .A2(n873), .ZN(n860) );
  NAND2_X1 U967 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U968 ( .A(n862), .B(KEYINPUT45), .Z(n863) );
  NOR2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n865), .B(n915), .ZN(n888) );
  XOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT106), .Z(n867) );
  XNOR2_X1 U972 ( .A(G162), .B(KEYINPUT108), .ZN(n866) );
  XNOR2_X1 U973 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U974 ( .A(KEYINPUT48), .B(n868), .ZN(n871) );
  XNOR2_X1 U975 ( .A(n869), .B(KEYINPUT105), .ZN(n870) );
  XNOR2_X1 U976 ( .A(n871), .B(n870), .ZN(n884) );
  NAND2_X1 U977 ( .A1(n872), .A2(G103), .ZN(n875) );
  NAND2_X1 U978 ( .A1(G139), .A2(n873), .ZN(n874) );
  NAND2_X1 U979 ( .A1(n875), .A2(n874), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G115), .A2(n876), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G127), .A2(n877), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U985 ( .A(KEYINPUT107), .B(n883), .Z(n921) );
  XOR2_X1 U986 ( .A(n884), .B(n921), .Z(n886) );
  XNOR2_X1 U987 ( .A(G164), .B(G160), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U989 ( .A(n888), .B(n887), .Z(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n892) );
  XOR2_X1 U991 ( .A(n892), .B(n891), .Z(n893) );
  NOR2_X1 U992 ( .A1(G37), .A2(n893), .ZN(G395) );
  XOR2_X1 U993 ( .A(n894), .B(G286), .Z(n896) );
  XOR2_X1 U994 ( .A(G301), .B(n994), .Z(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U996 ( .A1(G37), .A2(n897), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U998 ( .A(KEYINPUT110), .B(KEYINPUT49), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G401), .A2(n905), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(KEYINPUT109), .B(n900), .ZN(n901) );
  NOR2_X1 U1002 ( .A1(n902), .A2(n901), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(n905), .ZN(G319) );
  INV_X1 U1007 ( .A(n906), .ZN(G223) );
  XNOR2_X1 U1008 ( .A(G2090), .B(G162), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n907), .B(KEYINPUT111), .ZN(n908) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(KEYINPUT51), .B(n910), .ZN(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n920) );
  XOR2_X1 U1013 ( .A(G160), .B(G2084), .Z(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n928) );
  XOR2_X1 U1018 ( .A(G2072), .B(n921), .Z(n923) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(KEYINPUT50), .B(n924), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(KEYINPUT52), .B(n929), .ZN(n930) );
  XOR2_X1 U1025 ( .A(KEYINPUT55), .B(KEYINPUT112), .Z(n952) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n952), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n931), .A2(G29), .ZN(n1019) );
  XNOR2_X1 U1028 ( .A(KEYINPUT113), .B(G2090), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(G35), .ZN(n951) );
  XOR2_X1 U1030 ( .A(G34), .B(KEYINPUT115), .Z(n934) );
  XNOR2_X1 U1031 ( .A(G2084), .B(KEYINPUT54), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(n934), .B(n933), .ZN(n949) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(G33), .B(G2072), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1036 ( .A(G1991), .B(G25), .Z(n937) );
  NAND2_X1 U1037 ( .A1(n937), .A2(G28), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(G32), .B(n938), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1041 ( .A(G27), .B(n943), .Z(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT53), .B(n946), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT114), .B(n947), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n953), .B(n952), .ZN(n955) );
  XOR2_X1 U1048 ( .A(G29), .B(KEYINPUT116), .Z(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n956), .A2(G11), .ZN(n1017) );
  XOR2_X1 U1051 ( .A(G16), .B(KEYINPUT120), .Z(n985) );
  XOR2_X1 U1052 ( .A(G1986), .B(G24), .Z(n958) );
  XOR2_X1 U1053 ( .A(G1971), .B(G22), .Z(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G23), .B(G1976), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT58), .B(n961), .Z(n982) );
  XOR2_X1 U1058 ( .A(n962), .B(G5), .Z(n979) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G21), .ZN(n976) );
  XOR2_X1 U1060 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n974) );
  XOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT59), .Z(n963) );
  XNOR2_X1 U1062 ( .A(G4), .B(n963), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT121), .B(G20), .ZN(n964) );
  XOR2_X1 U1064 ( .A(n964), .B(G1956), .Z(n969) );
  XNOR2_X1 U1065 ( .A(G1981), .B(G6), .ZN(n966) );
  XOR2_X1 U1066 ( .A(G19), .B(n1004), .Z(n965) );
  NOR2_X1 U1067 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1068 ( .A(KEYINPUT122), .B(n967), .Z(n968) );
  NOR2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1070 ( .A(n970), .B(KEYINPUT123), .ZN(n971) );
  NOR2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1072 ( .A(n974), .B(n973), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(KEYINPUT125), .B(n977), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1076 ( .A(KEYINPUT126), .B(n980), .Z(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(KEYINPUT61), .B(n983), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n1014) );
  XNOR2_X1 U1080 ( .A(KEYINPUT56), .B(G16), .ZN(n1011) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G168), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(n988), .B(KEYINPUT57), .ZN(n1009) );
  XOR2_X1 U1084 ( .A(G301), .B(G1961), .Z(n993) );
  XOR2_X1 U1085 ( .A(G299), .B(G1956), .Z(n989) );
  XNOR2_X1 U1086 ( .A(n989), .B(KEYINPUT117), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n996) );
  XOR2_X1 U1089 ( .A(G1348), .B(n994), .Z(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(G1971), .A2(G303), .ZN(n997) );
  NAND2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(n1001), .B(KEYINPUT118), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1005), .B(n1004), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(KEYINPUT119), .B(n1012), .Z(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1015), .Z(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1020), .ZN(G150) );
  INV_X1 U1106 ( .A(G150), .ZN(G311) );
endmodule

