//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT96), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT15), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  NOR3_X1   g015(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT92), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(new_n218), .B2(new_n217), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n220), .A2(KEYINPUT93), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(KEYINPUT93), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n211), .B(new_n215), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT90), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n217), .B1(new_n224), .B2(new_n216), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(new_n224), .B2(new_n216), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n211), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT15), .A3(new_n212), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(KEYINPUT17), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT95), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT94), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n223), .A2(new_n231), .A3(new_n228), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n223), .B2(new_n228), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR4_X1   g035(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT95), .A4(KEYINPUT17), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n210), .B(new_n229), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n232), .A2(new_n233), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT97), .B1(new_n239), .B2(new_n210), .ZN(new_n240));
  OR4_X1    g039(.A1(KEYINPUT97), .A2(new_n232), .A3(new_n233), .A4(new_n210), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT98), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G169gat), .B(G197gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT12), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n244), .A2(new_n245), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n238), .A2(new_n242), .A3(KEYINPUT18), .A4(new_n243), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n210), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n243), .B(KEYINPUT13), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n255), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n244), .A2(new_n245), .B1(new_n258), .B2(new_n259), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n263), .B(new_n256), .C1(new_n246), .C2(new_n253), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G232gat), .A2(G233gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT41), .ZN(new_n268));
  XNOR2_X1  g067(.A(G134gat), .B(G162gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G85gat), .A2(G92gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT7), .ZN(new_n273));
  NAND2_X1  g072(.A1(G99gat), .A2(G106gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT8), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n273), .B(new_n275), .C1(G85gat), .C2(G92gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G99gat), .B(G106gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT101), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n229), .B(new_n279), .C1(new_n236), .C2(new_n237), .ZN(new_n280));
  XOR2_X1   g079(.A(G190gat), .B(G218gat), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n234), .A2(new_n278), .B1(KEYINPUT41), .B2(new_n267), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n282), .B1(new_n280), .B2(new_n283), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n271), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n286), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n270), .A3(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291));
  XOR2_X1   g090(.A(G57gat), .B(G64gat), .Z(new_n292));
  INV_X1    g091(.A(KEYINPUT9), .ZN(new_n293));
  INV_X1    g092(.A(G71gat), .ZN(new_n294));
  INV_X1    g093(.A(G78gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G71gat), .B(G78gat), .Z(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n210), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT100), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n291), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT99), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n301), .B(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G127gat), .B(G155gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G183gat), .B(G211gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n309), .B(new_n310), .Z(new_n311));
  AND2_X1   g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n306), .A2(new_n311), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n299), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n278), .A2(KEYINPUT10), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n278), .B(new_n319), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(KEYINPUT10), .ZN(new_n322));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n323), .B(KEYINPUT102), .Z(new_n324));
  AND2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n323), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n318), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n323), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n327), .A3(new_n317), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n290), .A2(new_n314), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n266), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n338));
  INV_X1    g137(.A(G134gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G127gat), .ZN(new_n340));
  INV_X1    g139(.A(G127gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G134gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT68), .ZN(new_n343));
  OR3_X1    g142(.A1(new_n341), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G120gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G113gat), .ZN(new_n347));
  INV_X1    g146(.A(G113gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G120gat), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT1), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n338), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n349), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n354), .A2(KEYINPUT69), .A3(new_n343), .A4(new_n344), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G141gat), .B(G148gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G155gat), .ZN(new_n359));
  INV_X1    g158(.A(G162gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(KEYINPUT2), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n358), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n362), .B(new_n361), .C1(new_n357), .C2(KEYINPUT2), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n340), .A2(new_n342), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT70), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT70), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n350), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n356), .A2(new_n368), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n368), .B1(new_n356), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n337), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n356), .A2(new_n368), .A3(new_n374), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n356), .A2(new_n374), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n365), .A2(new_n366), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n367), .A2(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n351), .A2(new_n355), .B1(new_n371), .B2(new_n373), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(new_n368), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n381), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n378), .B(new_n379), .C1(new_n390), .C2(new_n337), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n382), .A2(new_n367), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n380), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n394), .B2(new_n337), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n385), .A2(new_n384), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n380), .B(KEYINPUT4), .C1(new_n396), .C2(new_n388), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n375), .A2(new_n387), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n337), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n399), .B2(KEYINPUT81), .ZN(new_n400));
  XOR2_X1   g199(.A(G1gat), .B(G29gat), .Z(new_n401));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n400), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT6), .B1(new_n411), .B2(new_n405), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n407), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT83), .B(KEYINPUT6), .C1(new_n411), .C2(new_n405), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n417), .A2(KEYINPUT77), .ZN(new_n418));
  NAND2_X1  g217(.A1(G211gat), .A2(G218gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT22), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(KEYINPUT77), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G197gat), .B(G204gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT78), .ZN(new_n424));
  XOR2_X1   g223(.A(G211gat), .B(G218gat), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n426), .B1(new_n423), .B2(new_n424), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT25), .ZN(new_n432));
  AND2_X1   g231(.A1(G169gat), .A2(G176gat), .ZN(new_n433));
  INV_X1    g232(.A(G169gat), .ZN(new_n434));
  INV_X1    g233(.A(G176gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT23), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G183gat), .A2(G190gat), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT24), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G183gat), .ZN(new_n442));
  INV_X1    g241(.A(G190gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(G169gat), .A2(G176gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT23), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT64), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n438), .A2(new_n446), .A3(new_n448), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G169gat), .A2(G176gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n437), .B1(G169gat), .B2(G176gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n449), .A2(KEYINPUT25), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n439), .A2(new_n461), .A3(new_n440), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n439), .B2(new_n440), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n444), .B(new_n445), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n432), .A2(new_n452), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n442), .A2(KEYINPUT27), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G183gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n468), .A3(new_n443), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n469), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT28), .B1(new_n469), .B2(KEYINPUT67), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT26), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n453), .B1(new_n447), .B2(new_n472), .ZN(new_n473));
  NOR3_X1   g272(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n439), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n470), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n452), .A2(new_n432), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n469), .A2(KEYINPUT67), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT28), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n473), .A2(new_n474), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n484), .A2(new_n439), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT79), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n431), .B1(new_n478), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n431), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(KEYINPUT29), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n430), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n490), .A3(new_n493), .ZN(new_n496));
  INV_X1    g295(.A(new_n430), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n492), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  XOR2_X1   g298(.A(G8gat), .B(G36gat), .Z(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT80), .ZN(new_n501));
  XNOR2_X1  g300(.A(G64gat), .B(G92gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n495), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n495), .B2(new_n499), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n506));
  OR3_X1    g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n495), .A2(new_n499), .ZN(new_n508));
  INV_X1    g307(.A(new_n503), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n508), .A2(KEYINPUT30), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n416), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT71), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n465), .B2(new_n476), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n481), .A2(KEYINPUT71), .A3(new_n487), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n382), .ZN(new_n517));
  INV_X1    g316(.A(G227gat), .ZN(new_n518));
  INV_X1    g317(.A(G233gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n488), .A2(new_n514), .A3(new_n388), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT32), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g324(.A(G71gat), .B(G99gat), .Z(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G43gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(KEYINPUT33), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n522), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n523), .A2(new_n525), .A3(new_n537), .A4(new_n528), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n530), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n521), .ZN(new_n540));
  INV_X1    g339(.A(new_n520), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n539), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT75), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n530), .A2(new_n536), .A3(new_n545), .A4(new_n538), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT75), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n539), .A2(new_n550), .A3(new_n546), .ZN(new_n551));
  XNOR2_X1  g350(.A(G78gat), .B(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G22gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n384), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n428), .B2(new_n429), .ZN(new_n557));
  NAND2_X1  g356(.A1(G228gat), .A2(G233gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n423), .A2(new_n426), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT29), .B1(new_n423), .B2(new_n426), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT3), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n557), .B(new_n558), .C1(new_n368), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n422), .A2(new_n421), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n417), .A2(KEYINPUT77), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n424), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n425), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n566), .A2(new_n427), .B1(new_n384), .B2(new_n555), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n555), .A3(new_n427), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n383), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n569), .B2(new_n367), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n554), .B(new_n562), .C1(new_n570), .C2(new_n558), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT84), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n368), .B1(new_n568), .B2(new_n383), .ZN(new_n573));
  OAI211_X1 g372(.A(G228gat), .B(G233gat), .C1(new_n573), .C2(new_n567), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n554), .B1(new_n574), .B2(new_n562), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n553), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n562), .B1(new_n570), .B2(new_n558), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G22gat), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n578), .A2(KEYINPUT84), .A3(new_n571), .A4(new_n552), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT31), .B(G50gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n576), .A2(new_n579), .A3(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n548), .A2(new_n549), .A3(new_n551), .A4(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT35), .B1(new_n513), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n549), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT76), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n539), .A2(new_n589), .A3(new_n546), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n507), .A2(KEYINPUT86), .A3(new_n511), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT86), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n594), .B2(new_n510), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n409), .B1(new_n407), .B2(new_n412), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT35), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(new_n585), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n587), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n548), .A2(KEYINPUT36), .A3(new_n549), .A4(new_n551), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n591), .B2(KEYINPUT36), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT85), .ZN(new_n603));
  INV_X1    g402(.A(new_n584), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n581), .B1(new_n576), .B2(new_n579), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n583), .A2(KEYINPUT85), .A3(new_n584), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n513), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT39), .B1(new_n394), .B2(new_n337), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n337), .B2(new_n390), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT87), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n397), .A2(new_n398), .A3(new_n613), .A4(new_n337), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n614), .B2(new_n405), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n612), .A3(new_n405), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT88), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT40), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n407), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n616), .B2(new_n617), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n592), .A2(new_n595), .A3(new_n620), .A4(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT37), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n495), .A2(new_n626), .A3(new_n499), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n509), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n496), .A2(new_n498), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n626), .B1(new_n630), .B2(new_n430), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n497), .B1(new_n491), .B2(new_n494), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT38), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n504), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n628), .B1(KEYINPUT37), .B2(new_n508), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n597), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n625), .A2(new_n637), .A3(new_n585), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n602), .A2(new_n609), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n600), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n335), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n416), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G1gat), .ZN(G1324gat));
  INV_X1    g443(.A(new_n641), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n596), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT16), .B(G8gat), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT103), .ZN(new_n651));
  OAI221_X1 g450(.A(new_n651), .B1(new_n649), .B2(new_n648), .C1(new_n209), .C2(new_n646), .ZN(G1325gat));
  INV_X1    g451(.A(new_n591), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n645), .A2(G15gat), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G15gat), .B1(new_n645), .B2(new_n602), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n608), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  NOR3_X1   g458(.A1(new_n266), .A2(new_n314), .A3(new_n332), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n290), .B1(new_n600), .B2(new_n639), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n662), .A2(G29gat), .A3(new_n416), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT45), .Z(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  INV_X1    g464(.A(new_n290), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n640), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT104), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT104), .B1(new_n287), .B2(new_n289), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n665), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n639), .B2(new_n600), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n660), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT105), .B1(new_n673), .B2(new_n416), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G29gat), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n673), .A2(KEYINPUT105), .A3(new_n416), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n664), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT106), .Z(G1328gat));
  NOR3_X1   g477(.A1(new_n662), .A2(G36gat), .A3(new_n596), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT46), .ZN(new_n680));
  OAI21_X1  g479(.A(G36gat), .B1(new_n673), .B2(new_n596), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1329gat));
  OAI21_X1  g481(.A(G43gat), .B1(new_n673), .B2(new_n602), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n662), .A2(G43gat), .A3(new_n653), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n683), .A2(new_n688), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT47), .B1(new_n685), .B2(KEYINPUT107), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n690), .B(new_n692), .ZN(G1330gat));
  INV_X1    g492(.A(new_n673), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n608), .ZN(new_n695));
  INV_X1    g494(.A(new_n608), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n662), .A2(G50gat), .A3(new_n696), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n695), .A2(G50gat), .B1(KEYINPUT109), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(KEYINPUT48), .A2(G50gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n585), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n694), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n697), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(KEYINPUT48), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n698), .A2(KEYINPUT48), .B1(new_n701), .B2(new_n704), .ZN(G1331gat));
  INV_X1    g504(.A(new_n314), .ZN(new_n706));
  NOR4_X1   g505(.A1(new_n265), .A2(new_n666), .A3(new_n706), .A4(new_n333), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n640), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n416), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n596), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  AND2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n711), .B2(new_n712), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n708), .B2(new_n602), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n591), .A2(new_n294), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n708), .B2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g518(.A1(new_n708), .A2(new_n696), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n295), .ZN(G1335gat));
  NOR2_X1   g520(.A1(new_n265), .A2(new_n314), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n333), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n672), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n416), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT51), .B1(new_n661), .B2(new_n722), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n661), .A2(KEYINPUT51), .A3(new_n722), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n416), .A2(G85gat), .A3(new_n333), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  NOR3_X1   g532(.A1(new_n596), .A2(G92gat), .A3(new_n333), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n596), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n736), .B(new_n724), .C1(new_n667), .C2(new_n671), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G92gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n735), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n738), .A2(KEYINPUT110), .B1(new_n730), .B2(new_n734), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n737), .A2(new_n744), .A3(G92gat), .ZN(new_n745));
  AOI211_X1 g544(.A(KEYINPUT111), .B(new_n742), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n745), .A3(new_n735), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(KEYINPUT52), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n741), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(KEYINPUT113), .B(new_n741), .C1(new_n746), .C2(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1337gat));
  OAI21_X1  g554(.A(G99gat), .B1(new_n725), .B2(new_n602), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n653), .A2(G99gat), .A3(new_n333), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n731), .B2(new_n757), .ZN(G1338gat));
  NOR2_X1   g557(.A1(new_n725), .A2(new_n696), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT114), .B(G106gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n731), .A2(G106gat), .A3(new_n585), .A4(new_n333), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT53), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n764));
  NOR2_X1   g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766));
  INV_X1    g565(.A(new_n760), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n725), .B2(new_n585), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n765), .B2(new_n768), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n763), .B1(new_n769), .B2(new_n770), .ZN(G1339gat));
  NOR2_X1   g570(.A1(new_n668), .A2(new_n669), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n317), .B1(new_n325), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n330), .B(KEYINPUT54), .C1(new_n322), .C2(new_n324), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(KEYINPUT55), .A3(new_n775), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n331), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n262), .B2(new_n264), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n258), .A2(new_n259), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n243), .B1(new_n238), .B2(new_n242), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n251), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n261), .B2(new_n252), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(new_n333), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n772), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n785), .A2(new_n780), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n668), .B2(new_n669), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n314), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n265), .A2(new_n334), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n736), .A2(new_n416), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n793), .A2(new_n591), .A3(new_n696), .A4(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n795), .A2(new_n348), .A3(new_n266), .ZN(new_n796));
  NOR4_X1   g595(.A1(new_n792), .A2(new_n416), .A3(new_n736), .A4(new_n586), .ZN(new_n797));
  AOI21_X1  g596(.A(G113gat), .B1(new_n797), .B2(new_n265), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n796), .A2(new_n798), .ZN(G1340gat));
  NOR3_X1   g598(.A1(new_n795), .A2(new_n346), .A3(new_n333), .ZN(new_n800));
  AOI21_X1  g599(.A(G120gat), .B1(new_n797), .B2(new_n332), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(G1341gat));
  OAI21_X1  g601(.A(G127gat), .B1(new_n795), .B2(new_n706), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n797), .A2(new_n341), .A3(new_n314), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1342gat));
  NOR2_X1   g604(.A1(new_n792), .A2(new_n416), .ZN(new_n806));
  INV_X1    g605(.A(new_n586), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n666), .A2(new_n596), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n806), .A2(new_n339), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n810), .A2(KEYINPUT56), .ZN(new_n811));
  OAI21_X1  g610(.A(G134gat), .B1(new_n795), .B2(new_n290), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(KEYINPUT56), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(G1343gat));
  XNOR2_X1  g613(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n776), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n331), .A3(new_n779), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n262), .B2(new_n264), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n290), .B1(new_n818), .B2(new_n786), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT118), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n290), .C1(new_n818), .C2(new_n786), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n789), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n791), .B1(new_n823), .B2(new_n706), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT57), .B1(new_n824), .B2(new_n696), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n826), .B(new_n700), .C1(new_n790), .C2(new_n791), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n602), .A2(new_n794), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G141gat), .B1(new_n830), .B2(new_n266), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n602), .A2(new_n700), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n806), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n736), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n266), .A2(G141gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT58), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT119), .B1(new_n825), .B2(new_n829), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n825), .A2(KEYINPUT119), .A3(new_n829), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n265), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(KEYINPUT58), .A3(G141gat), .ZN(new_n843));
  NOR2_X1   g642(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n834), .B2(new_n836), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n838), .B1(new_n843), .B2(new_n845), .ZN(G1344gat));
  XOR2_X1   g645(.A(new_n791), .B(KEYINPUT121), .Z(new_n847));
  NAND2_X1  g646(.A1(new_n788), .A2(new_n666), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n819), .A2(KEYINPUT122), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n706), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT122), .B1(new_n819), .B2(new_n848), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n696), .A2(KEYINPUT57), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n700), .B1(new_n790), .B2(new_n791), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n852), .A2(new_n853), .B1(KEYINPUT57), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n855), .A2(new_n332), .A3(new_n828), .ZN(new_n856));
  INV_X1    g655(.A(G148gat), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT59), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n841), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(new_n839), .A3(new_n333), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n857), .A2(KEYINPUT59), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n834), .A2(new_n857), .A3(new_n332), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1345gat));
  NAND3_X1  g663(.A1(new_n834), .A2(new_n359), .A3(new_n314), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n859), .A2(new_n839), .A3(new_n706), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n359), .ZN(G1346gat));
  NOR3_X1   g666(.A1(new_n859), .A2(new_n839), .A3(new_n772), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n809), .A2(new_n360), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n868), .A2(new_n360), .B1(new_n833), .B2(new_n869), .ZN(G1347gat));
  NOR3_X1   g669(.A1(new_n653), .A2(new_n642), .A3(new_n596), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n793), .A2(new_n696), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT123), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n793), .A2(new_n874), .A3(new_n696), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n434), .A3(new_n266), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n792), .A2(new_n642), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n586), .A2(new_n596), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(G169gat), .B1(new_n881), .B2(new_n265), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n877), .A2(new_n882), .ZN(G1348gat));
  OAI21_X1  g682(.A(G176gat), .B1(new_n876), .B2(new_n333), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n435), .A3(new_n332), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1349gat));
  OAI21_X1  g685(.A(G183gat), .B1(new_n876), .B2(new_n706), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n881), .A2(new_n466), .A3(new_n468), .A4(new_n314), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT60), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n876), .B2(new_n290), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n880), .A2(G190gat), .A3(new_n772), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT124), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(G1351gat));
  AND2_X1   g699(.A1(new_n832), .A2(new_n736), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n878), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(G197gat), .B1(new_n903), .B2(new_n265), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n855), .A2(KEYINPUT125), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n855), .A2(KEYINPUT125), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n602), .A2(new_n416), .A3(new_n736), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n265), .A2(G197gat), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(G1352gat));
  XNOR2_X1  g710(.A(KEYINPUT126), .B(G204gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n332), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT62), .B1(new_n902), .B2(new_n913), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n902), .A2(KEYINPUT62), .A3(new_n913), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n908), .A2(new_n333), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n914), .B(new_n915), .C1(new_n916), .C2(new_n912), .ZN(G1353gat));
  OR3_X1    g716(.A1(new_n902), .A2(G211gat), .A3(new_n706), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n852), .A2(new_n853), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n907), .A2(new_n314), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n922), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT63), .B1(new_n922), .B2(G211gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT127), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n918), .B(new_n927), .C1(new_n923), .C2(new_n924), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1354gat));
  INV_X1    g728(.A(new_n772), .ZN(new_n930));
  AOI21_X1  g729(.A(G218gat), .B1(new_n903), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n666), .A2(G218gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n909), .B2(new_n932), .ZN(G1355gat));
endmodule


