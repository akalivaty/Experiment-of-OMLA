//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n188), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n191));
  XNOR2_X1  g005(.A(G143), .B(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G137), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT65), .A2(G134), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(KEYINPUT11), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT65), .A2(G134), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(G134), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(new_n202), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n193), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n192), .B2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n190), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n196), .A2(G137), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT65), .A2(G134), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n219), .A2(new_n220), .A3(new_n199), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n195), .A2(new_n197), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(G131), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n204), .B1(new_n198), .B2(new_n203), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n218), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n209), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT66), .B1(new_n227), .B2(G116), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(KEYINPUT2), .B(G113), .Z(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT28), .B1(new_n226), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n226), .A2(new_n236), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT68), .B(G237), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G953), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G210), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT70), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n244), .A3(G210), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT26), .B(G101), .Z(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n243), .A2(new_n249), .A3(new_n245), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(KEYINPUT71), .A3(new_n252), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n193), .A2(new_n205), .A3(new_n208), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n225), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G131), .B1(new_n221), .B2(new_n222), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n205), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n218), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n258), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT28), .A3(new_n236), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n239), .A2(new_n257), .A3(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(new_n266), .B(KEYINPUT74), .Z(new_n267));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n209), .A2(new_n225), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n264), .B2(new_n269), .ZN(new_n271));
  INV_X1    g085(.A(new_n236), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n264), .A2(new_n236), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n253), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n267), .A2(new_n268), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  AOI221_X4 g093(.A(new_n259), .B1(new_n211), .B2(new_n217), .C1(new_n261), .C2(new_n205), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT67), .B1(new_n262), .B2(new_n218), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n209), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n272), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n237), .A2(new_n285), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n276), .A2(new_n268), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n187), .B1(new_n278), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n270), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n282), .B2(KEYINPUT30), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n253), .B(new_n274), .C1(new_n293), .C2(new_n236), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT31), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n273), .A2(KEYINPUT31), .A3(new_n253), .A4(new_n274), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n257), .B1(new_n239), .B2(new_n265), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT32), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT72), .B1(new_n298), .B2(new_n300), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n302), .B(new_n299), .C1(new_n296), .C2(new_n297), .ZN(new_n309));
  OAI211_X1 g123(.A(KEYINPUT32), .B(new_n306), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT32), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n311), .A3(new_n310), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n291), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G210), .B1(G237), .B2(G902), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n319), .B(KEYINPUT89), .Z(new_n320));
  INV_X1    g134(.A(new_n234), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n235), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n227), .A3(G116), .ZN(new_n324));
  OAI211_X1 g138(.A(G113), .B(new_n324), .C1(new_n234), .C2(new_n323), .ZN(new_n325));
  INV_X1    g139(.A(G104), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT3), .B1(new_n326), .B2(G107), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n328));
  INV_X1    g142(.A(G107), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G104), .ZN(new_n330));
  INV_X1    g144(.A(G101), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(G107), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n327), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n326), .A2(G107), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n329), .A2(G104), .ZN(new_n335));
  OAI21_X1  g149(.A(G101), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n322), .A2(new_n325), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G122), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT86), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n330), .A3(new_n332), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G101), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n343), .A2(KEYINPUT4), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n272), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n343), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT83), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n348));
  OAI211_X1 g162(.A(KEYINPUT4), .B(new_n333), .C1(new_n343), .C2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n339), .B(new_n341), .C1(new_n345), .C2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n191), .B(new_n214), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n353));
  INV_X1    g167(.A(G125), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n211), .A2(new_n217), .A3(G125), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G224), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n353), .B1(new_n352), .B2(new_n354), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n322), .A2(new_n325), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n337), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n339), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n341), .B(KEYINPUT8), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT7), .ZN(new_n369));
  INV_X1    g183(.A(new_n360), .ZN(new_n370));
  OAI22_X1  g184(.A1(new_n357), .A2(new_n361), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n363), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n351), .B1(new_n372), .B2(KEYINPUT88), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(KEYINPUT88), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n339), .B1(new_n345), .B2(new_n350), .ZN(new_n375));
  INV_X1    g189(.A(new_n341), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n357), .A2(new_n361), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(new_n360), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n381), .A3(new_n376), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G902), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n320), .B1(new_n374), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n372), .A2(KEYINPUT88), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n372), .A2(KEYINPUT88), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n351), .ZN(new_n390));
  INV_X1    g204(.A(new_n320), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n390), .A2(new_n384), .A3(new_n391), .A4(new_n383), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n387), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT90), .B(new_n320), .C1(new_n374), .C2(new_n385), .ZN(new_n394));
  OAI21_X1  g208(.A(G214), .B1(G237), .B2(G902), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT85), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT20), .ZN(new_n399));
  NOR2_X1   g213(.A1(G475), .A2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n241), .A2(G214), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n212), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n241), .A2(G143), .A3(G214), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G131), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n204), .A3(new_n403), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n410));
  OR3_X1    g224(.A1(new_n354), .A2(KEYINPUT16), .A3(G140), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n410), .A2(G146), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(G146), .B1(new_n410), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n408), .B(new_n414), .C1(new_n406), .C2(new_n405), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n326), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n404), .A2(KEYINPUT18), .A3(G131), .ZN(new_n418));
  NAND2_X1  g232(.A1(KEYINPUT18), .A2(G131), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n402), .A2(new_n403), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n409), .A2(new_n189), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n409), .A2(new_n189), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n418), .B(new_n420), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n415), .A2(new_n417), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n405), .A2(new_n407), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n409), .B(KEYINPUT19), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n426), .A2(new_n189), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n412), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n425), .B(new_n429), .C1(new_n428), .C2(new_n427), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n417), .B1(new_n430), .B2(new_n423), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n399), .B(new_n400), .C1(new_n424), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n400), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n423), .ZN(new_n434));
  INV_X1    g248(.A(new_n417), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n415), .A2(new_n417), .A3(new_n423), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n417), .B1(new_n415), .B2(new_n423), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n384), .B1(new_n424), .B2(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT93), .B(G475), .Z(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(G234), .A2(G237), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(G952), .A3(new_n359), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(G902), .A3(G953), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(G898), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(G128), .B(G143), .Z(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n207), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n230), .A2(KEYINPUT14), .A3(G122), .ZN(new_n456));
  XNOR2_X1  g270(.A(G116), .B(G122), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(G107), .B(new_n456), .C1(new_n458), .C2(KEYINPUT14), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n455), .B(new_n459), .C1(G107), .C2(new_n458), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n457), .B(new_n329), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n212), .A3(G128), .ZN(new_n463));
  OAI211_X1 g277(.A(G134), .B(new_n463), .C1(new_n454), .C2(new_n462), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n461), .B(new_n464), .C1(new_n207), .C2(new_n454), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  INV_X1    g280(.A(G217), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n466), .A2(new_n467), .A3(G953), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n460), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n460), .B2(new_n465), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n384), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G478), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n471), .B(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n445), .A2(new_n453), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G469), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n193), .A2(new_n338), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n352), .A2(new_n337), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n262), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT84), .A2(KEYINPUT12), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n479), .A2(new_n482), .A3(new_n483), .A4(new_n262), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n218), .B(new_n344), .C1(new_n347), .C2(new_n349), .ZN(new_n488));
  INV_X1    g302(.A(new_n262), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n477), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n193), .A2(KEYINPUT10), .A3(new_n338), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n488), .A2(new_n489), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G110), .B(G140), .ZN(new_n494));
  INV_X1    g308(.A(G227), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(G953), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n494), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n487), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n262), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n498), .B1(new_n502), .B2(new_n493), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n476), .B(new_n384), .C1(new_n500), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n485), .A2(new_n493), .A3(new_n486), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n497), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n498), .A3(new_n493), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(G469), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n476), .A2(new_n384), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G221), .B1(new_n466), .B2(G902), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT82), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  OR3_X1    g329(.A1(new_n398), .A2(new_n475), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n467), .B1(G234), .B2(new_n384), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n412), .A2(new_n421), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n188), .A2(G119), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n227), .A2(G128), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT24), .B(G110), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT78), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n520), .B1(KEYINPUT77), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n521), .B(new_n528), .C1(new_n531), .C2(new_n520), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n526), .B1(G110), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n523), .B(KEYINPUT76), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT78), .B1(new_n534), .B2(new_n522), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n519), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(G110), .ZN(new_n537));
  OAI221_X1 g351(.A(new_n537), .B1(new_n522), .B2(new_n534), .C1(new_n412), .C2(new_n413), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(KEYINPUT80), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n359), .A2(G221), .A3(G234), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT79), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT22), .B(G137), .Z(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT80), .B1(new_n536), .B2(new_n538), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI211_X1 g360(.A(KEYINPUT80), .B(new_n543), .C1(new_n536), .C2(new_n538), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n384), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT25), .B(new_n384), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n518), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n546), .A2(new_n547), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n517), .A2(G902), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT81), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n318), .A2(new_n516), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(new_n331), .ZN(G3));
  AOI21_X1  g374(.A(G902), .B1(new_n303), .B2(new_n304), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G472), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n564));
  INV_X1    g378(.A(new_n515), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n563), .A2(new_n564), .A3(new_n314), .A4(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n314), .B1(new_n561), .B2(new_n187), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT94), .B1(new_n569), .B2(new_n566), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n460), .A2(new_n465), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT33), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n469), .B2(new_n470), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n469), .A2(new_n470), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT33), .A3(new_n574), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n576), .A2(new_n578), .A3(G478), .A4(new_n384), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT96), .B(G478), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n471), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n445), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n395), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n386), .B2(new_n392), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n584), .A2(new_n453), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n571), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G104), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  INV_X1    g405(.A(new_n586), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n452), .B(KEYINPUT99), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n438), .ZN(new_n596));
  INV_X1    g410(.A(new_n439), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT98), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n597), .B2(new_n596), .ZN(new_n599));
  INV_X1    g413(.A(new_n474), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n438), .A2(KEYINPUT98), .A3(new_n439), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n601), .A2(new_n444), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT100), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n571), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  INV_X1    g422(.A(new_n516), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n550), .A2(new_n551), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n517), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n536), .A2(new_n538), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT101), .Z(new_n613));
  NOR2_X1   g427(.A1(new_n543), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n555), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n609), .A2(new_n314), .A3(new_n563), .A4(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT37), .B(G110), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G12));
  INV_X1    g434(.A(new_n291), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n307), .A2(new_n312), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n314), .A2(KEYINPUT73), .A3(new_n315), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT102), .B(G900), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n448), .B1(new_n625), .B2(new_n450), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AND4_X1   g441(.A1(new_n586), .A2(new_n603), .A3(new_n617), .A4(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n624), .A2(new_n628), .A3(new_n565), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G128), .ZN(G30));
  AOI21_X1  g444(.A(new_n257), .B1(new_n274), .B2(new_n283), .ZN(new_n631));
  INV_X1    g445(.A(new_n275), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n632), .B2(new_n253), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n633), .B2(G902), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n622), .B2(new_n623), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n626), .B(KEYINPUT39), .Z(new_n636));
  NAND3_X1  g450(.A1(new_n565), .A2(KEYINPUT104), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n638));
  INV_X1    g452(.A(new_n636), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n638), .B1(new_n515), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(KEYINPUT40), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n637), .B2(new_n640), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n393), .A2(new_n394), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n393), .B2(new_n394), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n440), .A2(new_n444), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n600), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n617), .A2(new_n651), .A3(new_n585), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n635), .A2(new_n645), .A3(new_n649), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G143), .ZN(G45));
  AOI211_X1 g468(.A(new_n626), .B(new_n583), .C1(new_n440), .C2(new_n444), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n617), .A2(new_n586), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n624), .A2(new_n565), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  INV_X1    g474(.A(new_n500), .ZN(new_n661));
  INV_X1    g475(.A(new_n503), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n476), .B1(new_n663), .B2(new_n384), .ZN(new_n664));
  INV_X1    g478(.A(new_n504), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n664), .A2(new_n665), .A3(new_n513), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n624), .A2(new_n557), .A3(new_n587), .A4(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT41), .B(G113), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G15));
  INV_X1    g485(.A(new_n666), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n318), .A2(new_n558), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n605), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT106), .B(G116), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G18));
  NOR3_X1   g490(.A1(new_n657), .A2(new_n475), .A3(new_n672), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n624), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G119), .ZN(G21));
  AOI21_X1  g493(.A(new_n257), .B1(new_n288), .B2(KEYINPUT107), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(KEYINPUT107), .B2(new_n288), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n298), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n306), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n563), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n672), .A2(new_n651), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n557), .A3(new_n595), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G122), .ZN(G24));
  AND3_X1   g501(.A1(new_n655), .A2(new_n586), .A3(new_n666), .ZN(new_n688));
  AND4_X1   g502(.A1(new_n563), .A2(new_n688), .A3(new_n617), .A4(new_n683), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n354), .ZN(G27));
  AOI21_X1  g504(.A(new_n585), .B1(new_n393), .B2(new_n394), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n515), .B(KEYINPUT108), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n656), .A2(KEYINPUT42), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n624), .A2(new_n557), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n655), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n621), .A2(new_n316), .A3(new_n310), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n557), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT42), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n695), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n700), .B1(new_n695), .B2(new_n699), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G131), .ZN(G33));
  AND2_X1   g518(.A1(new_n603), .A2(new_n627), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n624), .A2(new_n557), .A3(new_n705), .A4(new_n693), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G134), .ZN(G36));
  NAND3_X1  g521(.A1(new_n440), .A2(new_n444), .A3(new_n582), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT43), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n440), .A2(new_n710), .A3(new_n444), .A4(new_n582), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n709), .A2(new_n617), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n569), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n712), .A2(KEYINPUT44), .A3(new_n569), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(KEYINPUT111), .A3(new_n691), .A4(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n506), .A2(new_n507), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n506), .A2(new_n507), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n476), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n722), .A3(KEYINPUT110), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT110), .B1(new_n719), .B2(new_n722), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n510), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n719), .A2(new_n722), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n509), .B1(new_n731), .B2(new_n723), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n728), .A2(new_n733), .A3(new_n504), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n514), .A3(new_n636), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n717), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n393), .A2(new_n394), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n395), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n713), .B2(new_n714), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT111), .B1(new_n740), .B2(new_n716), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n194), .ZN(G39));
  NOR3_X1   g557(.A1(new_n739), .A2(new_n557), .A3(new_n656), .ZN(new_n744));
  INV_X1    g558(.A(new_n733), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n504), .B1(new_n732), .B2(KEYINPUT46), .ZN(new_n746));
  OAI211_X1 g560(.A(KEYINPUT47), .B(new_n514), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT47), .B1(new_n734), .B2(new_n514), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n318), .B(new_n744), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G140), .ZN(G42));
  NAND3_X1  g565(.A1(new_n684), .A2(new_n617), .A3(new_n688), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n586), .A2(new_n650), .A3(new_n600), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n753), .A2(new_n515), .A3(new_n617), .A4(new_n626), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n635), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n629), .A2(new_n659), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n313), .A2(new_n317), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n515), .B1(new_n759), .B2(new_n621), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n689), .B1(new_n760), .B2(new_n628), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(KEYINPUT52), .A3(new_n659), .A4(new_n755), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n599), .A2(new_n602), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n600), .A2(new_n626), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n764), .A2(new_n691), .A3(new_n617), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n624), .A2(new_n565), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n684), .A2(new_n617), .A3(new_n655), .A4(new_n693), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n706), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n706), .A2(new_n767), .A3(new_n771), .A4(new_n768), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n398), .A2(new_n594), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n650), .A2(new_n474), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n568), .A2(new_n570), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n618), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n568), .A2(new_n570), .A3(new_n584), .A4(new_n774), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n779), .B2(new_n559), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n609), .A2(new_n624), .A3(new_n557), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n568), .A2(new_n570), .A3(new_n584), .A4(new_n774), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(KEYINPUT113), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n777), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n763), .A2(new_n773), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n686), .A2(new_n678), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n673), .B2(new_n605), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n703), .A2(new_n669), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n785), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n789), .B1(new_n785), .B2(new_n788), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(KEYINPUT54), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n695), .A2(new_n699), .A3(KEYINPUT53), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n669), .A2(new_n787), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n763), .A3(new_n784), .A4(new_n773), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n793), .B1(new_n792), .B2(KEYINPUT54), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n684), .A2(new_n557), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n709), .A2(new_n448), .A3(new_n711), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n649), .A2(new_n395), .A3(new_n672), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(KEYINPUT50), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n684), .A2(new_n617), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n739), .A2(new_n672), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n803), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n807), .A2(new_n808), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n635), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n557), .A3(new_n448), .A4(new_n810), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT116), .Z(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n445), .A3(new_n583), .ZN(new_n817));
  INV_X1    g631(.A(new_n804), .ZN(new_n818));
  INV_X1    g632(.A(new_n749), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n747), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n664), .A2(new_n665), .A3(new_n514), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n818), .B(new_n691), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n813), .A2(new_n817), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n811), .A2(new_n698), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT117), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n804), .A2(new_n592), .A3(new_n672), .ZN(new_n829));
  INV_X1    g643(.A(G952), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n829), .A2(new_n830), .A3(G953), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n828), .B(new_n833), .C1(new_n584), .C2(new_n816), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n823), .A2(new_n824), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n825), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n800), .A2(new_n801), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(G952), .A2(G953), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n557), .A2(new_n397), .A3(new_n514), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT112), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n664), .A2(new_n665), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT49), .Z(new_n842));
  OR4_X1    g656(.A1(new_n649), .A2(new_n840), .A3(new_n708), .A4(new_n842), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n837), .A2(new_n838), .B1(new_n635), .B2(new_n843), .ZN(G75));
  XOR2_X1   g658(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n845));
  AND2_X1   g659(.A1(new_n378), .A2(new_n382), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(new_n380), .Z(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n384), .B1(new_n791), .B2(new_n797), .ZN(new_n849));
  AOI211_X1 g663(.A(KEYINPUT56), .B(new_n848), .C1(new_n849), .C2(new_n320), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n791), .A2(new_n797), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(G902), .A3(new_n320), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n845), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n384), .B(new_n391), .C1(new_n791), .C2(new_n797), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n848), .B1(new_n856), .B2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n852), .A2(new_n853), .A3(new_n847), .ZN(new_n858));
  INV_X1    g672(.A(new_n845), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n359), .A2(G952), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n855), .A2(new_n860), .A3(new_n862), .ZN(G51));
  XNOR2_X1  g677(.A(new_n851), .B(new_n798), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n509), .B(KEYINPUT119), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT57), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n663), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n849), .A2(new_n731), .A3(new_n723), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(G54));
  AND3_X1   g683(.A1(new_n849), .A2(KEYINPUT58), .A3(G475), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n436), .A2(new_n437), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n862), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(G60));
  NAND2_X1  g687(.A1(new_n576), .A2(new_n578), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT120), .Z(new_n875));
  NAND2_X1  g689(.A1(G478), .A2(G902), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT59), .Z(new_n877));
  OR2_X1    g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n862), .B1(new_n864), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n877), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n800), .B2(new_n801), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n881), .B2(new_n875), .ZN(G63));
  NAND2_X1  g696(.A1(G217), .A2(G902), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT60), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n791), .B2(new_n797), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n615), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n886), .B(new_n862), .C1(new_n553), .C2(new_n885), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(G66));
  INV_X1    g703(.A(new_n451), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n359), .B1(new_n890), .B2(G224), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n784), .A2(new_n669), .A3(new_n787), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n359), .ZN(new_n893));
  INV_X1    g707(.A(G898), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n846), .B1(new_n894), .B2(G953), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n893), .B(new_n895), .ZN(G69));
  XNOR2_X1  g710(.A(new_n271), .B(new_n426), .ZN(new_n897));
  NAND2_X1  g711(.A1(G900), .A2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n750), .B1(new_n737), .B2(new_n741), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n698), .A2(new_n753), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n736), .A2(new_n901), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n659), .A2(new_n761), .A3(new_n902), .A4(new_n706), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n900), .A2(new_n703), .A3(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n897), .B(new_n898), .C1(new_n904), .C2(G953), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n761), .A2(new_n653), .A3(new_n659), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n761), .A2(KEYINPUT62), .A3(new_n653), .A4(new_n659), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n318), .A2(new_n558), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n584), .A2(new_n775), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n912), .A2(new_n739), .A3(new_n641), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n911), .A2(KEYINPUT121), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT121), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n899), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT122), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n910), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(G953), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n905), .B1(new_n922), .B2(new_n897), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n897), .A2(KEYINPUT123), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n359), .B(new_n924), .C1(G227), .C2(G900), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n923), .B(new_n925), .ZN(G72));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n927));
  INV_X1    g741(.A(new_n892), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n919), .A2(new_n928), .A3(new_n921), .ZN(new_n929));
  NAND2_X1  g743(.A1(G472), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT63), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT124), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n632), .A2(new_n276), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n931), .B1(new_n277), .B2(new_n294), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n792), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n632), .A2(new_n276), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n932), .B1(new_n904), .B2(new_n892), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(KEYINPUT125), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n941), .B(new_n932), .C1(new_n904), .C2(new_n892), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n861), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n935), .B(new_n937), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n927), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n943), .A2(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n943), .A2(new_n944), .ZN(new_n949));
  AOI22_X1  g763(.A1(new_n933), .A2(new_n934), .B1(new_n792), .B2(new_n936), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n947), .A2(new_n951), .ZN(G57));
endmodule


