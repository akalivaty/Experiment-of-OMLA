

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(KEYINPUT26), .ZN(n601) );
  INV_X1 U551 ( .A(KEYINPUT104), .ZN(n653) );
  XNOR2_X1 U552 ( .A(n653), .B(KEYINPUT31), .ZN(n654) );
  XNOR2_X1 U553 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U554 ( .A1(n678), .A2(n595), .ZN(n659) );
  INV_X1 U555 ( .A(KEYINPUT17), .ZN(n517) );
  XNOR2_X1 U556 ( .A(n517), .B(KEYINPUT66), .ZN(n518) );
  NOR2_X1 U557 ( .A1(G651), .A2(n574), .ZN(n783) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XNOR2_X2 U559 ( .A(n519), .B(n518), .ZN(n865) );
  NAND2_X1 U560 ( .A1(G138), .A2(n865), .ZN(n521) );
  INV_X1 U561 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U562 ( .A1(G2104), .A2(n522), .ZN(n868) );
  NAND2_X1 U563 ( .A1(G126), .A2(n868), .ZN(n520) );
  AND2_X1 U564 ( .A1(n521), .A2(n520), .ZN(n527) );
  AND2_X1 U565 ( .A1(n522), .A2(G2104), .ZN(n864) );
  NAND2_X1 U566 ( .A1(G102), .A2(n864), .ZN(n523) );
  XNOR2_X1 U567 ( .A(KEYINPUT91), .B(n523), .ZN(n525) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n869) );
  AND2_X1 U569 ( .A1(n869), .A2(G114), .ZN(n524) );
  NOR2_X1 U570 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U571 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U572 ( .A(n528), .B(KEYINPUT92), .Z(G164) );
  NAND2_X1 U573 ( .A1(n864), .A2(G101), .ZN(n529) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n529), .Z(n531) );
  NAND2_X1 U575 ( .A1(n868), .A2(G125), .ZN(n530) );
  NAND2_X1 U576 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U577 ( .A(n532), .B(KEYINPUT65), .ZN(n534) );
  NAND2_X1 U578 ( .A1(G113), .A2(n869), .ZN(n533) );
  NAND2_X1 U579 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U580 ( .A1(G137), .A2(n865), .ZN(n535) );
  XNOR2_X1 U581 ( .A(KEYINPUT67), .B(n535), .ZN(n536) );
  NOR2_X2 U582 ( .A1(n537), .A2(n536), .ZN(G160) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n786) );
  NAND2_X1 U584 ( .A1(G90), .A2(n786), .ZN(n540) );
  INV_X1 U585 ( .A(G651), .ZN(n544) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n574) );
  OR2_X1 U587 ( .A1(n544), .A2(n574), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT68), .B(n538), .Z(n788) );
  NAND2_X1 U589 ( .A1(G77), .A2(n788), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U591 ( .A(n541), .B(KEYINPUT9), .ZN(n543) );
  NAND2_X1 U592 ( .A1(G52), .A2(n783), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n549) );
  NOR2_X1 U594 ( .A1(G543), .A2(n544), .ZN(n546) );
  XNOR2_X1 U595 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n545) );
  XNOR2_X1 U596 ( .A(n546), .B(n545), .ZN(n782) );
  NAND2_X1 U597 ( .A1(n782), .A2(G64), .ZN(n547) );
  XOR2_X1 U598 ( .A(KEYINPUT70), .B(n547), .Z(n548) );
  NOR2_X1 U599 ( .A1(n549), .A2(n548), .ZN(G171) );
  NAND2_X1 U600 ( .A1(n786), .A2(G89), .ZN(n550) );
  XNOR2_X1 U601 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U602 ( .A1(G76), .A2(n788), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U604 ( .A(n553), .B(KEYINPUT5), .ZN(n558) );
  NAND2_X1 U605 ( .A1(G63), .A2(n782), .ZN(n555) );
  NAND2_X1 U606 ( .A1(G51), .A2(n783), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U609 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U610 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(G88), .A2(n786), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G75), .A2(n788), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U615 ( .A1(G62), .A2(n782), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G50), .A2(n783), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U618 ( .A1(n565), .A2(n564), .ZN(G166) );
  XNOR2_X1 U619 ( .A(KEYINPUT93), .B(G166), .ZN(G303) );
  NAND2_X1 U620 ( .A1(n788), .A2(G73), .ZN(n566) );
  XNOR2_X1 U621 ( .A(n566), .B(KEYINPUT2), .ZN(n573) );
  NAND2_X1 U622 ( .A1(G86), .A2(n786), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G48), .A2(n783), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U625 ( .A1(G61), .A2(n782), .ZN(n569) );
  XNOR2_X1 U626 ( .A(KEYINPUT87), .B(n569), .ZN(n570) );
  NOR2_X1 U627 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n573), .A2(n572), .ZN(G305) );
  NAND2_X1 U629 ( .A1(G74), .A2(G651), .ZN(n579) );
  NAND2_X1 U630 ( .A1(G49), .A2(n783), .ZN(n576) );
  NAND2_X1 U631 ( .A1(G87), .A2(n574), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U633 ( .A1(n782), .A2(n577), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U635 ( .A(n580), .B(KEYINPUT86), .ZN(G288) );
  AND2_X1 U636 ( .A1(G72), .A2(n788), .ZN(n584) );
  NAND2_X1 U637 ( .A1(G85), .A2(n786), .ZN(n582) );
  NAND2_X1 U638 ( .A1(G60), .A2(n782), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U640 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n783), .A2(G47), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n586), .A2(n585), .ZN(G290) );
  NAND2_X1 U643 ( .A1(G65), .A2(n782), .ZN(n588) );
  NAND2_X1 U644 ( .A1(G53), .A2(n783), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U646 ( .A(KEYINPUT72), .B(n589), .Z(n591) );
  NAND2_X1 U647 ( .A1(n786), .A2(G91), .ZN(n590) );
  NAND2_X1 U648 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U649 ( .A1(G78), .A2(n788), .ZN(n592) );
  XNOR2_X1 U650 ( .A(KEYINPUT71), .B(n592), .ZN(n593) );
  NOR2_X1 U651 ( .A1(n594), .A2(n593), .ZN(n1000) );
  NOR2_X1 U652 ( .A1(G1384), .A2(G164), .ZN(n678) );
  NAND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n677) );
  INV_X1 U654 ( .A(n677), .ZN(n595) );
  INV_X1 U655 ( .A(n659), .ZN(n642) );
  NAND2_X1 U656 ( .A1(n642), .A2(G2072), .ZN(n596) );
  XNOR2_X1 U657 ( .A(n596), .B(KEYINPUT27), .ZN(n598) );
  XNOR2_X1 U658 ( .A(G1956), .B(KEYINPUT101), .ZN(n912) );
  NOR2_X1 U659 ( .A1(n912), .A2(n642), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n598), .A2(n597), .ZN(n600) );
  NOR2_X1 U661 ( .A1(n1000), .A2(n600), .ZN(n599) );
  XOR2_X1 U662 ( .A(n599), .B(KEYINPUT28), .Z(n638) );
  NAND2_X1 U663 ( .A1(n1000), .A2(n600), .ZN(n636) );
  INV_X1 U664 ( .A(G1996), .ZN(n939) );
  NOR2_X1 U665 ( .A1(n659), .A2(n939), .ZN(n602) );
  XNOR2_X1 U666 ( .A(n602), .B(n601), .ZN(n604) );
  NAND2_X1 U667 ( .A1(n659), .A2(G1341), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n604), .A2(n603), .ZN(n616) );
  NAND2_X1 U669 ( .A1(n786), .A2(G81), .ZN(n605) );
  XNOR2_X1 U670 ( .A(n605), .B(KEYINPUT12), .ZN(n607) );
  NAND2_X1 U671 ( .A1(G68), .A2(n788), .ZN(n606) );
  NAND2_X1 U672 ( .A1(n607), .A2(n606), .ZN(n609) );
  XOR2_X1 U673 ( .A(KEYINPUT13), .B(KEYINPUT76), .Z(n608) );
  XNOR2_X1 U674 ( .A(n609), .B(n608), .ZN(n613) );
  NAND2_X1 U675 ( .A1(G56), .A2(n782), .ZN(n610) );
  XNOR2_X1 U676 ( .A(n610), .B(KEYINPUT14), .ZN(n611) );
  XNOR2_X1 U677 ( .A(n611), .B(KEYINPUT75), .ZN(n612) );
  NOR2_X1 U678 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U679 ( .A1(n783), .A2(G43), .ZN(n614) );
  NAND2_X1 U680 ( .A1(n615), .A2(n614), .ZN(n993) );
  NOR2_X1 U681 ( .A1(n616), .A2(n993), .ZN(n617) );
  XOR2_X1 U682 ( .A(n617), .B(KEYINPUT64), .Z(n632) );
  NAND2_X1 U683 ( .A1(n783), .A2(G54), .ZN(n625) );
  NAND2_X1 U684 ( .A1(G92), .A2(n786), .ZN(n619) );
  NAND2_X1 U685 ( .A1(G66), .A2(n782), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U687 ( .A(KEYINPUT78), .B(n620), .ZN(n623) );
  NAND2_X1 U688 ( .A1(G79), .A2(n788), .ZN(n621) );
  XNOR2_X1 U689 ( .A(KEYINPUT79), .B(n621), .ZN(n622) );
  NOR2_X1 U690 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U691 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U692 ( .A(KEYINPUT15), .B(n626), .Z(n773) );
  OR2_X1 U693 ( .A1(n632), .A2(n773), .ZN(n631) );
  AND2_X1 U694 ( .A1(n642), .A2(G2067), .ZN(n627) );
  XOR2_X1 U695 ( .A(n627), .B(KEYINPUT102), .Z(n629) );
  NAND2_X1 U696 ( .A1(n659), .A2(G1348), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U699 ( .A1(n632), .A2(n773), .ZN(n633) );
  NAND2_X1 U700 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U701 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U702 ( .A1(n638), .A2(n637), .ZN(n640) );
  XNOR2_X1 U703 ( .A(KEYINPUT29), .B(KEYINPUT103), .ZN(n639) );
  XNOR2_X1 U704 ( .A(n640), .B(n639), .ZN(n646) );
  INV_X1 U705 ( .A(G1961), .ZN(n924) );
  NAND2_X1 U706 ( .A1(n659), .A2(n924), .ZN(n644) );
  XNOR2_X1 U707 ( .A(G2078), .B(KEYINPUT25), .ZN(n641) );
  XNOR2_X1 U708 ( .A(n641), .B(KEYINPUT100), .ZN(n943) );
  NAND2_X1 U709 ( .A1(n642), .A2(n943), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U711 ( .A1(n647), .A2(G171), .ZN(n645) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n657) );
  NOR2_X1 U713 ( .A1(G171), .A2(n647), .ZN(n652) );
  NAND2_X1 U714 ( .A1(G8), .A2(n659), .ZN(n726) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n726), .ZN(n672) );
  NOR2_X1 U716 ( .A1(G2084), .A2(n659), .ZN(n668) );
  NOR2_X1 U717 ( .A1(n672), .A2(n668), .ZN(n648) );
  NAND2_X1 U718 ( .A1(G8), .A2(n648), .ZN(n649) );
  XNOR2_X1 U719 ( .A(KEYINPUT30), .B(n649), .ZN(n650) );
  NOR2_X1 U720 ( .A1(G168), .A2(n650), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n667) );
  NAND2_X1 U723 ( .A1(n667), .A2(G286), .ZN(n664) );
  NOR2_X1 U724 ( .A1(G1971), .A2(n726), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n658), .B(KEYINPUT106), .ZN(n661) );
  NOR2_X1 U726 ( .A1(n659), .A2(G2090), .ZN(n660) );
  NOR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U728 ( .A1(n662), .A2(G303), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U730 ( .A1(G8), .A2(n665), .ZN(n666) );
  XOR2_X1 U731 ( .A(KEYINPUT32), .B(n666), .Z(n674) );
  XOR2_X1 U732 ( .A(n667), .B(KEYINPUT105), .Z(n670) );
  NAND2_X1 U733 ( .A1(n668), .A2(G8), .ZN(n669) );
  NAND2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U737 ( .A(KEYINPUT107), .B(n675), .ZN(n721) );
  NOR2_X1 U738 ( .A1(G2090), .A2(G303), .ZN(n676) );
  NAND2_X1 U739 ( .A1(G8), .A2(n676), .ZN(n711) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n750) );
  XNOR2_X1 U741 ( .A(KEYINPUT97), .B(KEYINPUT36), .ZN(n691) );
  NAND2_X1 U742 ( .A1(n869), .A2(G116), .ZN(n679) );
  XNOR2_X1 U743 ( .A(n679), .B(KEYINPUT96), .ZN(n681) );
  NAND2_X1 U744 ( .A1(G128), .A2(n868), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U746 ( .A(n682), .B(KEYINPUT35), .ZN(n689) );
  XNOR2_X1 U747 ( .A(KEYINPUT34), .B(KEYINPUT95), .ZN(n687) );
  NAND2_X1 U748 ( .A1(n864), .A2(G104), .ZN(n683) );
  XNOR2_X1 U749 ( .A(n683), .B(KEYINPUT94), .ZN(n685) );
  NAND2_X1 U750 ( .A1(G140), .A2(n865), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U752 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U754 ( .A(n691), .B(n690), .ZN(n881) );
  XNOR2_X1 U755 ( .A(G2067), .B(KEYINPUT37), .ZN(n748) );
  NOR2_X1 U756 ( .A1(n881), .A2(n748), .ZN(n982) );
  NAND2_X1 U757 ( .A1(n750), .A2(n982), .ZN(n746) );
  NAND2_X1 U758 ( .A1(n869), .A2(G117), .ZN(n693) );
  NAND2_X1 U759 ( .A1(G141), .A2(n865), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n864), .A2(G105), .ZN(n694) );
  XOR2_X1 U762 ( .A(KEYINPUT38), .B(n694), .Z(n695) );
  NOR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n868), .A2(G129), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n875) );
  AND2_X1 U766 ( .A1(n875), .A2(G1996), .ZN(n974) );
  NAND2_X1 U767 ( .A1(G95), .A2(n864), .ZN(n700) );
  NAND2_X1 U768 ( .A1(G131), .A2(n865), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U770 ( .A1(G119), .A2(n868), .ZN(n702) );
  NAND2_X1 U771 ( .A1(G107), .A2(n869), .ZN(n701) );
  NAND2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n880) );
  INV_X1 U774 ( .A(G1991), .ZN(n740) );
  NOR2_X1 U775 ( .A1(n880), .A2(n740), .ZN(n968) );
  OR2_X1 U776 ( .A1(n974), .A2(n968), .ZN(n705) );
  NAND2_X1 U777 ( .A1(n750), .A2(n705), .ZN(n739) );
  NAND2_X1 U778 ( .A1(n746), .A2(n739), .ZN(n706) );
  XOR2_X1 U779 ( .A(KEYINPUT98), .B(n706), .Z(n729) );
  NOR2_X1 U780 ( .A1(G1981), .A2(G305), .ZN(n707) );
  XNOR2_X1 U781 ( .A(n707), .B(KEYINPUT24), .ZN(n708) );
  XNOR2_X1 U782 ( .A(n708), .B(KEYINPUT99), .ZN(n709) );
  NOR2_X1 U783 ( .A1(n709), .A2(n726), .ZN(n710) );
  NAND2_X1 U784 ( .A1(n729), .A2(n710), .ZN(n713) );
  AND2_X1 U785 ( .A1(n711), .A2(n713), .ZN(n712) );
  NAND2_X1 U786 ( .A1(n721), .A2(n712), .ZN(n717) );
  INV_X1 U787 ( .A(n713), .ZN(n715) );
  AND2_X1 U788 ( .A1(n726), .A2(n729), .ZN(n714) );
  OR2_X1 U789 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U790 ( .A1(n717), .A2(n716), .ZN(n735) );
  NOR2_X1 U791 ( .A1(G1976), .A2(G288), .ZN(n724) );
  NOR2_X1 U792 ( .A1(G1971), .A2(G303), .ZN(n718) );
  NOR2_X1 U793 ( .A1(n724), .A2(n718), .ZN(n1004) );
  INV_X1 U794 ( .A(KEYINPUT33), .ZN(n719) );
  AND2_X1 U795 ( .A1(n1004), .A2(n719), .ZN(n720) );
  NAND2_X1 U796 ( .A1(n721), .A2(n720), .ZN(n733) );
  INV_X1 U797 ( .A(n726), .ZN(n722) );
  NAND2_X1 U798 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  AND2_X1 U799 ( .A1(n722), .A2(n1003), .ZN(n723) );
  NOR2_X1 U800 ( .A1(KEYINPUT33), .A2(n723), .ZN(n728) );
  NAND2_X1 U801 ( .A1(n724), .A2(KEYINPUT33), .ZN(n725) );
  NOR2_X1 U802 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U803 ( .A1(n728), .A2(n727), .ZN(n731) );
  XOR2_X1 U804 ( .A(G1981), .B(G305), .Z(n995) );
  AND2_X1 U805 ( .A1(n995), .A2(n729), .ZN(n730) );
  AND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U807 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U809 ( .A(G1986), .B(G290), .ZN(n1011) );
  NAND2_X1 U810 ( .A1(n1011), .A2(n750), .ZN(n736) );
  NAND2_X1 U811 ( .A1(n737), .A2(n736), .ZN(n753) );
  NOR2_X1 U812 ( .A1(n875), .A2(G1996), .ZN(n738) );
  XNOR2_X1 U813 ( .A(n738), .B(KEYINPUT108), .ZN(n977) );
  INV_X1 U814 ( .A(n739), .ZN(n743) );
  AND2_X1 U815 ( .A1(n740), .A2(n880), .ZN(n967) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U817 ( .A1(n967), .A2(n741), .ZN(n742) );
  NOR2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n977), .A2(n744), .ZN(n745) );
  XNOR2_X1 U820 ( .A(n745), .B(KEYINPUT39), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n881), .A2(n748), .ZN(n983) );
  NAND2_X1 U823 ( .A1(n749), .A2(n983), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U826 ( .A(n754), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U827 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U828 ( .A1(n868), .A2(G123), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n755), .B(KEYINPUT18), .ZN(n757) );
  NAND2_X1 U830 ( .A1(G135), .A2(n865), .ZN(n756) );
  NAND2_X1 U831 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U832 ( .A(KEYINPUT82), .B(n758), .ZN(n762) );
  NAND2_X1 U833 ( .A1(G99), .A2(n864), .ZN(n760) );
  NAND2_X1 U834 ( .A1(G111), .A2(n869), .ZN(n759) );
  NAND2_X1 U835 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n970) );
  XNOR2_X1 U837 ( .A(n970), .B(G2096), .ZN(n763) );
  XNOR2_X1 U838 ( .A(n763), .B(KEYINPUT83), .ZN(n764) );
  OR2_X1 U839 ( .A1(G2100), .A2(n764), .ZN(G156) );
  INV_X1 U840 ( .A(G132), .ZN(G219) );
  INV_X1 U841 ( .A(G82), .ZN(G220) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U843 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U844 ( .A(G223), .ZN(n821) );
  NAND2_X1 U845 ( .A1(n821), .A2(G567), .ZN(n766) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n781) );
  OR2_X1 U848 ( .A1(n993), .A2(n781), .ZN(G153) );
  XNOR2_X1 U849 ( .A(G171), .B(KEYINPUT77), .ZN(G301) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n768) );
  INV_X1 U851 ( .A(G868), .ZN(n769) );
  NAND2_X1 U852 ( .A1(n773), .A2(n769), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(G284) );
  XNOR2_X1 U854 ( .A(n1000), .B(KEYINPUT73), .ZN(G299) );
  NOR2_X1 U855 ( .A1(G286), .A2(n769), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT80), .ZN(n772) );
  NOR2_X1 U857 ( .A1(G299), .A2(G868), .ZN(n771) );
  NOR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(G297) );
  NAND2_X1 U859 ( .A1(n781), .A2(G559), .ZN(n774) );
  INV_X1 U860 ( .A(n773), .ZN(n994) );
  NAND2_X1 U861 ( .A1(n774), .A2(n994), .ZN(n775) );
  XNOR2_X1 U862 ( .A(n775), .B(KEYINPUT81), .ZN(n776) );
  XOR2_X1 U863 ( .A(KEYINPUT16), .B(n776), .Z(G148) );
  NOR2_X1 U864 ( .A1(G868), .A2(n993), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G868), .A2(n994), .ZN(n777) );
  NOR2_X1 U866 ( .A1(G559), .A2(n777), .ZN(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U868 ( .A1(G559), .A2(n994), .ZN(n780) );
  XOR2_X1 U869 ( .A(n993), .B(n780), .Z(n801) );
  NAND2_X1 U870 ( .A1(n781), .A2(n801), .ZN(n794) );
  NAND2_X1 U871 ( .A1(G67), .A2(n782), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G55), .A2(n783), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n793) );
  NAND2_X1 U874 ( .A1(n786), .A2(G93), .ZN(n787) );
  XNOR2_X1 U875 ( .A(n787), .B(KEYINPUT84), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G80), .A2(n788), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U878 ( .A(KEYINPUT85), .B(n791), .Z(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n803) );
  XOR2_X1 U880 ( .A(n794), .B(n803), .Z(G145) );
  XOR2_X1 U881 ( .A(KEYINPUT88), .B(KEYINPUT19), .Z(n795) );
  XNOR2_X1 U882 ( .A(G305), .B(n795), .ZN(n796) );
  XNOR2_X1 U883 ( .A(G288), .B(n796), .ZN(n798) );
  XNOR2_X1 U884 ( .A(G290), .B(G166), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n798), .B(n797), .ZN(n799) );
  XOR2_X1 U886 ( .A(n803), .B(n799), .Z(n800) );
  XNOR2_X1 U887 ( .A(G299), .B(n800), .ZN(n890) );
  XNOR2_X1 U888 ( .A(n801), .B(n890), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n802), .A2(G868), .ZN(n805) );
  OR2_X1 U890 ( .A1(G868), .A2(n803), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n805), .A2(n804), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n806) );
  XNOR2_X1 U893 ( .A(n806), .B(KEYINPUT89), .ZN(n807) );
  XNOR2_X1 U894 ( .A(KEYINPUT20), .B(n807), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n808), .A2(G2090), .ZN(n809) );
  XNOR2_X1 U896 ( .A(KEYINPUT21), .B(n809), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n810), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U898 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U899 ( .A(KEYINPUT74), .B(G57), .Z(G237) );
  NOR2_X1 U900 ( .A1(G220), .A2(G219), .ZN(n811) );
  XOR2_X1 U901 ( .A(KEYINPUT22), .B(n811), .Z(n812) );
  NOR2_X1 U902 ( .A1(G218), .A2(n812), .ZN(n813) );
  NAND2_X1 U903 ( .A1(G96), .A2(n813), .ZN(n826) );
  AND2_X1 U904 ( .A1(G2106), .A2(n826), .ZN(n818) );
  NAND2_X1 U905 ( .A1(G108), .A2(G120), .ZN(n814) );
  NOR2_X1 U906 ( .A1(G237), .A2(n814), .ZN(n815) );
  NAND2_X1 U907 ( .A1(G69), .A2(n815), .ZN(n825) );
  NAND2_X1 U908 ( .A1(G567), .A2(n825), .ZN(n816) );
  XOR2_X1 U909 ( .A(KEYINPUT90), .B(n816), .Z(n817) );
  NOR2_X1 U910 ( .A1(n818), .A2(n817), .ZN(G319) );
  INV_X1 U911 ( .A(G319), .ZN(n820) );
  NAND2_X1 U912 ( .A1(G661), .A2(G483), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U917 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G108), .ZN(G238) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XOR2_X1 U927 ( .A(KEYINPUT42), .B(G2078), .Z(n828) );
  XNOR2_X1 U928 ( .A(G2090), .B(G2084), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U930 ( .A(n829), .B(G2100), .Z(n831) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U933 ( .A(G2096), .B(KEYINPUT43), .Z(n833) );
  XNOR2_X1 U934 ( .A(KEYINPUT109), .B(G2678), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U936 ( .A(n835), .B(n834), .Z(G227) );
  XOR2_X1 U937 ( .A(KEYINPUT110), .B(G1986), .Z(n837) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U940 ( .A(n838), .B(KEYINPUT41), .Z(n840) );
  XNOR2_X1 U941 ( .A(G1971), .B(G1976), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U943 ( .A(G1981), .B(G1956), .Z(n842) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1961), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U946 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2474), .B(KEYINPUT111), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U949 ( .A1(n868), .A2(G124), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U951 ( .A1(G136), .A2(n865), .ZN(n848) );
  NAND2_X1 U952 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U953 ( .A(KEYINPUT112), .B(n850), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G100), .A2(n864), .ZN(n852) );
  NAND2_X1 U955 ( .A1(G112), .A2(n869), .ZN(n851) );
  NAND2_X1 U956 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U958 ( .A(KEYINPUT113), .B(n855), .Z(G162) );
  NAND2_X1 U959 ( .A1(G130), .A2(n868), .ZN(n857) );
  NAND2_X1 U960 ( .A1(G118), .A2(n869), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G106), .A2(n864), .ZN(n859) );
  NAND2_X1 U963 ( .A1(G142), .A2(n865), .ZN(n858) );
  NAND2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U965 ( .A(KEYINPUT45), .B(n860), .Z(n861) );
  NOR2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n970), .B(n863), .ZN(n879) );
  NAND2_X1 U968 ( .A1(G103), .A2(n864), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G139), .A2(n865), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G127), .A2(n868), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G115), .A2(n869), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n962) );
  XOR2_X1 U976 ( .A(G162), .B(n962), .Z(n877) );
  XOR2_X1 U977 ( .A(G160), .B(n875), .Z(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(n886) );
  XNOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U983 ( .A(G164), .B(n884), .Z(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U985 ( .A1(G37), .A2(n887), .ZN(G395) );
  XNOR2_X1 U986 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n993), .B(G286), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U989 ( .A(n891), .B(n890), .Z(n893) );
  XNOR2_X1 U990 ( .A(G171), .B(n994), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U992 ( .A1(G37), .A2(n894), .ZN(G397) );
  XOR2_X1 U993 ( .A(G2451), .B(G2430), .Z(n896) );
  XNOR2_X1 U994 ( .A(G2438), .B(G2443), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n902) );
  XOR2_X1 U996 ( .A(G2435), .B(G2454), .Z(n898) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n900) );
  XOR2_X1 U999 ( .A(G2446), .B(G2427), .Z(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U1001 ( .A(n902), .B(n901), .Z(n903) );
  NAND2_X1 U1002 ( .A1(G14), .A2(n903), .ZN(n909) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n909), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1006 ( .A1(n906), .A2(n905), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(n909), .ZN(G401) );
  XOR2_X1 U1011 ( .A(KEYINPUT125), .B(G4), .Z(n911) );
  XNOR2_X1 U1012 ( .A(G1348), .B(KEYINPUT59), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(n911), .B(n910), .ZN(n916) );
  XOR2_X1 U1014 ( .A(n912), .B(G20), .Z(n914) );
  XNOR2_X1 U1015 ( .A(G6), .B(G1981), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(KEYINPUT124), .B(G1341), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(G19), .B(n917), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1021 ( .A(KEYINPUT60), .B(n920), .Z(n922) );
  XNOR2_X1 U1022 ( .A(G1966), .B(G21), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(KEYINPUT126), .B(n923), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n924), .B(G5), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(G1986), .B(G24), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(G1971), .B(G22), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(G1976), .B(G23), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(KEYINPUT127), .B(n929), .ZN(n930) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1033 ( .A(KEYINPUT58), .B(n932), .Z(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1035 ( .A(KEYINPUT61), .B(n935), .Z(n936) );
  NOR2_X1 U1036 ( .A1(G16), .A2(n936), .ZN(n961) );
  XOR2_X1 U1037 ( .A(KEYINPUT120), .B(G34), .Z(n938) );
  XNOR2_X1 U1038 ( .A(G2084), .B(KEYINPUT54), .ZN(n937) );
  XNOR2_X1 U1039 ( .A(n938), .B(n937), .ZN(n955) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n953) );
  XNOR2_X1 U1041 ( .A(G32), .B(n939), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n940), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n941) );
  NOR2_X1 U1045 ( .A1(n942), .A2(n941), .ZN(n947) );
  XOR2_X1 U1046 ( .A(n943), .B(G27), .Z(n945) );
  XNOR2_X1 U1047 ( .A(G1991), .B(G25), .ZN(n944) );
  NOR2_X1 U1048 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1051 ( .A(KEYINPUT53), .B(n950), .Z(n951) );
  XNOR2_X1 U1052 ( .A(n951), .B(KEYINPUT119), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(KEYINPUT121), .B(n956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(G29), .A2(n957), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(n958), .B(KEYINPUT55), .ZN(n959) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n959), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n991) );
  XOR2_X1 U1060 ( .A(G2072), .B(n962), .Z(n963) );
  XNOR2_X1 U1061 ( .A(KEYINPUT118), .B(n963), .ZN(n965) );
  XOR2_X1 U1062 ( .A(G2078), .B(G164), .Z(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(KEYINPUT50), .B(n966), .ZN(n987) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n972) );
  XOR2_X1 U1066 ( .A(G2084), .B(G160), .Z(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n980) );
  XOR2_X1 U1070 ( .A(G2090), .B(G162), .Z(n975) );
  XNOR2_X1 U1071 ( .A(KEYINPUT116), .B(n975), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1073 ( .A(KEYINPUT51), .B(n978), .Z(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT117), .B(n985), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(KEYINPUT52), .B(n988), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n989), .A2(G29), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n1019) );
  XOR2_X1 U1082 ( .A(G16), .B(KEYINPUT56), .Z(n1017) );
  XOR2_X1 U1083 ( .A(G1341), .B(KEYINPUT123), .Z(n992) );
  XNOR2_X1 U1084 ( .A(n993), .B(n992), .ZN(n1015) );
  XNOR2_X1 U1085 ( .A(G1348), .B(n994), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G168), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(KEYINPUT57), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1009) );
  XNOR2_X1 U1090 ( .A(G1956), .B(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(G1971), .A2(G303), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(KEYINPUT122), .B(n1007), .Z(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(G171), .B(G1961), .Z(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(n1020), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

