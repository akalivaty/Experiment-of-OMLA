//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G113), .ZN(new_n190));
  INV_X1    g004(.A(G113), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G113), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT71), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G116), .ZN(new_n199));
  INV_X1    g013(.A(G116), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n193), .A2(new_n194), .A3(new_n197), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(new_n196), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n199), .A3(new_n201), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n204), .A2(new_n188), .B1(new_n199), .B2(new_n201), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n194), .B1(new_n207), .B2(new_n197), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT75), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n202), .B1(new_n210), .B2(KEYINPUT71), .ZN(new_n211));
  INV_X1    g025(.A(new_n197), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT72), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n213), .A2(new_n214), .A3(new_n205), .A4(new_n203), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT65), .B1(new_n217), .B2(G146), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G146), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n221), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(G143), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n223), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT1), .B1(new_n217), .B2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n222), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT70), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n225), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT66), .A2(G131), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT66), .A2(G131), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(G137), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n238), .A2(new_n241), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT68), .B1(new_n243), .B2(G134), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n246), .A2(new_n242), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n243), .A2(KEYINPUT68), .A3(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  OR3_X1    g064(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n247), .B2(new_n250), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n235), .A2(new_n245), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n256), .B(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n226), .B2(new_n222), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n255), .A2(new_n257), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n264), .A2(new_n245), .A3(KEYINPUT73), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT73), .B1(new_n264), .B2(new_n245), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT74), .B(new_n262), .C1(new_n265), .C2(new_n266), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n216), .A2(new_n253), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n269), .A2(new_n253), .A3(new_n270), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(new_n216), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT28), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n253), .A2(new_n209), .A3(new_n215), .ZN(new_n276));
  INV_X1    g090(.A(new_n267), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G237), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G210), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n282), .B(KEYINPUT27), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G101), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n279), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n264), .A2(new_n245), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n259), .A2(new_n261), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(new_n254), .B2(new_n256), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT67), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n262), .A2(new_n296), .A3(new_n291), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n253), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n213), .A2(new_n205), .A3(new_n203), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n271), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT28), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n278), .A3(new_n285), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n269), .A2(KEYINPUT30), .A3(new_n253), .A4(new_n270), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT30), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n306), .A3(new_n299), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n271), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n286), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n303), .A2(new_n287), .A3(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT78), .B(G902), .Z(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n274), .A2(KEYINPUT77), .A3(new_n278), .A4(new_n288), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n290), .A2(new_n310), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G472), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n285), .B1(new_n302), .B2(new_n278), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n269), .A2(new_n270), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n317), .B(new_n285), .C1(new_n318), .C2(new_n276), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n317), .B1(new_n271), .B2(new_n285), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n307), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT31), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT31), .B(new_n307), .C1(new_n320), .C2(new_n321), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(G472), .A2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n326), .A2(KEYINPUT32), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT32), .ZN(new_n330));
  INV_X1    g144(.A(new_n316), .ZN(new_n331));
  INV_X1    g145(.A(new_n325), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n285), .B1(new_n318), .B2(new_n276), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n319), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT31), .B1(new_n335), .B2(new_n307), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n331), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n330), .B1(new_n337), .B2(new_n327), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n315), .B1(new_n329), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(G214), .B1(G237), .B2(G902), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G210), .B1(G237), .B2(G902), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n281), .A2(G224), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n344), .B(KEYINPUT93), .Z(new_n345));
  AND4_X1   g159(.A1(new_n218), .A2(new_n221), .A3(new_n222), .A4(new_n224), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n229), .B1(new_n227), .B2(new_n228), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n232), .A2(KEYINPUT70), .A3(new_n233), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G125), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n294), .A2(G125), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT94), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n351), .B2(new_n352), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n345), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  INV_X1    g172(.A(new_n345), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n354), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT5), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n364), .B(G113), .C1(KEYINPUT5), .C2(new_n199), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n205), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(new_n367), .B2(G107), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G104), .ZN(new_n371));
  INV_X1    g185(.A(G101), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(G107), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n368), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n370), .A2(G104), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n367), .A2(G107), .ZN(new_n376));
  OAI21_X1  g190(.A(G101), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n366), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n368), .A2(new_n371), .A3(new_n373), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G101), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT4), .A3(new_n374), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n383), .A3(G101), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n379), .B1(new_n385), .B2(new_n299), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G122), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n363), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n384), .B(new_n382), .C1(new_n206), .C2(new_n208), .ZN(new_n389));
  INV_X1    g203(.A(new_n379), .ZN(new_n390));
  AND4_X1   g204(.A1(new_n363), .A2(new_n389), .A3(new_n390), .A4(new_n387), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT6), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT91), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n386), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n387), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT6), .A4(new_n397), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n362), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT92), .B1(new_n393), .B2(new_n397), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n386), .A2(new_n363), .A3(new_n387), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n387), .B(KEYINPUT8), .Z(new_n405));
  NAND2_X1  g219(.A1(new_n366), .A2(new_n378), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(new_n390), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n359), .A2(KEYINPUT7), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n408), .A2(new_n351), .A3(new_n352), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n351), .B2(new_n352), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n343), .B1(new_n401), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n402), .B2(new_n403), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n400), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n361), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n342), .A3(new_n412), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n341), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G110), .B(G140), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT87), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n281), .A2(G227), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT10), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n254), .A2(new_n232), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n225), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n374), .A2(new_n377), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n385), .A2(new_n262), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n374), .A2(new_n377), .A3(KEYINPUT10), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n235), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT88), .B1(new_n349), .B2(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n265), .A2(new_n266), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n431), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n225), .B(new_n378), .C1(new_n230), .C2(new_n234), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n430), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n291), .A2(KEYINPUT12), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT73), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n291), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n264), .A2(new_n245), .A3(KEYINPUT73), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n430), .A2(new_n440), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n443), .B1(new_n447), .B2(KEYINPUT12), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n425), .B1(new_n439), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n432), .B1(new_n235), .B2(new_n434), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n349), .A2(KEYINPUT88), .A3(new_n433), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n430), .A2(new_n426), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n382), .A2(new_n384), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n294), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n450), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n438), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n431), .A2(new_n437), .A3(KEYINPUT89), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n439), .A2(new_n425), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n449), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G469), .B1(new_n462), .B2(G902), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT90), .B(G469), .C1(new_n462), .C2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n448), .ZN(new_n467));
  INV_X1    g281(.A(new_n439), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n431), .A2(new_n437), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n438), .B1(new_n469), .B2(new_n450), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n470), .B2(new_n459), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n467), .B1(new_n471), .B2(new_n425), .ZN(new_n472));
  INV_X1    g286(.A(G469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n312), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n466), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G221), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT9), .B(G234), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G902), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G122), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G116), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n200), .A2(G122), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(new_n370), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n217), .A2(G128), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT13), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n223), .A2(G143), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n487), .A2(new_n488), .ZN(new_n492));
  OAI21_X1  g306(.A(G134), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n487), .A2(new_n490), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n240), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n486), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n494), .B(new_n240), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n485), .A2(new_n370), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n484), .A2(KEYINPUT14), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n484), .A2(KEYINPUT14), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n483), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G107), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n478), .A2(G217), .A3(new_n281), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n496), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n496), .B2(new_n503), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT98), .B(new_n312), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G478), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT15), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n510), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n281), .A2(G952), .ZN(new_n514));
  INV_X1    g328(.A(G234), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(new_n280), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n281), .B(new_n312), .C1(G234), .C2(G237), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT21), .B(G898), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(G475), .A2(G902), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT97), .ZN(new_n523));
  XNOR2_X1  g337(.A(G113), .B(G122), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(G104), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n280), .A2(new_n281), .A3(G214), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n217), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n280), .A2(new_n281), .A3(G143), .A4(G214), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n238), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n238), .A3(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G140), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT16), .B1(new_n535), .B2(G125), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n350), .A2(G140), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT85), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT84), .A2(G125), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT85), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n540), .A3(G140), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT84), .B(G125), .C1(new_n535), .C2(KEYINPUT85), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n536), .B1(new_n543), .B2(KEYINPUT16), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n544), .A2(new_n220), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n535), .A2(G125), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n537), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT19), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n543), .B2(KEYINPUT19), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n549), .A2(KEYINPUT96), .A3(new_n220), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT96), .B1(new_n549), .B2(new_n220), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n534), .B(new_n545), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT18), .ZN(new_n554));
  INV_X1    g368(.A(G131), .ZN(new_n555));
  OAI22_X1  g369(.A1(new_n530), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n528), .A2(KEYINPUT95), .A3(new_n557), .A4(new_n529), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n537), .A2(new_n546), .A3(new_n220), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n543), .A2(G146), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n556), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n526), .B1(new_n552), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n544), .B(G146), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n532), .A2(new_n565), .A3(new_n533), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n530), .A2(KEYINPUT17), .A3(new_n531), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n525), .B(new_n561), .C1(new_n564), .C2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n523), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT20), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT20), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n572), .B(new_n523), .C1(new_n563), .C2(new_n569), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n564), .A2(new_n568), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n526), .B1(new_n575), .B2(new_n562), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n479), .B1(new_n576), .B2(new_n569), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G475), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n521), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AND4_X1   g394(.A1(new_n421), .A2(new_n475), .A3(new_n481), .A4(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT23), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n582), .A2(new_n198), .A3(G128), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT82), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n583), .A2(new_n584), .B1(new_n198), .B2(G128), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT83), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n587), .A2(new_n582), .B1(new_n223), .B2(G119), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n587), .B2(new_n582), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT24), .B(G110), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT80), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G119), .B(G128), .ZN(new_n594));
  OAI22_X1  g408(.A1(new_n590), .A2(G110), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n545), .A3(new_n559), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n590), .A2(G110), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT81), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n593), .A2(new_n598), .A3(new_n594), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n593), .B2(new_n594), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n596), .B1(new_n601), .B2(new_n564), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT22), .B(G137), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n476), .A2(new_n515), .A3(G953), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n603), .B(new_n604), .Z(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n596), .B(new_n605), .C1(new_n601), .C2(new_n564), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n312), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT25), .ZN(new_n610));
  OAI21_X1  g424(.A(G217), .B1(new_n311), .B2(new_n515), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT79), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT25), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n607), .A2(new_n614), .A3(new_n312), .A4(new_n608), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n610), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n607), .A2(new_n608), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n479), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT86), .Z(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n339), .A2(new_n581), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  OAI21_X1  g437(.A(KEYINPUT99), .B1(new_n326), .B2(new_n311), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n337), .A2(new_n625), .A3(new_n312), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n626), .A3(G472), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n337), .A2(new_n327), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n475), .A2(new_n481), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND4_X1   g444(.A1(new_n621), .A2(new_n627), .A3(new_n628), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n520), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n401), .A2(new_n343), .A3(new_n413), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n342), .B1(new_n419), .B2(new_n412), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n340), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n506), .A2(new_n507), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT33), .Z(new_n637));
  NOR2_X1   g451(.A1(new_n311), .A2(new_n509), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n509), .B1(new_n636), .B2(new_n311), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n574), .A2(new_n578), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n631), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  XNOR2_X1  g461(.A(new_n574), .B(KEYINPUT100), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n513), .A2(new_n578), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n635), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n631), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n627), .A2(new_n628), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n606), .A2(KEYINPUT36), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n602), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n602), .A2(new_n656), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n619), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n657), .A2(new_n619), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT101), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n661), .A2(new_n616), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT102), .B1(new_n655), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n661), .A2(new_n616), .A3(new_n663), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n627), .A2(new_n666), .A3(new_n628), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n581), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n517), .B1(new_n518), .B2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n650), .A2(new_n664), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n421), .A2(new_n475), .A3(new_n481), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n339), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n673), .B(KEYINPUT39), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n630), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT38), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n633), .B2(new_n634), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n414), .A2(new_n420), .A3(KEYINPUT38), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n513), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n574), .B2(new_n578), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n664), .A2(new_n340), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n335), .A2(new_n307), .B1(new_n286), .B2(new_n273), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n691), .B2(G902), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n329), .B2(new_n338), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n681), .A2(new_n689), .A3(new_n690), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  INV_X1    g509(.A(new_n673), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n641), .A2(new_n642), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n664), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n339), .A2(new_n676), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  AOI21_X1  g514(.A(new_n425), .B1(new_n460), .B2(new_n439), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n461), .A2(new_n448), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n312), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n473), .A2(KEYINPUT103), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n704), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n472), .A2(new_n312), .A3(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n705), .A2(new_n481), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n339), .A2(new_n621), .A3(new_n644), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  OAI21_X1  g525(.A(KEYINPUT32), .B1(new_n326), .B2(new_n328), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n337), .A2(new_n330), .A3(new_n327), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n712), .A2(new_n713), .B1(G472), .B2(new_n314), .ZN(new_n714));
  INV_X1    g528(.A(new_n621), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n705), .A2(new_n481), .A3(new_n707), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n651), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NAND4_X1  g533(.A1(new_n708), .A2(new_n421), .A3(new_n580), .A4(new_n667), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT104), .B1(new_n714), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n340), .B1(new_n633), .B2(new_n634), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n667), .A2(new_n574), .A3(new_n578), .A4(new_n521), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n723), .A3(new_n716), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n339), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NAND4_X1  g542(.A1(new_n708), .A2(new_n421), .A3(new_n632), .A4(new_n687), .ZN(new_n729));
  OAI21_X1  g543(.A(G472), .B1(new_n326), .B2(new_n311), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n279), .A2(new_n286), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n332), .B2(new_n336), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n327), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n621), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT105), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(G472), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n337), .B2(new_n312), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n324), .A2(new_n325), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n328), .B1(new_n738), .B2(new_n731), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n737), .A2(new_n715), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n687), .A2(new_n705), .A3(new_n481), .A4(new_n707), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n635), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n735), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  NOR3_X1   g560(.A1(new_n737), .A2(new_n664), .A3(new_n739), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n722), .A2(new_n716), .A3(new_n697), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NOR2_X1   g564(.A1(new_n714), .A2(new_n715), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n474), .A2(new_n463), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n481), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n414), .A2(new_n420), .A3(new_n340), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n697), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT42), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n714), .B2(new_n715), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n339), .A2(KEYINPUT106), .A3(new_n621), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n753), .A2(new_n754), .A3(new_n697), .A4(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n760), .A2(new_n761), .A3(KEYINPUT107), .A4(new_n763), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n758), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n555), .ZN(G33));
  NOR2_X1   g583(.A1(new_n650), .A2(new_n673), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT108), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n756), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n240), .ZN(G36));
  INV_X1    g587(.A(new_n754), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n641), .A2(new_n574), .A3(new_n578), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT43), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n641), .A2(new_n777), .A3(new_n574), .A4(new_n578), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n667), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n627), .B2(new_n628), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n774), .B1(new_n780), .B2(KEYINPUT44), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n780), .A2(KEYINPUT44), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n784), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT110), .B1(new_n786), .B2(new_n781), .ZN(new_n787));
  NAND2_X1  g601(.A1(G469), .A2(G902), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n462), .A2(KEYINPUT45), .ZN(new_n789));
  OAI21_X1  g603(.A(G469), .B1(new_n462), .B2(KEYINPUT45), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n474), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n791), .B2(new_n792), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n480), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n679), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT109), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n785), .A2(new_n787), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(KEYINPUT111), .B(G137), .Z(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G39));
  NOR4_X1   g615(.A1(new_n339), .A2(new_n621), .A3(new_n697), .A4(new_n754), .ZN(new_n802));
  XNOR2_X1  g616(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n796), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n796), .A2(new_n803), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(KEYINPUT113), .B(G140), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G42));
  INV_X1    g622(.A(new_n693), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n705), .A2(new_n707), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT49), .Z(new_n811));
  NOR4_X1   g625(.A1(new_n715), .A2(new_n775), .A3(new_n341), .A4(new_n480), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n811), .A3(new_n685), .A4(new_n812), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT114), .Z(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n716), .A2(new_n754), .A3(new_n715), .A4(new_n516), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n642), .A3(new_n641), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n776), .A2(new_n778), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(new_n517), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n708), .A3(new_n774), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n818), .B1(new_n747), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n740), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n685), .A2(new_n341), .A3(new_n708), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT50), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n825), .A2(KEYINPUT119), .A3(new_n827), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n825), .A2(KEYINPUT50), .A3(new_n827), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n830), .B2(new_n832), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n823), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n804), .A2(new_n805), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n810), .A2(new_n481), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n754), .B(new_n824), .C1(new_n840), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n815), .B1(new_n837), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n838), .B1(new_n481), .B2(new_n810), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n824), .A2(new_n754), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n815), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n823), .B(new_n848), .C1(new_n835), .C2(new_n836), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n760), .A2(new_n761), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n822), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT48), .Z(new_n852));
  NOR2_X1   g666(.A1(new_n722), .A2(new_n716), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  OAI221_X1 g668(.A(new_n514), .B1(new_n817), .B2(new_n643), .C1(new_n824), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n845), .A2(new_n849), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n651), .A2(new_n717), .B1(new_n721), .B2(new_n726), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n643), .B(KEYINPUT115), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n574), .A2(new_n578), .A3(new_n513), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT116), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n635), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n631), .A2(new_n862), .B1(new_n735), .B2(new_n744), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n709), .A2(new_n622), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n858), .A2(new_n863), .A3(new_n669), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n747), .A2(new_n757), .A3(new_n755), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n578), .A2(new_n667), .A3(new_n686), .A4(new_n696), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n630), .A2(new_n648), .A3(new_n774), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n868), .B2(new_n714), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n766), .A2(new_n767), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n751), .A2(new_n755), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n762), .B1(new_n872), .B2(new_n697), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n772), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n421), .A2(new_n687), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n752), .A2(new_n664), .A3(new_n481), .A4(new_n696), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n693), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n677), .A2(new_n699), .A3(new_n879), .A4(new_n749), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n712), .A2(new_n713), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n675), .B1(new_n883), .B2(new_n315), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n884), .A2(new_n674), .B1(new_n747), .B2(new_n748), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n699), .A4(new_n879), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n882), .A2(new_n886), .A3(KEYINPUT117), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n880), .A2(KEYINPUT117), .A3(new_n881), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n875), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n882), .A2(new_n886), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n870), .A2(new_n874), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT54), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n893), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n874), .A4(new_n870), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n857), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n814), .B1(new_n901), .B2(new_n902), .ZN(G75));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n896), .A2(new_n898), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n311), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(new_n342), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n418), .B(new_n361), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n909), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n904), .B(new_n911), .C1(new_n906), .C2(new_n342), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n281), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n910), .A2(new_n912), .A3(new_n914), .ZN(G51));
  XOR2_X1   g729(.A(new_n788), .B(KEYINPUT57), .Z(new_n916));
  INV_X1    g730(.A(new_n899), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n472), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n906), .A2(new_n789), .A3(new_n790), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(G54));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n923));
  NAND2_X1  g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n312), .B(new_n924), .C1(new_n896), .C2(new_n898), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n563), .A2(new_n569), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n914), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n924), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n311), .A2(new_n905), .A3(new_n926), .A4(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n923), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n926), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n906), .B2(new_n924), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n925), .A2(new_n926), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT121), .A4(new_n914), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(G60));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n637), .B1(new_n900), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n637), .B(new_n937), .C1(new_n917), .C2(new_n918), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n914), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n905), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n617), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n913), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n659), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n947), .B(KEYINPUT61), .C1(new_n948), .C2(new_n945), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n945), .A2(new_n948), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n943), .B1(new_n896), .B2(new_n898), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n914), .B1(new_n952), .B2(new_n617), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n950), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n949), .A2(new_n954), .ZN(G66));
  NAND2_X1  g769(.A1(G224), .A2(G953), .ZN(new_n956));
  OAI22_X1  g770(.A1(new_n865), .A2(G953), .B1(new_n519), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n399), .B(new_n400), .C1(G898), .C2(new_n281), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT122), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  AND2_X1   g774(.A1(new_n885), .A2(new_n699), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n694), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n964));
  AOI211_X1 g778(.A(new_n754), .B(new_n680), .C1(new_n861), .C2(new_n859), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n839), .A2(new_n802), .B1(new_n965), .B2(new_n751), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n963), .A2(new_n799), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n281), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n304), .A2(new_n306), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(new_n549), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n672), .A2(G953), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT123), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT124), .B1(new_n768), .B2(new_n772), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n874), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n798), .A2(new_n421), .A3(new_n687), .A4(new_n850), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n961), .A2(new_n806), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n978), .A2(new_n799), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n974), .B1(new_n981), .B2(new_n281), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n972), .B1(new_n982), .B2(new_n971), .ZN(new_n983));
  INV_X1    g797(.A(G227), .ZN(new_n984));
  OAI221_X1 g798(.A(G953), .B1(new_n984), .B2(new_n672), .C1(new_n971), .C2(KEYINPUT125), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n985), .B(new_n972), .C1(new_n982), .C2(new_n971), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(G72));
  NOR2_X1   g803(.A1(new_n308), .A2(new_n285), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n799), .A2(new_n979), .A3(new_n980), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n865), .B(new_n991), .C1(new_n977), .C2(new_n975), .ZN(new_n992));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n990), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n995), .B1(new_n322), .B2(new_n309), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT126), .Z(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n890), .B2(new_n894), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n994), .B1(new_n967), .B2(new_n865), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n286), .B1(new_n307), .B2(new_n271), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n913), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n996), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n996), .A2(new_n1002), .A3(KEYINPUT127), .A4(new_n999), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(G57));
endmodule


