//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G234), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT74), .A2(G140), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT74), .A2(G140), .ZN(new_n193));
  OAI21_X1  g007(.A(G125), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT75), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT76), .A2(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT76), .A2(G125), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(G140), .A3(new_n198), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT75), .B(G125), .C1(new_n192), .C2(new_n193), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(KEYINPUT16), .A3(new_n199), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n198), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT16), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(G146), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(KEYINPUT23), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT77), .B(G110), .Z(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT66), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G128), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT23), .A4(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT72), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT66), .B(G128), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT72), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT23), .A4(G119), .ZN(new_n222));
  AOI211_X1 g036(.A(new_n212), .B(new_n213), .C1(new_n219), .C2(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT24), .B(G110), .Z(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(G119), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(new_n210), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n205), .B(new_n208), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n210), .A3(new_n224), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n201), .A2(G146), .A3(new_n204), .ZN(new_n229));
  AOI21_X1  g043(.A(G146), .B1(new_n201), .B2(new_n204), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n212), .B1(new_n219), .B2(new_n222), .ZN(new_n232));
  OAI21_X1  g046(.A(G110), .B1(new_n232), .B2(KEYINPUT73), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT73), .ZN(new_n234));
  AOI211_X1 g048(.A(new_n234), .B(new_n212), .C1(new_n219), .C2(new_n222), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(KEYINPUT78), .B(new_n227), .C1(new_n231), .C2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G137), .ZN(new_n238));
  INV_X1    g052(.A(G953), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n239), .A2(G221), .A3(G234), .ZN(new_n240));
  XOR2_X1   g054(.A(new_n238), .B(new_n240), .Z(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n219), .A2(new_n222), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n234), .B1(new_n244), .B2(new_n212), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n232), .A2(KEYINPUT73), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(G110), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n201), .A2(new_n204), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n207), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n205), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n250), .A3(new_n228), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT78), .B1(new_n251), .B2(new_n227), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n243), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n227), .B1(new_n231), .B2(new_n236), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(new_n241), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n189), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n255), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n237), .A3(new_n242), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n256), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n189), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n191), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n190), .A2(G902), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT79), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT25), .B1(new_n263), .B2(new_n189), .ZN(new_n270));
  AOI211_X1 g084(.A(new_n259), .B(G902), .C1(new_n262), .C2(new_n256), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n190), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n267), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n209), .A2(G116), .ZN(new_n276));
  INV_X1    g090(.A(G116), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G119), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT2), .B(G113), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n281), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G143), .B(G146), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n207), .A2(G143), .ZN(new_n291));
  INV_X1    g105(.A(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G146), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n289), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n287), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G131), .ZN(new_n298));
  INV_X1    g112(.A(G137), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G134), .ZN(new_n300));
  AND2_X1   g114(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n300), .B(KEYINPUT65), .C1(new_n301), .C2(new_n302), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G137), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT11), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n300), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n298), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g127(.A(G131), .B(new_n311), .C1(new_n305), .C2(new_n306), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n297), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n298), .B1(new_n300), .B2(new_n309), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n311), .B1(new_n305), .B2(new_n306), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n298), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n286), .A2(new_n319), .A3(G128), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n319), .B1(G143), .B2(new_n207), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n294), .B(new_n321), .C1(new_n220), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT1), .B1(new_n292), .B2(G146), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n216), .A2(G128), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n214), .A2(KEYINPUT66), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n321), .B1(new_n328), .B2(new_n294), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n320), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n318), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n315), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(new_n315), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n285), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT26), .B(G101), .ZN(new_n336));
  INV_X1    g150(.A(G237), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n239), .A3(G210), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n336), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n285), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n315), .A2(new_n331), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n335), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT31), .ZN(new_n345));
  INV_X1    g159(.A(new_n341), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n342), .B1(new_n315), .B2(new_n331), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n348), .B1(new_n350), .B2(new_n343), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n346), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT31), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n335), .A2(new_n356), .A3(new_n341), .A4(new_n343), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n345), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G472), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n189), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT32), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(new_n362), .A3(new_n359), .A4(new_n189), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n315), .A2(new_n331), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT30), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n315), .A2(new_n331), .A3(new_n332), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n342), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n343), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n346), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n347), .B1(new_n368), .B2(new_n349), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n341), .A3(new_n353), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT70), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT71), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n350), .A2(new_n343), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT28), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n353), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n341), .A2(KEYINPUT29), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n376), .B(new_n189), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n352), .B1(new_n350), .B2(new_n343), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n382), .A2(new_n354), .A3(new_n380), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT71), .B1(new_n383), .B2(G902), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n369), .A2(new_n371), .A3(KEYINPUT70), .A4(new_n372), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n375), .A2(new_n381), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n361), .A2(new_n363), .B1(new_n386), .B2(G472), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n187), .B1(new_n275), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n361), .A2(new_n363), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(G472), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n391), .A2(KEYINPUT80), .A3(new_n269), .A4(new_n274), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n220), .A2(G143), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n292), .A2(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G134), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n308), .A3(new_n395), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G116), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n277), .A2(KEYINPUT14), .A3(G122), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n405), .A2(G107), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT97), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n404), .A2(KEYINPUT97), .A3(new_n406), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n399), .B(new_n402), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n400), .B(new_n401), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n398), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT13), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n395), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n394), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n395), .A2(new_n414), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n394), .A2(new_n413), .A3(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n412), .B1(new_n420), .B2(G134), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT9), .B(G234), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n422), .A2(new_n188), .A3(G953), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n410), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n420), .A2(G134), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n411), .A2(new_n398), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n428), .B2(new_n409), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n189), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT98), .ZN(new_n431));
  INV_X1    g245(.A(G478), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(KEYINPUT15), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(new_n409), .A3(new_n423), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n424), .B1(new_n410), .B2(new_n421), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT98), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n189), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n431), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G952), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(KEYINPUT99), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(KEYINPUT99), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n239), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(G234), .B2(G237), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n189), .B(new_n239), .C1(G234), .C2(G237), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(G898), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n448), .B(KEYINPUT100), .Z(new_n449));
  OR2_X1    g263(.A1(new_n430), .A2(new_n433), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n439), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT94), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n196), .A2(KEYINPUT94), .A3(new_n199), .A4(new_n200), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(G146), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n208), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n337), .A2(new_n239), .A3(G214), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(KEYINPUT93), .B2(new_n292), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT93), .B(G143), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(KEYINPUT18), .A2(G131), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G113), .B(G122), .ZN(new_n465));
  INV_X1    g279(.A(G104), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n461), .A2(G131), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT17), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n461), .A2(G131), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n461), .A2(KEYINPUT17), .A3(G131), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n471), .A2(new_n249), .A3(new_n205), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n464), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n467), .B1(new_n464), .B2(new_n473), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n189), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT95), .B(G475), .Z(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n229), .B1(new_n470), .B2(new_n468), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n454), .A2(KEYINPUT19), .A3(new_n455), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT19), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n206), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n207), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n480), .A2(new_n484), .B1(new_n457), .B2(new_n463), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n474), .B1(new_n485), .B2(new_n467), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n479), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n451), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G214), .B1(G237), .B2(G902), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G122), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n466), .A2(KEYINPUT3), .A3(G107), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n466), .A2(KEYINPUT81), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT81), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G104), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n501), .A3(G107), .ZN(new_n502));
  AOI21_X1  g316(.A(G107), .B1(new_n499), .B2(new_n501), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT3), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n498), .B(new_n502), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT4), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(G101), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n285), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT83), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT82), .B(G101), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n509), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n502), .A2(new_n511), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT81), .B(G104), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT3), .B1(new_n515), .B2(G107), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n514), .A2(KEYINPUT83), .A3(new_n516), .A4(new_n498), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n506), .B1(new_n505), .B2(G101), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n508), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G101), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n500), .A2(G104), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n466), .A2(KEYINPUT81), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n401), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n466), .A2(G107), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n276), .A2(new_n278), .A3(KEYINPUT5), .ZN(new_n527));
  OAI21_X1  g341(.A(G113), .B1(new_n276), .B2(KEYINPUT5), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n283), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n526), .B(new_n529), .C1(new_n513), .C2(new_n517), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n496), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n497), .B1(new_n524), .B2(KEYINPUT3), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT83), .B1(new_n532), .B2(new_n514), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n510), .A2(new_n509), .A3(new_n512), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n519), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n508), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n526), .B1(new_n513), .B2(new_n517), .ZN(new_n538));
  INV_X1    g352(.A(new_n529), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n495), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n531), .A2(new_n541), .A3(KEYINPUT6), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n543), .B(new_n496), .C1(new_n520), .C2(new_n530), .ZN(new_n544));
  INV_X1    g358(.A(new_n202), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n320), .B(new_n545), .C1(new_n324), .C2(new_n329), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n202), .B1(new_n290), .B2(new_n296), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT89), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n202), .C1(new_n290), .C2(new_n296), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n239), .A2(G224), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n551), .B(new_n552), .Z(new_n553));
  NAND3_X1  g367(.A1(new_n542), .A2(new_n544), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n542), .A2(KEYINPUT90), .A3(new_n553), .A4(new_n544), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G210), .B1(G237), .B2(G902), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n546), .B2(new_n547), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(new_n560), .ZN(new_n563));
  INV_X1    g377(.A(new_n526), .ZN(new_n564));
  INV_X1    g378(.A(new_n527), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n528), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n528), .A2(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n283), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n518), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n495), .B(KEYINPUT8), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n571), .B(new_n572), .C1(new_n538), .C2(new_n529), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n541), .A2(new_n563), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n574), .A2(new_n575), .A3(new_n189), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n574), .B2(new_n189), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n558), .A2(new_n559), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n559), .B1(new_n558), .B2(new_n578), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n493), .B(new_n494), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G469), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n294), .B1(new_n322), .B2(new_n214), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT85), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT85), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n294), .B(new_n585), .C1(new_n214), .C2(new_n322), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n586), .A3(new_n320), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n518), .A2(new_n564), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n538), .B2(new_n330), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n313), .A2(new_n314), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n593), .A2(KEYINPUT86), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(KEYINPUT86), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n294), .B1(new_n220), .B2(new_n322), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT67), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n323), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n597), .B1(new_n600), .B2(new_n320), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n588), .A2(new_n597), .B1(new_n538), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT84), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n507), .A2(new_n297), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n535), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n535), .B2(new_n604), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n602), .B(new_n590), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(G110), .B(G140), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n239), .A2(G227), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n589), .A2(KEYINPUT86), .A3(new_n593), .A4(new_n591), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n596), .A2(new_n607), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n591), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n611), .B1(new_n615), .B2(new_n607), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT87), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI211_X1 g432(.A(KEYINPUT87), .B(new_n611), .C1(new_n615), .C2(new_n607), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n582), .B(new_n189), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n582), .A2(new_n189), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n607), .A2(new_n611), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n596), .A2(new_n607), .A3(new_n612), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n615), .A2(new_n622), .B1(new_n623), .B2(new_n610), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n621), .B1(new_n624), .B2(G469), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G221), .ZN(new_n627));
  INV_X1    g441(.A(new_n422), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n189), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT88), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT88), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n626), .A2(new_n633), .A3(new_n630), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n581), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n393), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(new_n511), .Z(G3));
  AND2_X1   g451(.A1(new_n269), .A2(new_n274), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n358), .A2(new_n189), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(KEYINPUT101), .A3(new_n360), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n639), .A2(new_n642), .A3(G472), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n633), .B1(new_n626), .B2(new_n630), .ZN(new_n645));
  AOI211_X1 g459(.A(KEYINPUT88), .B(new_n629), .C1(new_n620), .C2(new_n625), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n638), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n431), .A2(new_n438), .ZN(new_n649));
  NAND2_X1  g463(.A1(KEYINPUT103), .A2(KEYINPUT33), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n436), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n652));
  OAI21_X1  g466(.A(new_n651), .B1(new_n436), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n432), .A2(G902), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  OAI22_X1  g469(.A1(new_n649), .A2(G478), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n492), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n449), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n494), .B1(new_n579), .B2(new_n580), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(KEYINPUT102), .B(new_n494), .C1(new_n579), .C2(new_n580), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n648), .A2(new_n659), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n466), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NAND2_X1  g482(.A1(new_n439), .A2(new_n450), .ZN(new_n669));
  INV_X1    g483(.A(new_n491), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n489), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n669), .A2(new_n671), .A3(new_n479), .A4(new_n449), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT105), .Z(new_n673));
  AND3_X1   g487(.A1(new_n648), .A2(new_n664), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT35), .B(G107), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NOR2_X1   g490(.A1(new_n242), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n254), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n266), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n272), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n272), .A2(KEYINPUT106), .A3(new_n679), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n682), .A2(new_n683), .B1(new_n641), .B2(new_n643), .ZN(new_n684));
  INV_X1    g498(.A(new_n581), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n684), .B(new_n685), .C1(new_n646), .C2(new_n645), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  NAND2_X1  g502(.A1(new_n632), .A2(new_n634), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n662), .A2(new_n663), .B1(new_n682), .B2(new_n683), .ZN(new_n690));
  INV_X1    g504(.A(new_n492), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n669), .ZN(new_n692));
  INV_X1    g506(.A(G900), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n444), .B1(new_n693), .B2(new_n445), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n391), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n689), .A2(new_n690), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XOR2_X1   g513(.A(new_n694), .B(KEYINPUT39), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n689), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n558), .A2(new_n578), .ZN(new_n704));
  INV_X1    g518(.A(new_n559), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n558), .A2(new_n559), .A3(new_n578), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT38), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n669), .A2(new_n492), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n494), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n682), .A2(new_n683), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n335), .A2(new_n343), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n346), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n189), .B1(new_n377), .B2(new_n341), .ZN(new_n717));
  OAI21_X1  g531(.A(G472), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n389), .A2(KEYINPUT107), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT107), .B1(new_n389), .B2(new_n718), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n712), .A2(new_n713), .A3(new_n721), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n702), .A2(new_n703), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n292), .ZN(G45));
  NOR2_X1   g538(.A1(new_n657), .A2(new_n694), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n689), .A2(new_n690), .A3(new_n391), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT108), .B(G146), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G48));
  NOR2_X1   g542(.A1(new_n275), .A2(new_n387), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n189), .B1(new_n618), .B2(new_n619), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n731), .A2(new_n630), .A3(new_n620), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n664), .A3(new_n659), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NAND4_X1  g549(.A1(new_n729), .A2(new_n673), .A3(new_n664), .A4(new_n732), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  AND4_X1   g551(.A1(new_n630), .A2(new_n731), .A3(new_n620), .A4(new_n493), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n664), .A2(new_n738), .A3(new_n391), .A4(new_n713), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT109), .B(G119), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G21));
  XOR2_X1   g555(.A(KEYINPUT110), .B(G472), .Z(new_n742));
  NAND2_X1  g556(.A1(new_n639), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n379), .A2(new_n346), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n345), .A3(new_n357), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n359), .A3(new_n189), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n265), .A3(new_n268), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n732), .A2(new_n748), .A3(new_n449), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT102), .B1(new_n708), .B2(new_n494), .ZN(new_n750));
  INV_X1    g564(.A(new_n663), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n711), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n664), .A2(new_n754), .A3(new_n711), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n749), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(G122), .Z(G24));
  INV_X1    g571(.A(new_n747), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n713), .A2(new_n725), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n731), .A2(new_n630), .A3(new_n620), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n662), .B2(new_n663), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  NOR2_X1   g577(.A1(new_n265), .A2(new_n268), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n391), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n706), .A2(new_n630), .A3(new_n494), .A4(new_n707), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n622), .A2(new_n615), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n623), .A2(new_n610), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT112), .A4(G469), .ZN(new_n770));
  INV_X1    g584(.A(new_n621), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n624), .A2(G469), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n767), .B1(new_n775), .B2(new_n620), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n766), .A2(KEYINPUT42), .A3(new_n725), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n773), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n620), .A3(new_n771), .A4(new_n770), .ZN(new_n779));
  INV_X1    g593(.A(new_n494), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n579), .A2(new_n580), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n630), .A3(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n782), .A2(new_n387), .A3(new_n275), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT113), .B1(new_n783), .B2(new_n725), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n729), .A2(new_n776), .A3(KEYINPUT113), .A4(new_n725), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n777), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT114), .B(G131), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G33));
  NAND2_X1  g604(.A1(new_n783), .A2(new_n695), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  OAI21_X1  g606(.A(G469), .B1(new_n624), .B2(KEYINPUT45), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(KEYINPUT45), .B2(new_n624), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n621), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n620), .B1(new_n795), .B2(KEYINPUT46), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n630), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n700), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n798), .A2(KEYINPUT115), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT115), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n781), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT43), .B1(new_n691), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n691), .A2(new_n656), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n641), .A2(new_n643), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n807), .A2(new_n808), .A3(new_n713), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n803), .B1(new_n809), .B2(KEYINPUT44), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(KEYINPUT44), .B2(new_n809), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n802), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  NAND3_X1  g627(.A1(new_n275), .A2(new_n387), .A3(new_n725), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT47), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n798), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n798), .A2(new_n815), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n781), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  NAND2_X1  g634(.A1(new_n731), .A2(new_n620), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT49), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT117), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(KEYINPUT49), .ZN(new_n824));
  INV_X1    g638(.A(new_n806), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n764), .A3(new_n630), .A4(new_n494), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n709), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n823), .A2(new_n721), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n807), .A2(new_n444), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n748), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n760), .A2(new_n494), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT122), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n830), .A2(new_n832), .A3(new_n709), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT50), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n803), .A2(new_n760), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n713), .A3(new_n758), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n721), .A2(new_n444), .A3(new_n638), .A4(new_n835), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n838), .A2(new_n492), .A3(new_n656), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n834), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n816), .B(new_n817), .C1(new_n630), .C2(new_n821), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(KEYINPUT123), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT123), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n830), .A2(new_n803), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n840), .B(KEYINPUT51), .C1(new_n842), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n841), .A2(new_n844), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n834), .A2(new_n847), .A3(new_n837), .A4(new_n839), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n836), .A2(new_n766), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT48), .Z(new_n852));
  NOR2_X1   g666(.A1(new_n838), .A2(new_n657), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n732), .B1(new_n750), .B2(new_n751), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n830), .A2(new_n854), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n852), .A2(new_n443), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n846), .A2(new_n850), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n391), .B(new_n695), .C1(new_n645), .C2(new_n646), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n713), .B1(new_n750), .B2(new_n751), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n713), .A2(new_n725), .A3(new_n758), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n859), .A2(new_n860), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n664), .A2(new_n391), .A3(new_n713), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n725), .B1(new_n645), .B2(new_n646), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n680), .A2(new_n629), .A3(new_n694), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n779), .ZN(new_n868));
  INV_X1    g682(.A(new_n720), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n389), .A2(KEYINPUT107), .A3(new_n718), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n754), .B1(new_n664), .B2(new_n711), .ZN(new_n872));
  AOI211_X1 g686(.A(KEYINPUT111), .B(new_n710), .C1(new_n662), .C2(new_n663), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n858), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n726), .A2(new_n698), .A3(new_n762), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n779), .B(new_n867), .C1(new_n719), .C2(new_n720), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n753), .B2(new_n755), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT52), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT120), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT52), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n696), .B1(new_n634), .B2(new_n632), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n882), .A2(new_n690), .B1(new_n759), .B2(new_n761), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n874), .A3(new_n858), .A4(new_n726), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n736), .A2(new_n733), .A3(new_n739), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n756), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n669), .A2(new_n492), .A3(new_n694), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n391), .A2(new_n781), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n689), .A2(new_n891), .A3(new_n713), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n759), .A2(new_n776), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n791), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n889), .A2(new_n788), .A3(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n660), .A2(new_n672), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n685), .B1(new_n645), .B2(new_n646), .ZN(new_n897));
  INV_X1    g711(.A(new_n684), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n647), .A2(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT118), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n808), .A2(new_n275), .ZN(new_n901));
  INV_X1    g715(.A(new_n896), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n689), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n686), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n708), .A2(new_n658), .A3(new_n494), .A4(new_n449), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n648), .A2(new_n907), .B1(new_n393), .B2(new_n635), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n900), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT119), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n900), .A2(new_n908), .A3(new_n911), .A4(new_n905), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n895), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n887), .A2(KEYINPUT53), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n862), .A2(KEYINPUT52), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n881), .A2(new_n884), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT54), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT53), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n881), .A2(new_n885), .A3(new_n884), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n885), .B1(new_n881), .B2(new_n884), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n889), .A2(new_n788), .A3(new_n894), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n904), .B1(new_n903), .B2(new_n686), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n689), .A2(new_n901), .A3(new_n907), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n636), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n911), .B1(new_n927), .B2(new_n905), .ZN(new_n928));
  INV_X1    g742(.A(new_n912), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n919), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT54), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n913), .A2(KEYINPUT53), .A3(new_n916), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n918), .A2(KEYINPUT121), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n936), .B(KEYINPUT54), .C1(new_n914), .C2(new_n917), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n857), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(G952), .A2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n828), .B1(new_n938), .B2(new_n939), .ZN(G75));
  NAND2_X1  g754(.A1(new_n931), .A2(new_n933), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(G210), .A3(G902), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT56), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n542), .A2(new_n544), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n553), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT55), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n942), .B2(new_n943), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n239), .A2(G952), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G51));
  AOI21_X1  g764(.A(KEYINPUT53), .B1(new_n887), .B2(new_n913), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n910), .A2(new_n912), .ZN(new_n952));
  AND4_X1   g766(.A1(KEYINPUT53), .A2(new_n952), .A3(new_n923), .A4(new_n916), .ZN(new_n953));
  OAI211_X1 g767(.A(G902), .B(new_n794), .C1(new_n951), .C2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT124), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n621), .B(KEYINPUT57), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n951), .A2(new_n953), .A3(KEYINPUT54), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n618), .A2(new_n619), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n949), .B1(new_n955), .B2(new_n961), .ZN(G54));
  AND2_X1   g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n941), .A2(G902), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  INV_X1    g779(.A(new_n486), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n949), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n964), .B2(new_n966), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n965), .B1(new_n964), .B2(new_n966), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(G60));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT59), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n653), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n957), .B2(new_n958), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n968), .ZN(new_n976));
  INV_X1    g790(.A(new_n973), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n935), .A2(new_n937), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n653), .B2(new_n978), .ZN(G63));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n941), .A2(new_n678), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n931), .B2(new_n933), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n983), .B(new_n968), .C1(new_n263), .C2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n984), .A2(new_n263), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n968), .A4(new_n983), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(G66));
  INV_X1    g804(.A(G224), .ZN(new_n991));
  OAI21_X1  g805(.A(G953), .B1(new_n446), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n952), .A2(new_n889), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(G953), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n944), .B1(G898), .B2(new_n239), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(G69));
  OR3_X1    g810(.A1(new_n239), .A2(KEYINPUT127), .A3(G900), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT127), .B1(new_n239), .B2(G900), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n819), .A2(new_n791), .A3(new_n866), .ZN(new_n999));
  INV_X1    g813(.A(new_n788), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n766), .B1(new_n872), .B2(new_n873), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n802), .B1(new_n811), .B2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n997), .B(new_n998), .C1(new_n1003), .C2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n481), .A2(new_n483), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT126), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n365), .A2(new_n366), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1006), .B(new_n1007), .Z(new_n1008));
  NAND2_X1  g822(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G227), .A2(G900), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(G953), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1008), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n723), .A2(new_n876), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT62), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n692), .A2(new_n657), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n1015), .B(new_n701), .C1(new_n388), .C2(new_n392), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n781), .B1(new_n818), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n812), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1012), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1009), .A2(new_n1011), .A3(new_n1020), .ZN(new_n1021));
  OAI211_X1 g835(.A(G953), .B(new_n1010), .C1(new_n1004), .C2(new_n1012), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(G72));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n1019), .B2(new_n993), .ZN(new_n1027));
  INV_X1    g841(.A(new_n716), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n968), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1026), .B1(new_n1003), .B2(new_n993), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n1030), .A2(new_n341), .A3(new_n714), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n914), .A2(new_n917), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n369), .A2(new_n344), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1032), .A2(new_n1026), .A3(new_n1033), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1029), .A2(new_n1031), .A3(new_n1034), .ZN(G57));
endmodule


