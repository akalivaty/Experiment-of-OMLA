//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  XOR2_X1   g020(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  AND3_X1   g047(.A1(new_n464), .A2(new_n470), .A3(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n471), .A2(G136), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g055(.A(G114), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT70), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G114), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n482), .A2(new_n484), .A3(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n461), .B1(new_n489), .B2(new_n490), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n466), .A2(new_n467), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n496), .A2(G138), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n500), .A3(new_n461), .A4(new_n493), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n492), .B1(new_n498), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n511), .A3(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n504), .B2(new_n506), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n509), .A2(new_n511), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n519));
  NOR4_X1   g094(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n519), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT72), .B(G651), .ZN(new_n522));
  OAI211_X1 g097(.A(G543), .B(new_n521), .C1(new_n522), .C2(new_n515), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT73), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n519), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n526), .A2(new_n527), .A3(G50), .A4(G543), .ZN(new_n528));
  AOI211_X1 g103(.A(new_n514), .B(new_n520), .C1(new_n525), .C2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n521), .B1(new_n522), .B2(new_n515), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n509), .A2(new_n511), .ZN(new_n534));
  INV_X1    g109(.A(new_n523), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT74), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  AOI22_X1  g116(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n507), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n531), .A2(new_n517), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n535), .A2(G52), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n517), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(new_n522), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT75), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n544), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n535), .A2(G43), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n517), .B(KEYINPUT77), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G651), .B1(G91), .B2(new_n544), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n523), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G299));
  XOR2_X1   g149(.A(new_n547), .B(KEYINPUT78), .Z(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G301));
  NAND2_X1  g151(.A1(new_n525), .A2(new_n528), .ZN(new_n577));
  INV_X1    g152(.A(new_n514), .ZN(new_n578));
  INV_X1    g153(.A(new_n520), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G303));
  OAI21_X1  g155(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n581));
  INV_X1    g156(.A(G49), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n526), .A2(new_n534), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n581), .B1(new_n582), .B2(new_n523), .C1(new_n583), .C2(new_n584), .ZN(G288));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT79), .B1(new_n523), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n526), .A2(new_n588), .A3(G48), .A4(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n544), .A2(G86), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n509), .A2(new_n511), .A3(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n507), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n544), .A2(G85), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  XOR2_X1   g173(.A(KEYINPUT80), .B(G47), .Z(new_n599));
  OAI221_X1 g174(.A(new_n597), .B1(new_n507), .B2(new_n598), .C1(new_n523), .C2(new_n599), .ZN(G290));
  AND3_X1   g175(.A1(new_n526), .A2(G92), .A3(new_n534), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT10), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n535), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n566), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n575), .B2(new_n609), .ZN(G284));
  OAI21_X1  g186(.A(new_n610), .B1(new_n575), .B2(new_n609), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  XOR2_X1   g190(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g191(.A(new_n608), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n499), .A2(new_n462), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n471), .A2(G135), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT82), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n475), .A2(G123), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G111), .C2(new_n461), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n629), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n627), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n651), .A2(G14), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT85), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(KEYINPUT18), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  AOI21_X1  g235(.A(KEYINPUT18), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT86), .ZN(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n665), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n674), .A2(new_n671), .A3(new_n669), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n669), .A2(new_n665), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n676), .A2(new_n673), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n672), .B(new_n675), .C1(new_n677), .C2(new_n671), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT87), .B(KEYINPUT88), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1991), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1996), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n683), .B(new_n685), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  OAI21_X1  g263(.A(KEYINPUT23), .B1(new_n614), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(G20), .ZN(new_n690));
  MUX2_X1   g265(.A(KEYINPUT23), .B(new_n689), .S(new_n690), .Z(new_n691));
  INV_X1    g266(.A(G1956), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G2090), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT89), .B(G29), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G35), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n695), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT29), .Z(new_n698));
  OAI21_X1  g273(.A(new_n693), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT97), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n471), .A2(G141), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT93), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT26), .Z(new_n705));
  AOI22_X1  g280(.A1(new_n475), .A2(G129), .B1(G105), .B2(new_n462), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G29), .B2(G32), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT94), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n688), .A2(G21), .ZN(new_n714));
  INV_X1    g289(.A(G1966), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n714), .B1(KEYINPUT95), .B2(new_n715), .C1(G168), .C2(new_n688), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT95), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  NAND2_X1  g293(.A1(G171), .A2(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G5), .B2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G1961), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(G160), .A2(G29), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT24), .B(G34), .Z(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n695), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n720), .B2(new_n721), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G33), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT25), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n471), .A2(G139), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n731), .B(new_n732), .C1(new_n461), .C2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n729), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT92), .B(G2072), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n722), .A2(new_n728), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G164), .A2(new_n695), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G27), .B2(new_n695), .ZN(new_n741));
  INV_X1    g316(.A(G2078), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n710), .B2(new_n711), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G28), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n746), .B2(G28), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n636), .B2(new_n695), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n749), .B1(new_n742), .B2(new_n741), .C1(new_n725), .C2(new_n726), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n713), .A2(new_n718), .A3(new_n739), .A4(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT31), .B(G11), .Z(new_n753));
  OR3_X1    g328(.A1(new_n752), .A2(KEYINPUT96), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT96), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n471), .A2(G140), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n475), .A2(G128), .ZN(new_n757));
  NOR2_X1   g332(.A1(G104), .A2(G2105), .ZN(new_n758));
  OAI21_X1  g333(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G29), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n762));
  INV_X1    g337(.A(G26), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n695), .B2(new_n763), .ZN(new_n764));
  OR3_X1    g339(.A1(new_n695), .A2(new_n762), .A3(new_n763), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n761), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2067), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n688), .A2(G4), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n617), .B2(new_n688), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1348), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n767), .B(new_n770), .C1(new_n694), .C2(new_n698), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n754), .A2(new_n755), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n701), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n688), .A2(G23), .ZN(new_n774));
  INV_X1    g349(.A(G288), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n688), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT33), .ZN(new_n777));
  INV_X1    g352(.A(G1976), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  MUX2_X1   g354(.A(G6), .B(G305), .S(G16), .Z(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n688), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n688), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n779), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT34), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n695), .A2(G25), .ZN(new_n790));
  OR2_X1    g365(.A1(G95), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT90), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n471), .A2(G131), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n475), .A2(G119), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(new_n695), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT35), .B(G1991), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n688), .A2(G24), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G290), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1986), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n805), .A2(new_n806), .A3(KEYINPUT91), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n789), .A2(new_n801), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n688), .A2(G19), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n557), .B2(new_n688), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1341), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n808), .A2(new_n809), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n773), .A2(new_n810), .A3(new_n813), .A4(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  AOI22_X1  g391(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(new_n507), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n544), .A2(G93), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n535), .A2(G55), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT100), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT37), .ZN(new_n824));
  INV_X1    g399(.A(new_n821), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n557), .A2(KEYINPUT99), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(KEYINPUT99), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n556), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n618), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT39), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n824), .B1(new_n836), .B2(G860), .ZN(G145));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n707), .B(new_n760), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n498), .A2(new_n501), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n475), .A2(G126), .B1(new_n485), .B2(new_n487), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n839), .A2(new_n842), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n734), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n845), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n847), .A2(new_n735), .A3(new_n843), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n625), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n471), .A2(G142), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n475), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n796), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n856), .A2(new_n857), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n850), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n862), .A2(new_n625), .A3(new_n858), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n838), .B1(new_n849), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n846), .A2(new_n848), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n864), .A3(KEYINPUT103), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT102), .B1(new_n849), .B2(new_n865), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n867), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n866), .B(new_n868), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n636), .B(G162), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G160), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n867), .B2(new_n864), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n869), .B2(new_n871), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n880));
  XNOR2_X1  g455(.A(G303), .B(G288), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G305), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G290), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n882), .A2(G290), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(G290), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(KEYINPUT105), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n880), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n883), .A2(KEYINPUT42), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT106), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n608), .B(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(KEYINPUT104), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(new_n614), .B2(new_n608), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n893), .B1(new_n897), .B2(KEYINPUT41), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n831), .B(new_n620), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n892), .B2(new_n899), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n890), .A2(KEYINPUT106), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n891), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n891), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g479(.A(G868), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n821), .A2(new_n609), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(G295));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n906), .ZN(G331));
  NAND2_X1  g483(.A1(G171), .A2(G286), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n575), .B2(G286), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n826), .A3(new_n830), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n831), .B(new_n909), .C1(G286), .C2(new_n575), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(new_n892), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n898), .B2(new_n913), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n885), .A2(new_n888), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT41), .B1(new_n894), .B2(new_n896), .ZN(new_n918));
  INV_X1    g493(.A(new_n892), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n918), .B(new_n913), .C1(KEYINPUT41), .C2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT107), .B1(new_n913), .B2(new_n892), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n911), .A2(new_n912), .A3(new_n922), .A4(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n888), .A3(new_n885), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n917), .A2(new_n925), .A3(KEYINPUT43), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n915), .A2(new_n916), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT43), .B1(new_n927), .B2(new_n917), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n917), .A2(new_n925), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n927), .B2(new_n917), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(G397));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G164), .B2(G1384), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n464), .A2(G40), .A3(new_n470), .A4(new_n472), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G2067), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n760), .B(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT108), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n940), .B1(new_n943), .B2(new_n708), .ZN(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT125), .B(KEYINPUT46), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n951));
  XNOR2_X1  g526(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n939), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT48), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n707), .B(new_n945), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n943), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n797), .A2(new_n800), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n796), .A2(new_n799), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n955), .B1(new_n960), .B2(new_n940), .ZN(new_n961));
  INV_X1    g536(.A(new_n959), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n957), .A2(new_n962), .B1(G2067), .B2(new_n760), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n939), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n952), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT63), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT109), .B1(new_n842), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n971), .B(G1384), .C1(new_n840), .C2(new_n841), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n968), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n840), .B2(new_n841), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n938), .B1(new_n975), .B2(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n694), .A3(new_n976), .ZN(new_n977));
  AND4_X1   g552(.A1(G40), .A2(new_n464), .A3(new_n470), .A4(new_n472), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n785), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n977), .A2(new_n985), .A3(new_n982), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(G8), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  NOR3_X1   g566(.A1(G166), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n984), .A2(KEYINPUT114), .A3(G8), .A4(new_n986), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n989), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n971), .B1(G164), .B2(G1384), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n974), .A2(KEYINPUT109), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n991), .B1(new_n999), .B2(new_n978), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n1002), .A2(new_n590), .A3(new_n591), .A4(new_n595), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n594), .B1(new_n587), .B2(new_n589), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n1004), .B2(new_n591), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1001), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G305), .A2(G1981), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1002), .A3(new_n591), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(KEYINPUT49), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1000), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT113), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1000), .A2(new_n1006), .A3(new_n1012), .A4(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n978), .B1(new_n970), .B2(new_n972), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n775), .A2(G1976), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(G8), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n775), .A2(G1976), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1015), .A2(KEYINPUT112), .A3(new_n1020), .A4(G8), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1014), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n997), .A2(new_n936), .A3(new_n998), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n938), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1966), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n973), .A2(new_n726), .A3(new_n976), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(G8), .A3(G168), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1026), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n967), .B1(new_n996), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT111), .B1(new_n992), .B2(new_n993), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n990), .B1(G166), .B2(new_n991), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n1038));
  NAND3_X1  g613(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n984), .A2(G8), .A3(new_n1041), .A4(new_n986), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n997), .A2(KEYINPUT50), .A3(new_n998), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n974), .A2(new_n968), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n694), .A4(new_n978), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n991), .B1(new_n1045), .B2(new_n982), .ZN(new_n1046));
  INV_X1    g621(.A(new_n994), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n967), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1042), .B1(new_n1033), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1014), .A2(new_n1025), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n775), .A2(new_n778), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1000), .B1(new_n1053), .B2(new_n1003), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1035), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT61), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1043), .A2(new_n978), .A3(new_n1044), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n980), .A2(new_n981), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT56), .B(G2072), .Z(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT115), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1059), .A2(new_n692), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n1064));
  XNOR2_X1  g639(.A(G299), .B(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1058), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n937), .A2(new_n945), .A3(new_n978), .A4(new_n979), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT118), .B(G1341), .Z(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT58), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1015), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1028), .A2(KEYINPUT117), .A3(new_n945), .A4(new_n937), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1074), .A2(KEYINPUT59), .A3(new_n557), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1348), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT50), .B1(new_n997), .B2(new_n998), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n978), .B1(new_n968), .B2(new_n974), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n938), .B1(new_n997), .B2(new_n998), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n941), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n602), .A2(KEYINPUT120), .A3(new_n603), .A4(new_n607), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n608), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n973), .A2(new_n976), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1089), .A2(new_n1077), .B1(new_n941), .B2(new_n1081), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1090), .A2(KEYINPUT60), .A3(new_n1083), .A4(new_n1086), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT60), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1088), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1059), .A2(new_n692), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT61), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1065), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1074), .A2(new_n557), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1098), .A2(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1063), .A2(new_n1065), .A3(new_n1058), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1076), .A2(new_n1095), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1065), .B(KEYINPUT116), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1063), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1090), .A2(new_n608), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT51), .B(G8), .C1(new_n1032), .C2(G286), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1031), .ZN(new_n1112));
  OAI21_X1  g687(.A(G8), .B1(new_n1112), .B2(new_n1029), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G286), .A2(G8), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1032), .A2(G8), .A3(G286), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1089), .A2(new_n721), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1028), .A2(new_n742), .A3(new_n937), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(G2078), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1027), .A2(new_n1028), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1119), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n575), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n981), .B2(new_n938), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n937), .A2(KEYINPUT123), .A3(new_n978), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n979), .A4(new_n1123), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1089), .B2(new_n721), .ZN(new_n1132));
  AOI211_X1 g707(.A(KEYINPUT122), .B(G1961), .C1(new_n973), .C2(new_n976), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1122), .B(new_n1130), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1126), .B1(new_n1134), .B2(new_n575), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1117), .A2(new_n1118), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1045), .A2(new_n982), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n994), .B1(new_n1138), .B2(new_n991), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1042), .A2(new_n1139), .A3(new_n1014), .A4(new_n1025), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1125), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1134), .A2(G171), .B1(new_n1141), .B2(G301), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1140), .B1(KEYINPUT54), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1110), .A2(new_n1137), .A3(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1056), .A2(new_n1144), .A3(KEYINPUT124), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT124), .B1(new_n1056), .B2(new_n1144), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1140), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n575), .B(new_n1125), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1145), .A2(new_n1146), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n960), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(G1986), .B2(G290), .ZN(new_n1156));
  INV_X1    g731(.A(new_n953), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n940), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n966), .B1(new_n1154), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g734(.A(G401), .B1(new_n875), .B2(new_n877), .ZN(new_n1161));
  INV_X1    g735(.A(G319), .ZN(new_n1162));
  OR2_X1    g736(.A1(G227), .A2(new_n1162), .ZN(new_n1163));
  AND2_X1   g737(.A1(new_n1163), .A2(KEYINPUT127), .ZN(new_n1164));
  NOR2_X1   g738(.A1(new_n1163), .A2(KEYINPUT127), .ZN(new_n1165));
  NOR3_X1   g739(.A1(G229), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI211_X1 g740(.A(new_n1161), .B(new_n1166), .C1(new_n932), .C2(new_n933), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


