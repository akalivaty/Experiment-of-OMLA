//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n640, new_n641, new_n643, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1274,
    new_n1275, new_n1276;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND3_X1   g033(.A1(new_n458), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n459));
  AOI21_X1  g034(.A(KEYINPUT66), .B1(new_n458), .B2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G101), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT65), .B1(new_n462), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n463), .A2(new_n466), .A3(new_n458), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT67), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n461), .B(new_n472), .C1(new_n468), .C2(new_n469), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n467), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND4_X1  g057(.A1(new_n463), .A2(new_n466), .A3(G2105), .A4(new_n467), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n458), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n468), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n476), .A2(new_n467), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n458), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n497), .A2(KEYINPUT68), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n495), .B1(new_n502), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI211_X1 g088(.A(G50), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n515), .A2(new_n516), .B1(new_n512), .B2(new_n513), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT69), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n505), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n508), .A2(new_n524), .A3(G88), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n526), .A3(new_n514), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n511), .B1(new_n520), .B2(new_n527), .ZN(G166));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n524), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n534), .B1(new_n508), .B2(new_n537), .ZN(G168));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n506), .A2(new_n507), .B1(new_n522), .B2(new_n523), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G90), .B1(new_n530), .B2(G52), .ZN(new_n541));
  OAI21_X1  g116(.A(G64), .B1(new_n516), .B2(new_n515), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n505), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n539), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g121(.A(G52), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n517), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g124(.A1(new_n549), .A2(new_n544), .A3(KEYINPUT70), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n546), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n506), .B2(new_n507), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g132(.A(G43), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n508), .A2(new_n524), .A3(G81), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(KEYINPUT71), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g144(.A(KEYINPUT71), .B(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n530), .A2(G53), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n540), .A2(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(G65), .B1(new_n516), .B2(new_n515), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT72), .B1(new_n576), .B2(G651), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n578));
  AOI211_X1 g153(.A(new_n578), .B(new_n505), .C1(new_n574), .C2(new_n575), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n572), .B(new_n573), .C1(new_n577), .C2(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n537), .A2(new_n508), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(new_n531), .A3(new_n533), .ZN(G286));
  INV_X1    g157(.A(new_n527), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n526), .B1(new_n525), .B2(new_n514), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n509), .A2(new_n510), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n583), .A2(new_n584), .B1(new_n505), .B2(new_n585), .ZN(G303));
  NAND2_X1  g161(.A1(new_n540), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n530), .A2(G49), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT73), .ZN(G288));
  AOI22_X1  g166(.A1(new_n540), .A2(G86), .B1(new_n530), .B2(G48), .ZN(new_n592));
  OAI21_X1  g167(.A(G61), .B1(new_n516), .B2(new_n515), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(KEYINPUT74), .B1(G73), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n595), .B(G61), .C1(new_n516), .C2(new_n515), .ZN(new_n596));
  AOI211_X1 g171(.A(KEYINPUT75), .B(new_n505), .C1(new_n594), .C2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n593), .A2(KEYINPUT74), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n599), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n598), .B1(new_n601), .B2(G651), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n592), .B1(new_n597), .B2(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(new_n530), .A2(G47), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n508), .A2(new_n524), .A3(G85), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT77), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n508), .A2(G60), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n612));
  NAND2_X1  g187(.A1(G72), .A2(G543), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G60), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n506), .B2(new_n507), .ZN(new_n616));
  INV_X1    g191(.A(new_n613), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT76), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n614), .A2(G651), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n610), .A2(new_n619), .ZN(G290));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(G301), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G92), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n517), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n540), .A2(G92), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n530), .A2(G54), .ZN(new_n628));
  INV_X1    g203(.A(G66), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n506), .B2(new_n507), .ZN(new_n630));
  AND2_X1   g205(.A1(G79), .A2(G543), .ZN(new_n631));
  OAI21_X1  g206(.A(G651), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT79), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n622), .B1(new_n621), .B2(new_n634), .ZN(G284));
  AOI21_X1  g210(.A(new_n622), .B1(new_n621), .B2(new_n634), .ZN(G321));
  NAND2_X1  g211(.A1(G299), .A2(new_n621), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n621), .B2(G168), .ZN(G297));
  OAI21_X1  g213(.A(new_n637), .B1(new_n621), .B2(G168), .ZN(G280));
  INV_X1    g214(.A(new_n634), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n640), .A2(G559), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(G860), .B2(new_n634), .ZN(G148));
  NAND2_X1  g217(.A1(new_n560), .A2(new_n621), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n641), .B2(new_n621), .ZN(G323));
  XOR2_X1   g219(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n645));
  XNOR2_X1  g220(.A(G323), .B(new_n645), .ZN(G282));
  OR2_X1    g221(.A1(new_n459), .A2(new_n460), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(new_n493), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G123), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n458), .A2(G111), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n655));
  OAI22_X1  g230(.A1(new_n483), .A2(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(G135), .B2(new_n488), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n652), .A2(new_n658), .ZN(G156));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n665), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G14), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT82), .ZN(G401));
  XNOR2_X1  g251(.A(G2084), .B(G2090), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2072), .B(G2078), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT83), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n680), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n677), .B(new_n681), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n677), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT18), .Z(new_n688));
  NOR2_X1   g263(.A1(new_n680), .A2(new_n677), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n685), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2096), .B(G2100), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G227));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT85), .ZN(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT86), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT19), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT20), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(new_n702), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n697), .A2(new_n699), .ZN(new_n706));
  MUX2_X1   g281(.A(new_n702), .B(new_n705), .S(new_n706), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n704), .A2(KEYINPUT87), .A3(new_n707), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n712), .B1(new_n710), .B2(new_n711), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n695), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(new_n695), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n717), .A2(new_n718), .A3(new_n713), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(G1981), .B(G1986), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n716), .A2(new_n719), .A3(new_n721), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(G229));
  NOR2_X1   g300(.A1(G5), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G171), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G2078), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n732), .A2(G2078), .ZN(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n736), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(G1966), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(G28), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n730), .B1(new_n740), .B2(G28), .ZN(new_n742));
  AND2_X1   g317(.A1(KEYINPUT31), .A2(G11), .ZN(new_n743));
  NOR2_X1   g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n657), .B2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n738), .A2(G1966), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n739), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n730), .A2(G33), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT25), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(new_n458), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n751), .B(new_n753), .C1(G139), .C2(new_n488), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(new_n730), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2072), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n734), .A2(new_n735), .A3(new_n748), .A4(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT96), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n647), .A2(new_n758), .A3(G105), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n647), .B2(G105), .ZN(new_n760));
  INV_X1    g335(.A(G129), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n483), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT97), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT26), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(KEYINPUT26), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n766), .A2(new_n767), .B1(G141), .B2(new_n488), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT98), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n763), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n730), .A2(G32), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT27), .B(G1996), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n730), .B1(KEYINPUT24), .B2(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(KEYINPUT24), .B2(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n481), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2084), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n757), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(KEYINPUT99), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT99), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n757), .A2(new_n786), .A3(new_n779), .A4(new_n783), .ZN(new_n787));
  NOR2_X1   g362(.A1(G4), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n634), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT92), .B(G1348), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT93), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n730), .A2(G26), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT28), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n488), .A2(G140), .ZN(new_n795));
  INV_X1    g370(.A(G128), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n458), .A2(G116), .ZN(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n798));
  OAI22_X1  g373(.A1(new_n483), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n794), .B1(new_n800), .B2(new_n730), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT95), .B(G2067), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G16), .A2(G19), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n561), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT94), .B(G1341), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n792), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n730), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n730), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT29), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(G2090), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(G2090), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n736), .A2(G20), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT23), .Z(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G299), .B2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G1956), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n808), .A2(new_n812), .A3(new_n813), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n785), .A2(new_n787), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(G16), .A2(G22), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G166), .B2(G16), .ZN(new_n822));
  INV_X1    g397(.A(G1971), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT32), .B(G1981), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n736), .A2(G6), .ZN(new_n826));
  INV_X1    g401(.A(new_n592), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n601), .A2(G651), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT75), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n505), .B1(new_n594), .B2(new_n596), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n598), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n826), .B1(new_n832), .B2(new_n736), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n736), .A2(G23), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n590), .B2(new_n736), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT33), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(G1976), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(G1976), .ZN(new_n838));
  OAI221_X1 g413(.A(new_n824), .B1(new_n825), .B2(new_n833), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n833), .A2(new_n825), .ZN(new_n840));
  OR3_X1    g415(.A1(new_n839), .A2(KEYINPUT34), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n736), .A2(G24), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G290), .B2(G16), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT90), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G1986), .ZN(new_n845));
  OR2_X1    g420(.A1(G95), .A2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n847));
  INV_X1    g422(.A(G131), .ZN(new_n848));
  INV_X1    g423(.A(G119), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n847), .B1(new_n468), .B2(new_n848), .C1(new_n849), .C2(new_n483), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT88), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n851), .A2(G29), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n730), .A2(G25), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G1991), .Z(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n845), .B1(new_n857), .B2(KEYINPUT89), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n857), .A2(KEYINPUT89), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT34), .B1(new_n839), .B2(new_n840), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n841), .A2(new_n858), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT91), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT36), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n864), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n820), .B1(new_n865), .B2(new_n866), .ZN(G311));
  INV_X1    g442(.A(G311), .ZN(G150));
  OAI211_X1 g443(.A(G55), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n869));
  INV_X1    g444(.A(G93), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n517), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  INV_X1    g447(.A(G67), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n506), .B2(new_n507), .ZN(new_n874));
  NAND2_X1  g449(.A1(G80), .A2(G543), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(G651), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n871), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G81), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n558), .B1(new_n517), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(G56), .B1(new_n516), .B2(new_n515), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n505), .B1(new_n881), .B2(new_n555), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT101), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n557), .A2(new_n884), .A3(new_n558), .A4(new_n559), .ZN(new_n885));
  OAI21_X1  g460(.A(G67), .B1(new_n516), .B2(new_n515), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n505), .B1(new_n886), .B2(new_n875), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT100), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n878), .A2(new_n883), .A3(new_n885), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n508), .A2(new_n524), .A3(G93), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n869), .B(new_n890), .C1(new_n887), .C2(KEYINPUT100), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n877), .A2(new_n872), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n560), .B(KEYINPUT101), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT38), .Z(new_n895));
  NAND2_X1  g470(.A1(new_n634), .A2(G559), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n898));
  INV_X1    g473(.A(G860), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n891), .A2(new_n892), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n902), .A2(new_n899), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(G145));
  AND2_X1   g480(.A1(new_n773), .A2(new_n754), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n754), .A2(new_n769), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G130), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n483), .A2(new_n909), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n458), .A2(KEYINPUT102), .A3(G118), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT102), .B1(new_n458), .B2(G118), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n910), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G142), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n649), .B(new_n916), .C1(new_n917), .C2(new_n468), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n648), .B(KEYINPUT12), .Z(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n917), .B2(new_n468), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n850), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n918), .B2(new_n921), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n800), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n850), .ZN(new_n928));
  INV_X1    g503(.A(new_n800), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n923), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n495), .A2(new_n500), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n926), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n908), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n931), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n924), .A2(new_n925), .A3(new_n800), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n929), .B1(new_n928), .B2(new_n923), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n939), .B(new_n932), .C1(new_n906), .C2(new_n907), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n481), .B(new_n657), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(G162), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  INV_X1    g520(.A(new_n943), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n935), .A2(new_n940), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g524(.A(new_n633), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT103), .B1(G299), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n576), .A2(G651), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n578), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n576), .A2(KEYINPUT72), .A3(G651), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n953), .A2(new_n954), .B1(G91), .B2(new_n540), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n955), .A2(new_n633), .A3(new_n956), .A4(new_n572), .ZN(new_n957));
  NAND2_X1  g532(.A1(G299), .A2(new_n950), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n951), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT41), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n572), .A3(new_n633), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n958), .A3(KEYINPUT41), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n958), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n641), .B(new_n894), .Z(new_n966));
  MUX2_X1   g541(.A(new_n964), .B(new_n965), .S(new_n966), .Z(new_n967));
  NOR2_X1   g542(.A1(G166), .A2(KEYINPUT104), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n969), .B(new_n511), .C1(new_n520), .C2(new_n527), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n832), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G303), .A2(new_n969), .ZN(new_n972));
  NAND2_X1  g547(.A1(G166), .A2(KEYINPUT104), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(G305), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n976));
  INV_X1    g551(.A(new_n609), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT77), .B1(new_n604), .B2(new_n605), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n976), .B(new_n619), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n610), .B2(new_n619), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n975), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n971), .A3(new_n974), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT42), .Z(new_n987));
  AND2_X1   g562(.A1(new_n967), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n967), .A2(new_n987), .ZN(new_n989));
  OAI21_X1  g564(.A(G868), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(G868), .B2(new_n902), .ZN(G295));
  OAI21_X1  g566(.A(new_n990), .B1(G868), .B2(new_n902), .ZN(G331));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n995));
  OAI21_X1  g570(.A(G168), .B1(new_n546), .B2(new_n550), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n541), .A2(new_n545), .A3(new_n539), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT70), .B1(new_n549), .B2(new_n544), .ZN(new_n998));
  NAND3_X1  g573(.A1(G286), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n894), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(new_n999), .A3(new_n889), .A4(new_n893), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n961), .A2(new_n1003), .A3(new_n963), .ZN(new_n1004));
  INV_X1    g579(.A(new_n965), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n995), .B(new_n945), .C1(new_n1007), .C2(new_n986), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1004), .A2(new_n1006), .B1(new_n985), .B2(new_n984), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n945), .B1(new_n1007), .B2(new_n986), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT105), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n994), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1000), .A2(new_n894), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n999), .A2(new_n996), .B1(new_n889), .B2(new_n893), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT41), .B(new_n959), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(new_n985), .A3(new_n984), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n965), .B1(new_n1003), .B2(KEYINPUT41), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n945), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1020), .A2(KEYINPUT43), .A3(new_n1009), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n993), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT43), .B1(new_n1020), .B2(new_n1009), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT106), .B(KEYINPUT43), .C1(new_n1020), .C2(new_n1009), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1011), .A2(new_n994), .A3(new_n1013), .ZN(new_n1028));
  AND4_X1   g603(.A1(KEYINPUT107), .A2(new_n1027), .A3(KEYINPUT44), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n993), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT107), .B1(new_n1030), .B2(new_n1028), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1022), .B1(new_n1029), .B2(new_n1031), .ZN(G397));
  OAI211_X1 g607(.A(new_n955), .B(new_n572), .C1(KEYINPUT117), .C2(KEYINPUT57), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT117), .B(new_n573), .C1(new_n577), .C2(new_n579), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n1035));
  NAND3_X1  g610(.A1(G299), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n493), .A2(new_n494), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n497), .A2(KEYINPUT68), .A3(new_n499), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT68), .B1(new_n497), .B2(new_n499), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G40), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n479), .B2(G2105), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n471), .A2(new_n473), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n495), .B2(new_n500), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT50), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1046), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n817), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G1384), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n495), .B2(new_n500), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(new_n471), .A3(new_n473), .A4(new_n1048), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1054), .B1(G164), .B2(G1384), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1037), .B1(new_n1053), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1053), .A2(new_n1037), .A3(new_n1061), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1063), .A2(new_n634), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1065));
  INV_X1    g640(.A(new_n500), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1384), .B1(new_n1040), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT109), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1044), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT109), .B1(new_n1050), .B2(KEYINPUT50), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1065), .A2(new_n1069), .A3(new_n1070), .A4(new_n1049), .ZN(new_n1071));
  INV_X1    g646(.A(G2067), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n471), .A2(new_n473), .A3(new_n1048), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n1050), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1071), .A2(new_n790), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1062), .B1(new_n1064), .B2(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n634), .A2(KEYINPUT60), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n634), .A2(KEYINPUT60), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1075), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT61), .B1(new_n1062), .B2(KEYINPUT121), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1053), .A2(new_n1061), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1037), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1063), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n1063), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1082), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT45), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1092), .A2(new_n1057), .A3(G1996), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(G1341), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1074), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n561), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1091), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1102), .A3(new_n1099), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT120), .B1(new_n1097), .B2(KEYINPUT59), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1100), .A2(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1077), .B1(new_n1090), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G8), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G168), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT51), .B1(new_n1108), .B2(KEYINPUT122), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1065), .A2(new_n1070), .A3(new_n1069), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1073), .A2(G2084), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1055), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(G164), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1043), .A2(KEYINPUT115), .A3(new_n1055), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1115), .A2(new_n1049), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1966), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1111), .A2(new_n1112), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1109), .B(new_n1110), .C1(new_n1120), .C2(new_n1107), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1110), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1112), .A2(new_n1065), .A3(new_n1070), .A4(new_n1069), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(G8), .B(new_n1122), .C1(new_n1125), .C2(G286), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1121), .A2(new_n1126), .B1(new_n1108), .B2(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(G2078), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1058), .A2(new_n1128), .A3(new_n1059), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1071), .A2(new_n728), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1128), .A2(KEYINPUT53), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n936), .B2(new_n1055), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1049), .A3(new_n1116), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1130), .A2(new_n1129), .B1(new_n1071), .B2(new_n728), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1118), .A2(new_n1133), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(G301), .A3(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1137), .A2(new_n1140), .A3(KEYINPUT54), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n823), .B1(new_n1092), .B2(new_n1057), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT110), .B(G2090), .Z(new_n1143));
  OAI21_X1  g718(.A(new_n1142), .B1(new_n1052), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G8), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G166), .A2(new_n1107), .ZN(new_n1146));
  NOR2_X1   g721(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1142), .B1(new_n1071), .B2(new_n1143), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(new_n1151), .A3(G8), .ZN(new_n1155));
  INV_X1    g730(.A(G1981), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1156), .B(new_n592), .C1(new_n597), .C2(new_n602), .ZN(new_n1157));
  OAI21_X1  g732(.A(G1981), .B1(new_n827), .B2(new_n830), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(KEYINPUT49), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT113), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT49), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT113), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1157), .A2(new_n1164), .A3(KEYINPUT49), .A4(new_n1158), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1074), .A2(new_n1107), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1160), .A2(new_n1163), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n590), .A2(G1976), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1168), .B(G8), .C1(new_n1073), .C2(new_n1050), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT52), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(KEYINPUT112), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(G1976), .ZN(new_n1174));
  NAND3_X1  g749(.A1(G288), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1153), .A2(new_n1155), .A3(new_n1167), .A4(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1127), .A2(new_n1141), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  AOI21_X1  g755(.A(G301), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1181));
  AND4_X1   g756(.A1(G301), .A2(new_n1131), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g760(.A(KEYINPUT123), .B(new_n1180), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1106), .A2(new_n1179), .A3(new_n1187), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1167), .A2(new_n1177), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1189), .A2(new_n1181), .A3(new_n1155), .A4(new_n1153), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1127), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1125), .A2(new_n1108), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1195), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1127), .B2(new_n1191), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1192), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1167), .A2(new_n1177), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT114), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT114), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1167), .A2(new_n1202), .A3(new_n1177), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1155), .ZN(new_n1205));
  INV_X1    g780(.A(G288), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1167), .A2(new_n1174), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1157), .ZN(new_n1208));
  AOI22_X1  g783(.A1(new_n1204), .A2(new_n1205), .B1(new_n1166), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT116), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1203), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1202), .B1(new_n1167), .B2(new_n1177), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1154), .A2(G8), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(new_n1152), .ZN(new_n1215));
  AOI211_X1 g790(.A(new_n1107), .B(G286), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1215), .A2(new_n1216), .A3(KEYINPUT63), .A4(new_n1155), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1210), .B1(new_n1213), .B2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1125), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1205), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1204), .A2(KEYINPUT116), .A3(new_n1215), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1216), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1222), .B1(new_n1178), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1218), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1188), .A2(new_n1199), .A3(new_n1209), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n800), .A2(new_n1072), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n929), .A2(G2067), .ZN(new_n1228));
  OAI211_X1 g803(.A(new_n1227), .B(new_n1228), .C1(new_n773), .C2(G1996), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n1116), .A2(new_n1073), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1230), .A2(G1996), .A3(new_n769), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT108), .ZN(new_n1232));
  OR2_X1    g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1234));
  AOI22_X1  g809(.A1(new_n1229), .A2(new_n1230), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g810(.A(new_n850), .B(new_n856), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1230), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g813(.A(G290), .B(G1986), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1238), .B1(new_n1230), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1226), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1242));
  INV_X1    g817(.A(new_n1230), .ZN(new_n1243));
  NOR2_X1   g818(.A1(new_n851), .A2(new_n856), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1235), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g820(.A(new_n1243), .B1(new_n1245), .B2(new_n1227), .ZN(new_n1246));
  INV_X1    g821(.A(KEYINPUT125), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1228), .A2(new_n1227), .ZN(new_n1249));
  OAI21_X1  g824(.A(new_n1230), .B1(new_n1249), .B2(new_n769), .ZN(new_n1250));
  NOR3_X1   g825(.A1(new_n1243), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1251));
  INV_X1    g826(.A(KEYINPUT46), .ZN(new_n1252));
  INV_X1    g827(.A(G1996), .ZN(new_n1253));
  AOI21_X1  g828(.A(new_n1252), .B1(new_n1230), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g829(.A(new_n1250), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g830(.A(new_n1255), .B(KEYINPUT47), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1248), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g832(.A(KEYINPUT126), .ZN(new_n1258));
  AOI21_X1  g833(.A(new_n1258), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1259));
  NOR3_X1   g834(.A1(new_n1243), .A2(G1986), .A3(G290), .ZN(new_n1260));
  XOR2_X1   g835(.A(new_n1260), .B(KEYINPUT48), .Z(new_n1261));
  OAI21_X1  g836(.A(new_n1261), .B1(new_n1238), .B2(KEYINPUT126), .ZN(new_n1262));
  OAI22_X1  g837(.A1(new_n1259), .A2(new_n1262), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1263));
  OAI21_X1  g838(.A(new_n1242), .B1(new_n1257), .B2(new_n1263), .ZN(new_n1264));
  OR2_X1    g839(.A1(new_n1262), .A2(new_n1259), .ZN(new_n1265));
  AND2_X1   g840(.A1(new_n1245), .A2(new_n1227), .ZN(new_n1266));
  OAI21_X1  g841(.A(KEYINPUT125), .B1(new_n1266), .B2(new_n1243), .ZN(new_n1267));
  INV_X1    g842(.A(new_n1256), .ZN(new_n1268));
  AOI21_X1  g843(.A(new_n1268), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1269));
  NAND4_X1  g844(.A1(new_n1265), .A2(new_n1267), .A3(new_n1269), .A4(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g845(.A1(new_n1264), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g846(.A1(new_n1241), .A2(new_n1271), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g847(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1274));
  OAI211_X1 g848(.A(new_n693), .B(G319), .C1(new_n674), .C2(new_n673), .ZN(new_n1275));
  AOI21_X1  g849(.A(new_n1275), .B1(new_n723), .B2(new_n724), .ZN(new_n1276));
  AND3_X1   g850(.A1(new_n1274), .A2(new_n1276), .A3(new_n948), .ZN(G308));
  NAND3_X1  g851(.A1(new_n1274), .A2(new_n1276), .A3(new_n948), .ZN(G225));
endmodule


