//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT65), .Z(new_n231));
  OAI21_X1  g0031(.A(new_n220), .B1(KEYINPUT1), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  OR2_X1    g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(G1698), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n254), .B1(new_n255), .B2(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(new_n263), .A3(G274), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G179), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n265), .A2(new_n273), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n207), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(G20), .B2(new_n203), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n213), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n285), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n206), .A2(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G50), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(G50), .B2(new_n288), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n276), .A2(G169), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n275), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G244), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n269), .B1(new_n296), .B2(new_n272), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n253), .A2(G232), .ZN(new_n298));
  INV_X1    g0098(.A(G107), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n298), .B1(new_n299), .B2(new_n258), .C1(new_n223), .C2(new_n260), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n297), .B1(new_n300), .B2(new_n264), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G20), .A2(G77), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT15), .B(G87), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n304), .B1(new_n277), .B2(new_n281), .C1(new_n278), .C2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n306), .A2(new_n285), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n290), .A2(G77), .A3(new_n291), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G77), .B2(new_n288), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n303), .B(new_n311), .C1(G169), .C2(new_n301), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n300), .A2(new_n264), .ZN(new_n313));
  INV_X1    g0113(.A(new_n297), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(G190), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n310), .C1(new_n316), .C2(new_n301), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n287), .A2(new_n293), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n319), .B(KEYINPUT9), .Z(new_n320));
  NAND2_X1  g0120(.A1(new_n274), .A2(G200), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n276), .A2(G190), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT10), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT10), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n320), .A2(new_n321), .A3(new_n325), .A4(new_n322), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n295), .B(new_n318), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n277), .B1(new_n206), .B2(G20), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n290), .B1(new_n289), .B2(new_n277), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT68), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT16), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT7), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n258), .B2(G20), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n222), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G58), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n222), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n338), .B2(new_n201), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n280), .A2(G159), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n332), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT7), .B1(new_n252), .B2(new_n207), .ZN(new_n343));
  NOR4_X1   g0143(.A1(new_n250), .A2(new_n251), .A3(new_n333), .A4(G20), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n345), .A2(KEYINPUT16), .A3(new_n339), .A4(new_n340), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n346), .A3(new_n285), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n270), .A2(G1698), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n348), .B1(G223), .B2(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G87), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n263), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n269), .B1(new_n235), .B2(new_n272), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n316), .B1(new_n351), .B2(new_n354), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT17), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n331), .A2(new_n347), .A3(new_n358), .A4(new_n361), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n331), .A2(new_n347), .A3(new_n358), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT69), .B(KEYINPUT17), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT18), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n331), .A2(new_n347), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n352), .B2(new_n355), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n351), .A2(new_n354), .A3(new_n302), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n366), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n371), .B1(new_n347), .B2(new_n331), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n366), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n365), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT14), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT13), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n235), .A2(G1698), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n381), .B1(G226), .B2(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n264), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n269), .B1(new_n223), .B2(new_n272), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n380), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n263), .B1(new_n382), .B2(new_n383), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n389), .A2(new_n386), .A3(KEYINPUT13), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n379), .B(G169), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n380), .A2(KEYINPUT66), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n385), .B2(new_n387), .ZN(new_n393));
  INV_X1    g0193(.A(new_n392), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n389), .A2(new_n386), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(G179), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT67), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n385), .A2(new_n387), .A3(new_n380), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT13), .B1(new_n389), .B2(new_n386), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n368), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n401), .B2(new_n379), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n388), .B2(new_n390), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT67), .A3(KEYINPUT14), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n397), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n289), .A2(new_n222), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT12), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n255), .B2(new_n278), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n290), .A2(G68), .A3(new_n291), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT11), .B1(new_n410), .B2(new_n285), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(G200), .B1(new_n388), .B2(new_n390), .ZN(new_n418));
  OAI21_X1  g0218(.A(G190), .B1(new_n393), .B2(new_n395), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(new_n415), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n327), .A2(new_n378), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT70), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT70), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n327), .A2(new_n424), .A3(new_n378), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G283), .ZN(new_n427));
  INV_X1    g0227(.A(G97), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(new_n207), .C1(G33), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G116), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G20), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n285), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT20), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n206), .A2(G33), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n288), .A2(new_n435), .A3(new_n213), .A4(new_n284), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n289), .A2(KEYINPUT76), .A3(new_n430), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT76), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n288), .B2(G116), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n437), .A2(G116), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(G264), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n443));
  INV_X1    g0243(.A(G1698), .ZN(new_n444));
  OAI211_X1 g0244(.A(G257), .B(new_n444), .C1(new_n250), .C2(new_n251), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n256), .A2(G303), .A3(new_n257), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n302), .B1(new_n447), .B2(new_n264), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n206), .B(G45), .C1(new_n266), .C2(KEYINPUT5), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(KEYINPUT71), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT71), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n267), .A2(G1), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G41), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(G270), .B(new_n263), .C1(new_n452), .C2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT75), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n263), .A2(G274), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n451), .A2(KEYINPUT71), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n454), .A2(new_n453), .A3(new_n456), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n450), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n458), .A2(new_n463), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT75), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n449), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT77), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n447), .A2(new_n264), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n466), .B2(new_n464), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n442), .A2(KEYINPUT21), .A3(G169), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n459), .B1(new_n458), .B2(new_n463), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT21), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n477), .B(new_n368), .C1(new_n434), .C2(new_n441), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT77), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n467), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT78), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n442), .A2(G169), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n471), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n476), .A2(KEYINPUT78), .A3(G169), .A4(new_n442), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n477), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n442), .B1(new_n476), .B2(G200), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n353), .B2(new_n476), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n480), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(G244), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n489));
  OAI211_X1 g0289(.A(G238), .B(new_n444), .C1(new_n250), .C2(new_n251), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G116), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n264), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n225), .B1(new_n267), .B2(G1), .ZN(new_n494));
  INV_X1    g0294(.A(G274), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n206), .A2(new_n495), .A3(G45), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n263), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n368), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n492), .B2(new_n264), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n302), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT19), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n207), .B1(new_n383), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G97), .A2(G107), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n224), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n207), .B(G68), .C1(new_n250), .C2(new_n251), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n503), .B1(new_n278), .B2(new_n428), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n285), .B1(new_n289), .B2(new_n305), .ZN(new_n511));
  INV_X1    g0311(.A(new_n305), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n437), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n500), .A2(new_n502), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT73), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n437), .A2(new_n516), .A3(G87), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT73), .B1(new_n436), .B2(new_n224), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n511), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n316), .B1(new_n493), .B2(new_n498), .ZN(new_n521));
  AOI211_X1 g0321(.A(new_n353), .B(new_n497), .C1(new_n492), .C2(new_n264), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT74), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT72), .ZN(new_n525));
  OAI21_X1  g0325(.A(G107), .B1(new_n343), .B2(new_n344), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  AND2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n505), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n299), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n286), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n288), .A2(G97), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n437), .B2(G97), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n525), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(G20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n280), .A2(G77), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n299), .B1(new_n334), .B2(new_n335), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n285), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(KEYINPUT72), .A3(new_n535), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(new_n263), .C1(new_n452), .C2(new_n457), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n544), .A2(new_n463), .ZN(new_n545));
  OAI211_X1 g0345(.A(G244), .B(new_n444), .C1(new_n250), .C2(new_n251), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n444), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n427), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n264), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n545), .A2(G179), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n368), .B1(new_n545), .B2(new_n552), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n537), .B(new_n543), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n499), .A2(G200), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n501), .A2(G190), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n556), .A2(new_n511), .A3(new_n557), .A4(new_n519), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT74), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n500), .A2(new_n502), .A3(new_n514), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n533), .A2(new_n536), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n545), .A2(G190), .A3(new_n552), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n544), .A2(new_n463), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n264), .B2(new_n551), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n562), .B(new_n563), .C1(new_n565), .C2(new_n316), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n524), .A2(new_n555), .A3(new_n561), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n289), .A2(new_n299), .ZN(new_n568));
  NOR2_X1   g0368(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n568), .B2(new_n569), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n570), .A2(new_n572), .B1(G107), .B2(new_n437), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n207), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT22), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n258), .A2(new_n577), .A3(new_n207), .A4(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n278), .A2(new_n430), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT79), .B1(new_n207), .B2(G107), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT23), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT23), .ZN(new_n583));
  OAI211_X1 g0383(.A(KEYINPUT79), .B(new_n583), .C1(new_n207), .C2(G107), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT24), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT24), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n579), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n574), .B1(new_n590), .B2(new_n285), .ZN(new_n591));
  OAI211_X1 g0391(.A(G264), .B(new_n263), .C1(new_n452), .C2(new_n457), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT82), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n461), .A2(new_n450), .A3(new_n462), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT82), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(G264), .A4(new_n263), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n258), .A2(G257), .A3(G1698), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n258), .A2(G250), .A3(new_n444), .ZN(new_n598));
  INV_X1    g0398(.A(G33), .ZN(new_n599));
  AND2_X1   g0399(.A1(KEYINPUT81), .A2(G294), .ZN(new_n600));
  NOR2_X1   g0400(.A1(KEYINPUT81), .A2(G294), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n593), .A2(new_n596), .B1(new_n264), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(G200), .B1(new_n604), .B2(new_n463), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n264), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n592), .A3(new_n463), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n591), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n593), .A2(new_n596), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(G179), .A3(new_n463), .A4(new_n606), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(G169), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n579), .A2(new_n588), .A3(new_n585), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n588), .B1(new_n579), .B2(new_n585), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n285), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n573), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n567), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n426), .A2(new_n488), .A3(new_n620), .ZN(G372));
  AND3_X1   g0421(.A1(new_n367), .A2(new_n372), .A3(new_n366), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(new_n373), .ZN(new_n623));
  INV_X1    g0423(.A(new_n312), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n406), .A2(new_n416), .B1(new_n420), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n365), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n324), .A2(new_n326), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n295), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n426), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n542), .A2(new_n535), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n553), .B2(new_n554), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT83), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n499), .A2(new_n635), .A3(new_n368), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT83), .B1(new_n501), .B2(G169), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n514), .A2(new_n502), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n523), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  OAI211_X1 g0441(.A(KEYINPUT85), .B(new_n631), .C1(new_n553), .C2(new_n554), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n634), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n638), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n555), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n641), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT84), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n640), .A2(new_n555), .A3(new_n566), .ZN(new_n653));
  INV_X1    g0453(.A(new_n609), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n545), .A2(new_n552), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G169), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n302), .B2(new_n656), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n537), .A2(new_n543), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n316), .B1(new_n545), .B2(new_n552), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n631), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n658), .A2(new_n659), .B1(new_n563), .B2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n662), .A2(KEYINPUT84), .A3(new_n609), .A4(new_n640), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n480), .A2(new_n485), .A3(new_n618), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n655), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n651), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n629), .B1(new_n630), .B2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(G213), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n442), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n488), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n480), .A2(new_n485), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n677), .B2(new_n674), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n673), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n591), .A2(new_n680), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n619), .A2(new_n681), .B1(new_n618), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT86), .Z(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n677), .A2(new_n673), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n611), .A2(new_n612), .B1(new_n616), .B2(new_n573), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n680), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n684), .A2(new_n686), .A3(new_n688), .ZN(G399));
  NOR2_X1   g0489(.A1(new_n506), .A2(G116), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT87), .ZN(new_n691));
  INV_X1    g0491(.A(new_n210), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n691), .A2(new_n693), .A3(new_n206), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n217), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  AOI21_X1  g0496(.A(new_n673), .B1(new_n651), .B2(new_n665), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n648), .A2(new_n649), .A3(new_n641), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n634), .A2(new_n640), .A3(new_n642), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n698), .B(new_n644), .C1(new_n699), .C2(new_n641), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n653), .A2(new_n654), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(new_n664), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n680), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  MUX2_X1   g0503(.A(new_n697), .B(new_n703), .S(KEYINPUT29), .Z(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n610), .A2(new_n463), .A3(new_n606), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n316), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n607), .A2(G190), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n687), .B1(new_n709), .B2(new_n591), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n648), .A3(new_n662), .A4(new_n680), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n480), .A2(new_n485), .A3(new_n487), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT89), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT89), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n488), .A2(new_n620), .A3(new_n714), .A4(new_n680), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n466), .A2(new_n464), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n448), .A2(new_n501), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n717), .A2(new_n565), .A3(new_n604), .A4(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n718), .B1(new_n466), .B2(new_n464), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n545), .A2(KEYINPUT30), .A3(new_n552), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n604), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n501), .A2(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n476), .A2(new_n706), .A3(new_n656), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n680), .B1(new_n728), .B2(KEYINPUT88), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT88), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n722), .A2(new_n730), .A3(new_n725), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n680), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n732), .A2(new_n733), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n705), .B1(new_n716), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n704), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n696), .B1(new_n737), .B2(G1), .ZN(G364));
  AND2_X1   g0538(.A1(new_n207), .A2(G13), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G45), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(G1), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n693), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n692), .A2(new_n252), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G355), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G116), .B2(new_n210), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n692), .A2(new_n258), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n267), .B2(new_n217), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n245), .A2(new_n267), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(G20), .B1(KEYINPUT91), .B2(G169), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(KEYINPUT91), .A2(G169), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n213), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n744), .B1(new_n752), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT92), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n207), .A2(G179), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G159), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NAND2_X1  g0569(.A1(G20), .A2(G179), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(new_n353), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n769), .B1(G68), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n771), .A2(new_n765), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n258), .B1(new_n775), .B2(new_n255), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n770), .A2(new_n353), .A3(G200), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(G58), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n771), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n353), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G50), .A2(new_n780), .B1(new_n782), .B2(G87), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n764), .A2(new_n353), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n299), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n353), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n207), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(G97), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n774), .A2(new_n778), .A3(new_n783), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n252), .B1(new_n775), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n777), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n792), .B(new_n795), .C1(G329), .C2(new_n767), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G326), .A2(new_n780), .B1(new_n782), .B2(G303), .ZN(new_n797));
  INV_X1    g0597(.A(new_n602), .ZN(new_n798));
  INV_X1    g0598(.A(new_n784), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n788), .A2(new_n798), .B1(new_n799), .B2(G283), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n772), .B1(new_n802), .B2(KEYINPUT93), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(KEYINPUT93), .B2(new_n802), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n790), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n756), .ZN(new_n807));
  INV_X1    g0607(.A(new_n759), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n763), .B1(new_n806), .B2(new_n807), .C1(new_n678), .C2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n678), .A2(G330), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n679), .A2(new_n811), .A3(new_n744), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  NAND2_X1  g0614(.A1(new_n311), .A2(new_n673), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n312), .A2(new_n317), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT96), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT96), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n312), .A2(new_n317), .A3(new_n818), .A4(new_n815), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n624), .A2(new_n673), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OR3_X1    g0621(.A1(new_n697), .A2(KEYINPUT97), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT97), .B1(new_n697), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n817), .A2(new_n819), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n697), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n822), .A2(new_n736), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT98), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n716), .A2(new_n735), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G330), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n744), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n757), .ZN(new_n834));
  INV_X1    g0634(.A(new_n744), .ZN(new_n835));
  INV_X1    g0635(.A(new_n775), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n836), .A2(G159), .B1(G143), .B2(new_n777), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  INV_X1    g0638(.A(new_n780), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n279), .B2(new_n772), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n784), .A2(new_n222), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n252), .B(new_n844), .C1(G132), .C2(new_n767), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n788), .A2(G58), .B1(new_n782), .B2(G50), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n842), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G303), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n839), .A2(new_n848), .B1(new_n781), .B2(new_n299), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G87), .B2(new_n799), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n258), .B1(G294), .B2(new_n777), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G311), .A2(new_n767), .B1(new_n836), .B2(G116), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT95), .B(G283), .Z(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n788), .A2(G97), .B1(new_n854), .B2(new_n773), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n807), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n756), .A2(new_n757), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n835), .B(new_n857), .C1(new_n255), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n834), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n832), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G384));
  OR2_X1    g0662(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(G116), .A3(new_n214), .A4(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT36), .Z(new_n866));
  NOR3_X1   g0666(.A1(new_n216), .A2(new_n255), .A3(new_n338), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n867), .A2(KEYINPUT99), .B1(new_n202), .B2(G68), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n206), .B(G13), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n375), .A2(new_n363), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT101), .ZN(new_n874));
  INV_X1    g0674(.A(new_n671), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n367), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT37), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n671), .B1(new_n331), .B2(new_n347), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n878), .B2(new_n874), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n367), .A2(new_n372), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n331), .A2(new_n347), .A3(new_n358), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n879), .B1(new_n882), .B2(new_n878), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n876), .B1(new_n623), .B2(new_n365), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n872), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n347), .A2(new_n329), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n372), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n875), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n881), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n873), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(KEYINPUT38), .B(new_n894), .C1(new_n378), .C2(new_n889), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n886), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n889), .B1(new_n623), .B2(new_n365), .ZN(new_n899));
  AOI22_X1  g0699(.A1(KEYINPUT37), .A2(new_n890), .B1(new_n873), .B2(new_n892), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n872), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n898), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n417), .A2(new_n673), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n903), .A2(new_n905), .B1(new_n623), .B2(new_n875), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n312), .A2(new_n673), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n697), .B2(new_n824), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n404), .A2(new_n402), .ZN(new_n910));
  INV_X1    g0710(.A(new_n397), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n911), .A3(new_n420), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n415), .A2(new_n680), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT100), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n913), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n420), .B(new_n915), .C1(new_n405), .C2(new_n415), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT100), .B1(new_n912), .B2(new_n913), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n909), .A2(new_n902), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n906), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n426), .A2(new_n704), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n629), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n922), .B(new_n924), .Z(new_n925));
  AND2_X1   g0725(.A1(new_n720), .A2(new_n721), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n727), .A2(new_n725), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT88), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND4_X1   g0728(.A1(KEYINPUT31), .A2(new_n928), .A3(new_n673), .A4(new_n731), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT31), .B1(new_n729), .B2(new_n731), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n716), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n630), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n821), .B1(new_n917), .B2(new_n918), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n713), .A2(new_n715), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n732), .A2(new_n733), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n731), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n936), .B(new_n902), .C1(new_n937), .C2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n886), .B2(new_n895), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n932), .A2(new_n944), .A3(new_n936), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n705), .B1(new_n934), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n934), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n925), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n206), .B2(new_n739), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n925), .A2(new_n948), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n871), .B1(new_n950), .B2(new_n951), .ZN(G367));
  NOR2_X1   g0752(.A1(new_n632), .A2(new_n680), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT103), .Z(new_n954));
  OAI21_X1  g0754(.A(new_n662), .B1(new_n562), .B2(new_n680), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n683), .A2(new_n685), .A3(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n958));
  INV_X1    g0758(.A(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n555), .B1(new_n959), .B2(new_n618), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n680), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n520), .A2(new_n673), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n640), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n644), .B2(new_n964), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT102), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n968), .B(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n684), .A2(new_n959), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n693), .B(KEYINPUT41), .Z(new_n976));
  NAND2_X1  g0776(.A1(new_n686), .A2(new_n688), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n959), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n686), .A2(new_n688), .A3(new_n956), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n982), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n683), .B(new_n685), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(new_n679), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n737), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n981), .B1(new_n979), .B2(new_n985), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n987), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n976), .B1(new_n993), .B2(new_n737), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n975), .B1(new_n994), .B2(new_n743), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n761), .B1(new_n692), .B2(new_n512), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n748), .A2(new_n241), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n835), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n781), .A2(new_n430), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n999), .A2(KEYINPUT46), .B1(new_n602), .B2(new_n772), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT46), .B2(new_n999), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1002), .A2(KEYINPUT106), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(KEYINPUT106), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n258), .B1(new_n767), .B2(G317), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n848), .B2(new_n793), .C1(new_n775), .C2(new_n853), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n788), .A2(G107), .B1(new_n799), .B2(G97), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n791), .B2(new_n839), .ZN(new_n1008));
  NOR4_X1   g0808(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT107), .Z(new_n1010));
  INV_X1    g0810(.A(G143), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n839), .A2(new_n1011), .B1(new_n784), .B2(new_n255), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n258), .B1(new_n775), .B2(new_n202), .C1(new_n793), .C2(new_n279), .ZN(new_n1013));
  INV_X1    g0813(.A(G159), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n787), .A2(new_n222), .B1(new_n772), .B2(new_n1014), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n781), .A2(new_n337), .B1(new_n766), .B2(new_n838), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT108), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1010), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  OAI221_X1 g0820(.A(new_n998), .B1(new_n808), .B2(new_n966), .C1(new_n1020), .C2(new_n807), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n995), .A2(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n989), .A2(new_n743), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n238), .A2(new_n267), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1024), .A2(new_n748), .B1(new_n691), .B2(new_n745), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n277), .A2(G50), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT50), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n267), .B1(new_n222), .B2(new_n255), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n691), .B(new_n1028), .C1(new_n1027), .C2(new_n1026), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1025), .A2(new_n1029), .B1(G107), .B2(new_n210), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n835), .B1(new_n1030), .B2(new_n760), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n787), .A2(new_n305), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n255), .B2(new_n781), .C1(new_n277), .C2(new_n772), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n252), .B1(G50), .B2(new_n777), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n222), .B2(new_n775), .C1(new_n279), .C2(new_n766), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n839), .A2(new_n1014), .B1(new_n784), .B2(new_n428), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n788), .A2(new_n854), .B1(new_n782), .B2(new_n798), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n836), .A2(G303), .B1(G317), .B2(new_n777), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n791), .B2(new_n772), .C1(new_n794), .C2(new_n839), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT109), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT49), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n258), .B1(new_n767), .B2(G326), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n430), .B2(new_n784), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1045), .B2(KEYINPUT49), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1038), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1050), .A2(KEYINPUT110), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n756), .B1(new_n1050), .B2(KEYINPUT110), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1031), .B1(new_n683), .B2(new_n808), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n990), .A2(new_n693), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n989), .A2(new_n737), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1023), .B(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(G393));
  NAND3_X1  g0856(.A1(new_n980), .A2(new_n684), .A3(new_n986), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n679), .B(new_n683), .C1(new_n979), .C2(new_n985), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n743), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n749), .A2(new_n248), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n760), .B1(new_n428), .B2(new_n210), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n744), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n780), .A2(G150), .B1(G159), .B2(new_n777), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT51), .Z(new_n1064));
  OAI221_X1 g0864(.A(new_n258), .B1(new_n766), .B2(new_n1011), .C1(new_n277), .C2(new_n775), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n787), .A2(new_n255), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n784), .A2(new_n224), .B1(new_n772), .B2(new_n202), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G68), .C2(new_n782), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G294), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n252), .B1(new_n775), .B2(new_n1071), .C1(new_n794), .C2(new_n766), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n785), .B(new_n1072), .C1(new_n782), .C2(new_n854), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n787), .A2(new_n430), .B1(new_n772), .B2(new_n848), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT111), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT111), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n780), .A2(G317), .B1(G311), .B2(new_n777), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1070), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT112), .Z(new_n1081));
  AOI21_X1  g0881(.A(new_n1062), .B1(new_n1081), .B2(new_n756), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n956), .B2(new_n808), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n993), .A2(new_n693), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n991), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1059), .B(new_n1083), .C1(new_n1084), .C2(new_n1085), .ZN(G390));
  NOR2_X1   g0886(.A1(new_n933), .A2(new_n705), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n426), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n923), .A3(new_n629), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n705), .B(new_n833), .C1(new_n931), .C2(new_n716), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n920), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n680), .B(new_n824), .C1(new_n700), .C2(new_n702), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n907), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT113), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(KEYINPUT113), .A3(new_n1094), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n932), .A2(G330), .A3(new_n821), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(KEYINPUT114), .A3(new_n919), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n736), .A2(new_n936), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1092), .A2(new_n1098), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n919), .B1(new_n830), .B2(new_n833), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n932), .A2(G330), .A3(new_n936), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n909), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1089), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n905), .B1(new_n908), .B2(new_n919), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n903), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1097), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1111), .A2(new_n1095), .A3(new_n919), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n904), .B1(new_n886), .B2(new_n895), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1110), .B(new_n1101), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1096), .A2(new_n920), .A3(new_n1097), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1116), .A2(new_n1113), .B1(new_n1109), .B2(new_n903), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1117), .B2(new_n1104), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1108), .A2(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1117), .A2(new_n1104), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n1107), .A3(new_n1115), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1121), .A3(new_n693), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1120), .A2(KEYINPUT115), .A3(new_n743), .A4(new_n1115), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT115), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n743), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n903), .A2(new_n757), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n835), .B1(new_n277), .B2(new_n858), .ZN(new_n1129));
  INV_X1    g0929(.A(G132), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n793), .A2(new_n1130), .B1(new_n775), .B2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n788), .A2(G159), .B1(new_n773), .B2(G137), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n839), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1132), .B(new_n1135), .C1(G125), .C2(new_n767), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n781), .A2(new_n279), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT53), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n258), .B1(new_n784), .B2(new_n202), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1139), .A2(KEYINPUT116), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(KEYINPUT116), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n252), .B1(new_n781), .B2(new_n224), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT117), .Z(new_n1144));
  AOI22_X1  g0944(.A1(G294), .A2(new_n767), .B1(new_n836), .B2(G97), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n430), .B2(new_n793), .ZN(new_n1146));
  INV_X1    g0946(.A(G283), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n839), .A2(new_n1147), .B1(new_n299), .B2(new_n772), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1146), .A2(new_n1148), .A3(new_n844), .A4(new_n1067), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1136), .A2(new_n1142), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1128), .B(new_n1129), .C1(new_n807), .C2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1122), .A2(new_n1127), .A3(new_n1151), .ZN(G378));
  INV_X1    g0952(.A(new_n295), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n319), .B(new_n671), .C1(new_n628), .C2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n319), .A2(new_n671), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n295), .B(new_n1155), .C1(new_n324), .C2(new_n326), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n1154), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n945), .A2(G330), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n935), .B1(new_n931), .B2(new_n716), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT40), .B1(new_n1163), .B2(new_n902), .ZN(new_n1164));
  OAI21_X1  g0964(.A(KEYINPUT119), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n705), .B1(new_n1163), .B2(new_n944), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT119), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n943), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1161), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n943), .B2(new_n1166), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1161), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT120), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n922), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n922), .ZN(new_n1175));
  OAI211_X1 g0975(.A(KEYINPUT120), .B(new_n1175), .C1(new_n1169), .C2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1171), .A2(new_n757), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n858), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n744), .B1(new_n1179), .B2(G50), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n839), .A2(new_n430), .B1(new_n784), .B2(new_n337), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G97), .B2(new_n773), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n252), .A2(new_n266), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n793), .A2(new_n299), .B1(new_n766), .B2(new_n1147), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n512), .C2(new_n836), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n788), .A2(G68), .B1(new_n782), .B2(G77), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT58), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1183), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n780), .A2(G125), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1130), .B2(new_n772), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n836), .A2(G137), .B1(G128), .B2(new_n777), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n781), .B2(new_n1131), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(G150), .C2(new_n788), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n799), .A2(G159), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1188), .B(new_n1189), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT118), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n807), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1180), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1177), .A2(new_n743), .B1(new_n1178), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1089), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1101), .B1(new_n1111), .B2(new_n1095), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT114), .B1(new_n1099), .B2(new_n919), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1210), .A2(new_n1100), .B1(new_n909), .B2(new_n1105), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1207), .B1(new_n1118), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n922), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n943), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1171), .B1(new_n1215), .B2(new_n1170), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1165), .A2(new_n1161), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1175), .A3(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1212), .A2(KEYINPUT57), .A3(new_n1214), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n693), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1206), .B1(new_n1213), .B2(new_n1220), .ZN(G375));
  NAND2_X1  g1021(.A1(new_n919), .A2(new_n757), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n744), .B1(new_n1179), .B2(G68), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n781), .A2(new_n428), .B1(new_n766), .B2(new_n848), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT121), .Z(new_n1225));
  OAI221_X1 g1025(.A(new_n252), .B1(new_n775), .B2(new_n299), .C1(new_n793), .C2(new_n1147), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1033), .B1(new_n255), .B2(new_n784), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n839), .A2(new_n1071), .B1(new_n430), .B2(new_n772), .ZN(new_n1228));
  OR4_X1    g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n337), .A2(new_n784), .B1(new_n781), .B2(new_n1014), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n258), .B1(new_n775), .B2(new_n279), .C1(new_n1134), .C2(new_n766), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(G50), .C2(new_n788), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT122), .Z(new_n1233));
  NAND2_X1  g1033(.A1(new_n777), .A2(G137), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n772), .B2(new_n1131), .C1(new_n839), .C2(new_n1130), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1229), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1223), .B1(new_n1236), .B2(new_n756), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1222), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1211), .B2(new_n1125), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n976), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1102), .A2(new_n1106), .A3(new_n1089), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1108), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(G381));
  OR2_X1    g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(G390), .A2(new_n1245), .A3(G384), .A4(G381), .ZN(new_n1246));
  INV_X1    g1046(.A(G378), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1246), .A2(new_n1021), .A3(new_n995), .A4(new_n1247), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(G375), .ZN(G407));
  NAND2_X1  g1049(.A1(new_n672), .A2(G213), .ZN(new_n1250));
  OR3_X1    g1050(.A1(G375), .A2(G378), .A3(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(G407), .A2(G213), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT123), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT123), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(G407), .A2(new_n1254), .A3(G213), .A4(new_n1251), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(G409));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1250), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1214), .A2(new_n1218), .A3(new_n743), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1178), .A2(new_n1205), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1259), .A2(KEYINPUT124), .A3(new_n1260), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1175), .B1(new_n1265), .B2(KEYINPUT120), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1176), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1241), .B(new_n1212), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1263), .A2(new_n1264), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1247), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1206), .B(G378), .C1(new_n1213), .C2(new_n1220), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1258), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1258), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1106), .A2(new_n1102), .A3(new_n1089), .A4(KEYINPUT60), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1275), .A2(new_n693), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1242), .B1(new_n1107), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(G384), .A3(new_n1240), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1279), .B2(new_n1240), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1274), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1279), .A2(new_n1240), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n861), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1280), .A3(new_n1273), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1257), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1285), .A2(new_n1280), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n1258), .B(new_n1292), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1291), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(KEYINPUT126), .B(new_n1257), .C1(new_n1272), .C2(new_n1287), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1290), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1293), .A2(new_n1294), .A3(new_n1291), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(new_n813), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G390), .B1(new_n995), .B2(new_n1021), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n995), .A2(G390), .A3(new_n1021), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1302), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1299), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1304), .A2(new_n1300), .A3(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1298), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1292), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1250), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1293), .A2(KEYINPUT63), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1250), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1287), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT125), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1272), .A2(new_n1318), .A3(new_n1287), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1313), .B(new_n1314), .C1(new_n1317), .C2(new_n1319), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1297), .A2(new_n1308), .B1(new_n1320), .B2(new_n1307), .ZN(G405));
  XNOR2_X1  g1121(.A(G375), .B(G378), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1310), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(new_n1307), .ZN(G402));
endmodule


