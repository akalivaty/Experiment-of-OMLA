//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203));
  AOI21_X1  g002(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n204));
  OR2_X1    g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n207), .A2(KEYINPUT69), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT69), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n203), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT29), .ZN(new_n213));
  AND2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(G155gat), .B2(G162gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G141gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G155gat), .B(G162gat), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT2), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n220), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n212), .B1(new_n213), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n212), .A2(new_n235), .A3(new_n213), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n210), .A2(new_n211), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT81), .B1(new_n237), .B2(KEYINPUT29), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n231), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n234), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n212), .A2(new_n213), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n231), .B1(new_n244), .B2(new_n232), .ZN(new_n245));
  INV_X1    g044(.A(new_n242), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n245), .A2(new_n246), .A3(new_n234), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n202), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  INV_X1    g048(.A(new_n202), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n249), .B(new_n250), .C1(new_n242), .C2(new_n241), .ZN(new_n251));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G22gat), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n248), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n253), .B1(new_n248), .B2(new_n251), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT27), .B(G183gat), .ZN(new_n259));
  INV_X1    g058(.A(G190gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G183gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT27), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT27), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G183gat), .ZN(new_n265));
  AND4_X1   g064(.A1(new_n258), .A2(new_n263), .A3(new_n265), .A4(new_n260), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n257), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(new_n265), .A3(new_n260), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT64), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n259), .A2(new_n258), .A3(new_n260), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT28), .ZN(new_n271));
  INV_X1    g070(.A(G169gat), .ZN(new_n272));
  INV_X1    g071(.A(G176gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n274), .A2(KEYINPUT26), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(KEYINPUT26), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n262), .B2(new_n260), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n267), .A2(new_n271), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  NAND2_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(new_n260), .ZN(new_n283));
  OAI21_X1  g082(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n275), .A2(KEYINPUT23), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n288), .B2(new_n275), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n281), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n282), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n260), .B2(new_n282), .ZN(new_n292));
  INV_X1    g091(.A(new_n275), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n274), .B2(new_n287), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n294), .A4(new_n286), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G120gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT65), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G120gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n301), .A3(G113gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n298), .A2(G113gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT66), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT65), .B(G120gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n303), .B1(new_n307), .B2(G113gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT66), .ZN(new_n309));
  INV_X1    g108(.A(G134gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G127gat), .ZN(new_n311));
  INV_X1    g110(.A(G127gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G134gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n306), .A2(new_n309), .A3(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G113gat), .B(G120gat), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n314), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(new_n313), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n297), .B(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G227gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT32), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT33), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(G15gat), .B(G43gat), .Z(new_n330));
  XNOR2_X1  g129(.A(G71gat), .B(G99gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n332), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n326), .B(KEYINPUT32), .C1(new_n328), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT34), .B1(new_n325), .B2(KEYINPUT67), .ZN(new_n337));
  INV_X1    g136(.A(new_n323), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n337), .B1(new_n338), .B2(new_n324), .ZN(new_n339));
  INV_X1    g138(.A(new_n337), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n323), .A2(new_n325), .A3(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n339), .A2(new_n341), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(new_n333), .A3(new_n335), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT87), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT35), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(KEYINPUT87), .A3(new_n345), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n256), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT70), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n297), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n280), .A2(KEYINPUT70), .A3(new_n296), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT29), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT71), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n280), .A2(KEYINPUT70), .A3(new_n296), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT70), .B1(new_n280), .B2(new_n296), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n213), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT71), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n356), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n297), .A2(new_n357), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n358), .A2(new_n212), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n359), .A2(new_n360), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n357), .A2(KEYINPUT29), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n366), .A2(new_n357), .B1(new_n297), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n237), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G8gat), .B(G36gat), .Z(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT72), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n365), .A2(KEYINPUT30), .A3(new_n369), .A4(new_n374), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n365), .A2(new_n369), .A3(new_n374), .ZN(new_n379));
  XOR2_X1   g178(.A(KEYINPUT75), .B(KEYINPUT30), .Z(new_n380));
  AND2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT82), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n383), .A2(new_n376), .A3(new_n384), .A4(new_n377), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT0), .ZN(new_n388));
  XNOR2_X1  g187(.A(G57gat), .B(G85gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n322), .A2(new_n392), .A3(new_n233), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n316), .B1(new_n308), .B2(KEYINPUT66), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n302), .A2(KEYINPUT66), .A3(new_n304), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n231), .B(new_n321), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT4), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n398), .B2(KEYINPUT4), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(KEYINPUT77), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n317), .A2(new_n405), .A3(new_n231), .A4(new_n321), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT4), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n395), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n397), .A2(new_n305), .A3(new_n315), .ZN(new_n410));
  INV_X1    g209(.A(new_n321), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n240), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n412), .A3(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(new_n394), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n409), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n398), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n393), .B2(KEYINPUT4), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n404), .B2(new_n406), .ZN(new_n424));
  NOR4_X1   g223(.A1(new_n422), .A2(new_n424), .A3(KEYINPUT5), .A4(new_n414), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n391), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427));
  INV_X1    g226(.A(new_n402), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n400), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n394), .B(new_n393), .C1(new_n429), .C2(new_n407), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT78), .B1(new_n415), .B2(KEYINPUT5), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT5), .ZN(new_n432));
  AOI211_X1 g231(.A(new_n417), .B(new_n432), .C1(new_n413), .C2(new_n414), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n425), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n390), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n426), .A2(new_n427), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n390), .B1(new_n434), .B2(new_n435), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT6), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n351), .A2(new_n386), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n434), .A2(new_n390), .A3(new_n435), .ZN(new_n443));
  NOR2_X1   g242(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n443), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n438), .A2(new_n445), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n383), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n378), .A2(KEYINPUT74), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT74), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n376), .A2(new_n451), .A3(new_n377), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n442), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n336), .A2(KEYINPUT68), .A3(new_n342), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n342), .B1(new_n336), .B2(KEYINPUT68), .ZN(new_n456));
  NOR4_X1   g255(.A1(new_n254), .A2(new_n455), .A3(new_n255), .A4(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n376), .A2(new_n451), .A3(new_n377), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n451), .B1(new_n376), .B2(new_n377), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n426), .A2(new_n444), .A3(new_n436), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n381), .B1(new_n461), .B2(new_n447), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT80), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n454), .A2(new_n457), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n441), .B1(new_n464), .B2(KEYINPUT35), .ZN(new_n465));
  INV_X1    g264(.A(new_n256), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT80), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT80), .B1(new_n460), .B2(new_n462), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT36), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n455), .A2(new_n456), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT36), .B1(new_n343), .B2(new_n345), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n365), .A2(new_n474), .A3(new_n369), .ZN(new_n475));
  INV_X1    g274(.A(new_n374), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n365), .B2(new_n369), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT38), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n370), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT38), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n375), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n358), .A2(new_n237), .A3(new_n363), .A4(new_n364), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n474), .B1(new_n368), .B2(new_n212), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n480), .A2(new_n374), .B1(new_n485), .B2(new_n475), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n479), .A2(new_n486), .A3(new_n437), .A4(new_n439), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n487), .A2(new_n256), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n413), .A2(new_n414), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n490), .A2(KEYINPUT39), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n414), .B1(new_n422), .B2(new_n424), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n414), .B(new_n494), .C1(new_n422), .C2(new_n424), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n495), .A2(new_n496), .A3(new_n390), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n495), .B2(new_n390), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT86), .B1(KEYINPUT85), .B2(KEYINPUT40), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n500), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n493), .B(new_n502), .C1(new_n497), .C2(new_n498), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n426), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n386), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n473), .B1(new_n488), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n465), .B1(new_n469), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(G197gat), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT11), .B(G169gat), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT12), .Z(new_n514));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT89), .ZN(new_n516));
  AND2_X1   g315(.A1(G29gat), .A2(G36gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT88), .ZN(new_n518));
  NOR2_X1   g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n521), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n522), .A2(new_n523), .B1(new_n525), .B2(new_n515), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT16), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(G1gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G1gat), .B2(new_n528), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n527), .B2(KEYINPUT17), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(KEYINPUT18), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n527), .B(new_n533), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n539), .B(KEYINPUT13), .Z(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT18), .B1(new_n538), .B2(new_n539), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n514), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n545), .ZN(new_n547));
  INV_X1    g346(.A(new_n514), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n540), .A4(new_n543), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(KEYINPUT90), .B(new_n514), .C1(new_n544), .C2(new_n545), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  INV_X1    g356(.A(G92gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT94), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n555), .B1(new_n565), .B2(new_n527), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n537), .A2(new_n569), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT96), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G134gat), .B(G162gat), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n574), .B(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(G57gat), .A2(G64gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G57gat), .A2(G64gat), .ZN(new_n580));
  AND2_X1   g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(KEYINPUT9), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(new_n581), .ZN(new_n584));
  XNOR2_X1  g383(.A(G71gat), .B(G78gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n533), .B1(new_n586), .B2(new_n587), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT93), .ZN(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT92), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n592), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n565), .A2(new_n586), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n563), .A2(new_n564), .ZN(new_n604));
  INV_X1    g403(.A(new_n564), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n560), .B2(new_n562), .ZN(new_n606));
  OR3_X1    g405(.A1(new_n604), .A2(new_n586), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n565), .A2(KEYINPUT97), .A3(new_n586), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT10), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n602), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n602), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n615), .A3(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR4_X1   g424(.A1(new_n554), .A2(new_n578), .A3(new_n601), .A4(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n509), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n461), .A2(new_n447), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G1gat), .ZN(G1324gat));
  INV_X1    g430(.A(new_n627), .ZN(new_n632));
  INV_X1    g431(.A(new_n386), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT16), .B(G8gat), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n532), .B1(new_n627), .B2(new_n386), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT42), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(KEYINPUT42), .B2(new_n635), .ZN(G1325gat));
  OR2_X1    g437(.A1(new_n471), .A2(new_n472), .ZN(new_n639));
  OAI21_X1  g438(.A(G15gat), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n348), .A2(new_n350), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(G15gat), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n632), .B2(new_n642), .ZN(G1326gat));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n466), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT43), .B(G22gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  INV_X1    g445(.A(new_n577), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n574), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n649));
  INV_X1    g448(.A(new_n441), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n469), .A2(new_n507), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n554), .A2(new_n625), .A3(new_n600), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n628), .A2(G29gat), .ZN(new_n656));
  OR3_X1    g455(.A1(new_n655), .A2(KEYINPUT98), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT98), .B1(new_n655), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT45), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n661), .B(KEYINPUT44), .C1(new_n508), .C2(new_n648), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT99), .B1(new_n653), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n256), .B1(new_n454), .B2(new_n463), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n504), .B1(new_n382), .B2(new_n385), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n487), .A2(new_n256), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n639), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT100), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n469), .A2(new_n507), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n651), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n663), .A3(new_n578), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n648), .B1(new_n673), .B2(new_n651), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(KEYINPUT101), .A3(new_n663), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n665), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n654), .ZN(new_n681));
  OAI21_X1  g480(.A(G29gat), .B1(new_n681), .B2(new_n628), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n660), .A2(new_n682), .ZN(G1328gat));
  NOR3_X1   g482(.A1(new_n655), .A2(G36gat), .A3(new_n633), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT102), .ZN(new_n687));
  OAI21_X1  g486(.A(G36gat), .B1(new_n681), .B2(new_n633), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT103), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(G1329gat));
  INV_X1    g490(.A(G43gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n655), .B2(new_n641), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n473), .A2(G43gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n681), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT47), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n697), .B(new_n693), .C1(new_n681), .C2(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1330gat));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n653), .A2(new_n466), .A3(new_n654), .ZN(new_n701));
  INV_X1    g500(.A(G50gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n466), .A2(G50gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n681), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT48), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n703), .B(new_n707), .C1(new_n681), .C2(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1331gat));
  NOR2_X1   g508(.A1(new_n578), .A2(new_n601), .ZN(new_n710));
  AND4_X1   g509(.A1(new_n554), .A2(new_n674), .A3(new_n710), .A4(new_n625), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n628), .B(KEYINPUT105), .Z(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n386), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT49), .B(G64gat), .Z(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n715), .B2(new_n717), .ZN(G1333gat));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n473), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n641), .A2(G71gat), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n719), .A2(G71gat), .B1(new_n711), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g521(.A1(new_n711), .A2(new_n466), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g523(.A1(new_n553), .A2(new_n600), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n674), .A2(new_n578), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n678), .A2(KEYINPUT51), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n730), .A2(new_n557), .A3(new_n629), .A4(new_n625), .ZN(new_n731));
  INV_X1    g530(.A(new_n725), .ZN(new_n732));
  INV_X1    g531(.A(new_n625), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n664), .A2(new_n662), .B1(new_n675), .B2(new_n676), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n679), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n629), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n731), .B1(new_n738), .B2(new_n557), .ZN(G1336gat));
  NAND3_X1  g538(.A1(new_n680), .A2(new_n386), .A3(new_n734), .ZN(new_n740));
  AOI211_X1 g539(.A(KEYINPUT106), .B(KEYINPUT51), .C1(new_n678), .C2(new_n725), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT51), .B1(new_n678), .B2(new_n725), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n465), .B1(new_n670), .B2(new_n672), .ZN(new_n743));
  NOR4_X1   g542(.A1(new_n743), .A2(new_n727), .A3(new_n648), .A4(new_n732), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n741), .B1(new_n745), .B2(KEYINPUT106), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n633), .A2(G92gat), .A3(new_n733), .ZN(new_n747));
  AOI22_X1  g546(.A1(G92gat), .A2(new_n740), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n558), .B1(new_n737), .B2(new_n386), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n633), .A2(G92gat), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n730), .A2(new_n751), .A3(new_n625), .A4(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n625), .B(new_n752), .C1(new_n742), .C2(new_n744), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT107), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n755), .A3(new_n749), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n756), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n680), .A2(new_n473), .A3(new_n734), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n680), .A2(KEYINPUT108), .A3(new_n473), .A4(new_n734), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT109), .B(G99gat), .Z(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  OR4_X1    g563(.A1(new_n641), .A2(new_n745), .A3(new_n733), .A4(new_n763), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n680), .A2(new_n466), .A3(new_n734), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT110), .B(G106gat), .Z(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n733), .A2(G106gat), .A3(new_n256), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT111), .Z(new_n771));
  AOI21_X1  g570(.A(KEYINPUT53), .B1(new_n730), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n767), .A2(new_n768), .B1(new_n746), .B2(new_n771), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n611), .A2(new_n602), .A3(new_n613), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(KEYINPUT54), .A3(new_n614), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n621), .B1(new_n614), .B2(KEYINPUT54), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n781), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n783), .A2(KEYINPUT55), .A3(new_n779), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n553), .A2(new_n782), .A3(new_n623), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n538), .A2(new_n539), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n541), .A2(new_n542), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n513), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(new_n549), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n625), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n578), .B1(new_n785), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n783), .A2(new_n779), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n622), .B1(new_n794), .B2(new_n777), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n578), .A2(new_n795), .A3(new_n784), .A4(new_n791), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n601), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n710), .A2(KEYINPUT112), .A3(new_n554), .A4(new_n733), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n554), .A2(new_n648), .A3(new_n600), .A4(new_n733), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n804), .A2(new_n457), .A3(new_n712), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(new_n633), .ZN(new_n806));
  AOI21_X1  g605(.A(G113gat), .B1(new_n806), .B2(new_n553), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n641), .A2(new_n466), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n809), .A2(new_n628), .A3(new_n386), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n553), .A2(G113gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(G1340gat));
  AOI21_X1  g611(.A(new_n298), .B1(new_n810), .B2(new_n625), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT114), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n806), .A2(new_n307), .A3(new_n625), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1341gat));
  INV_X1    g615(.A(new_n810), .ZN(new_n817));
  OAI21_X1  g616(.A(G127gat), .B1(new_n817), .B2(new_n601), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n806), .A2(new_n312), .A3(new_n600), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1342gat));
  OAI21_X1  g619(.A(G134gat), .B1(new_n817), .B2(new_n648), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n648), .A2(new_n386), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n310), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n826));
  OAI221_X1 g625(.A(new_n821), .B1(KEYINPUT56), .B2(new_n823), .C1(new_n825), .C2(new_n826), .ZN(G1343gat));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT121), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT122), .Z(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n386), .A2(new_n628), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n639), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n804), .A2(new_n466), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT116), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837));
  AOI211_X1 g636(.A(new_n837), .B(KEYINPUT57), .C1(new_n804), .C2(new_n466), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n793), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n796), .B1(new_n793), .B2(new_n840), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT118), .B(new_n601), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n803), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n785), .A2(new_n792), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n648), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT117), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n796), .A3(new_n841), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT118), .B1(new_n849), .B2(new_n601), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT57), .B(new_n466), .C1(new_n845), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n833), .B1(new_n839), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n221), .B1(new_n852), .B2(new_n553), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n804), .A2(new_n712), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n473), .A2(new_n256), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT120), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n854), .B2(KEYINPUT119), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n855), .A2(new_n633), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n554), .A2(G141gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n828), .A2(KEYINPUT121), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n831), .B1(new_n853), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n862), .B1(new_n859), .B2(new_n860), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n554), .B(new_n833), .C1(new_n839), .C2(new_n851), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n866), .B(new_n830), .C1(new_n867), .C2(new_n221), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(G1344gat));
  NAND3_X1  g668(.A1(new_n859), .A2(new_n223), .A3(new_n625), .ZN(new_n870));
  AOI211_X1 g669(.A(KEYINPUT59), .B(new_n223), .C1(new_n852), .C2(new_n625), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n798), .A2(new_n800), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT123), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(KEYINPUT123), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n874), .A2(new_n835), .A3(new_n466), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n834), .A2(KEYINPUT57), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n833), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n625), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n872), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n870), .B1(new_n871), .B2(new_n881), .ZN(G1345gat));
  AOI21_X1  g681(.A(new_n227), .B1(new_n852), .B2(new_n600), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n601), .A2(G155gat), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n859), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT124), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n601), .B(new_n833), .C1(new_n839), .C2(new_n851), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n888), .B(new_n885), .C1(new_n889), .C2(new_n227), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(G1346gat));
  NAND4_X1  g690(.A1(new_n855), .A2(new_n858), .A3(new_n228), .A4(new_n822), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n852), .A2(new_n578), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n228), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n712), .A2(new_n633), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n804), .A2(new_n808), .A3(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(new_n272), .A3(new_n554), .ZN(new_n897));
  AOI211_X1 g696(.A(new_n629), .B(new_n633), .C1(new_n798), .C2(new_n803), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(new_n457), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n553), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(new_n272), .ZN(G1348gat));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n273), .A3(new_n625), .ZN(new_n902));
  OAI21_X1  g701(.A(G176gat), .B1(new_n896), .B2(new_n733), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1349gat));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n259), .A3(new_n600), .ZN(new_n905));
  OAI21_X1  g704(.A(G183gat), .B1(new_n896), .B2(new_n601), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n905), .A2(new_n906), .B1(KEYINPUT125), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n896), .B2(new_n648), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT61), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n899), .A2(new_n260), .A3(new_n578), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1351gat));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n856), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n553), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n639), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n876), .A2(new_n877), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n553), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  NAND3_X1  g721(.A1(new_n878), .A2(new_n625), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G204gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n915), .A2(G204gat), .A3(new_n733), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1353gat));
  OR3_X1    g726(.A1(new_n915), .A2(G211gat), .A3(new_n601), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n920), .A2(new_n600), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1354gat));
  AOI21_X1  g731(.A(G218gat), .B1(new_n916), .B2(new_n578), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n578), .A2(G218gat), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT126), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n920), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1355gat));
endmodule


