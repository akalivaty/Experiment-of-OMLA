//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n206), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n211), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n207), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n220), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AOI21_X1  g0050(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G238), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT66), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(G1), .B(G13), .C1(new_n259), .C2(new_n252), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT66), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n258), .A2(new_n260), .A3(new_n263), .A4(G274), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT13), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n235), .A2(G1698), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n267), .B(new_n268), .C1(G226), .C2(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G97), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n251), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n265), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n256), .A2(new_n264), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n260), .B1(new_n269), .B2(new_n270), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT13), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(new_n276), .A3(G179), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n266), .B1(new_n265), .B2(new_n272), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT13), .ZN(new_n279));
  OAI21_X1  g0079(.A(G169), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n280), .B2(KEYINPUT14), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT72), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT14), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n273), .B2(new_n276), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT72), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n281), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G68), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT12), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT67), .B1(new_n207), .B2(new_n259), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT67), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n294), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n293), .A2(new_n213), .A3(new_n295), .A4(new_n289), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n214), .A2(G1), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(G68), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n292), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n296), .A2(new_n222), .A3(new_n298), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT70), .B1(new_n291), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n214), .A2(G33), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n227), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n293), .A2(new_n213), .A3(new_n295), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(KEYINPUT11), .A3(new_n309), .ZN(new_n313));
  AND4_X1   g0113(.A1(new_n302), .A2(new_n304), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n288), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(G200), .B1(new_n278), .B2(new_n279), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n273), .A2(new_n276), .A3(G190), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT71), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n255), .A2(G244), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n264), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n267), .A2(G238), .A3(G1698), .ZN(new_n325));
  INV_X1    g0125(.A(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n267), .A2(G232), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n325), .B(new_n327), .C1(new_n229), .C2(new_n267), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n324), .B1(new_n251), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G20), .A2(G77), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  INV_X1    g0133(.A(new_n305), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT15), .B(G87), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n332), .B1(new_n333), .B2(new_n334), .C1(new_n307), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n289), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n336), .A2(new_n309), .B1(new_n227), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n297), .A2(G77), .A3(new_n299), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n331), .B(new_n340), .C1(G169), .C2(new_n329), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n299), .A2(G50), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n296), .A2(new_n342), .B1(G50), .B2(new_n289), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n305), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n333), .A2(KEYINPUT68), .ZN(new_n345));
  INV_X1    g0145(.A(G58), .ZN(new_n346));
  OR3_X1    g0146(.A1(new_n346), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n348), .B2(new_n307), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n309), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n343), .B1(new_n350), .B2(KEYINPUT69), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(KEYINPUT69), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G222), .A2(G1698), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n326), .A2(G223), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n267), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n251), .C1(G77), .C2(new_n267), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n255), .A2(G226), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n264), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n284), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G179), .B2(new_n360), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n340), .B1(new_n329), .B2(G190), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n329), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n322), .A2(new_n341), .A3(new_n363), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n360), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n352), .A2(KEYINPUT9), .A3(new_n353), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT9), .ZN(new_n373));
  INV_X1    g0173(.A(new_n353), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(new_n351), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n371), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT9), .B1(new_n352), .B2(new_n353), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n351), .A3(new_n373), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT10), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(new_n371), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n315), .B(new_n367), .C1(new_n377), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n309), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G33), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n385), .B1(new_n214), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n391), .B(G20), .C1(new_n386), .C2(new_n388), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n346), .A2(new_n222), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n394), .B2(new_n201), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n305), .A2(G159), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n384), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT75), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT73), .ZN(new_n403));
  OR3_X1    g0203(.A1(new_n387), .A2(KEYINPUT73), .A3(G33), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(new_n214), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n222), .B1(new_n405), .B2(KEYINPUT7), .ZN(new_n406));
  INV_X1    g0206(.A(new_n385), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(new_n403), .A3(new_n214), .A4(new_n404), .ZN(new_n408));
  AOI211_X1 g0208(.A(new_n401), .B(new_n402), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(KEYINPUT7), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(G68), .A3(new_n408), .ZN(new_n411));
  INV_X1    g0211(.A(new_n402), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT75), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n400), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n260), .A2(G232), .A3(new_n262), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n264), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G226), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G223), .B2(G1698), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n404), .B2(new_n403), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n259), .A2(new_n224), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n251), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n365), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(G190), .B2(new_n423), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n348), .A2(new_n298), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n297), .B1(new_n337), .B2(new_n348), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n414), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n416), .A2(new_n422), .A3(new_n330), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n264), .A2(new_n415), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n387), .A2(KEYINPUT73), .A3(G33), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n267), .B2(KEYINPUT73), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n434), .A2(new_n419), .B1(new_n259), .B2(new_n224), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n432), .B1(new_n251), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n431), .B(KEYINPUT76), .C1(new_n436), .C2(G169), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT76), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n438), .A3(new_n330), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n414), .A2(new_n427), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT18), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT77), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n414), .A2(new_n427), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n437), .A2(new_n439), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT18), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n440), .A2(KEYINPUT77), .A3(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n430), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n383), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n206), .A2(new_n326), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n210), .A2(G1698), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n403), .B2(new_n404), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G294), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT86), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT86), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n458), .C1(new_n434), .C2(new_n456), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n462), .A3(new_n251), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n261), .B(G45), .C1(new_n252), .C2(KEYINPUT5), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT79), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G41), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n468), .A2(KEYINPUT79), .A3(new_n261), .A4(G45), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n466), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n260), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT87), .B1(new_n472), .B2(new_n211), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n464), .A2(new_n465), .B1(KEYINPUT5), .B2(new_n252), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(G274), .A3(new_n260), .A4(new_n469), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n251), .B1(new_n474), .B2(new_n469), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT87), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(G264), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n463), .A2(new_n473), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n284), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(G179), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n289), .A2(G107), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n482), .B(KEYINPUT25), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n261), .A2(G33), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n297), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n229), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n487));
  AND4_X1   g0287(.A1(new_n214), .A2(new_n267), .A3(new_n487), .A4(G87), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n403), .A2(new_n404), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(new_n214), .A3(G87), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(KEYINPUT22), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n214), .B2(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n229), .A2(KEYINPUT23), .A3(G20), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n493), .A2(new_n494), .B1(new_n496), .B2(new_n214), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT24), .B1(new_n491), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT24), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  AOI21_X1  g0301(.A(G20), .B1(new_n403), .B2(new_n404), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(G87), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n500), .B(new_n497), .C1(new_n503), .C2(new_n488), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n486), .B1(new_n505), .B2(new_n309), .ZN(new_n506));
  OR3_X1    g0306(.A1(new_n481), .A2(new_n506), .A3(KEYINPUT88), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n384), .B1(new_n499), .B2(new_n504), .ZN(new_n508));
  OAI221_X1 g0308(.A(new_n480), .B1(G179), .B2(new_n479), .C1(new_n508), .C2(new_n486), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n479), .A2(new_n365), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n477), .B1(new_n476), .B2(G264), .ZN(new_n512));
  AND4_X1   g0312(.A1(new_n477), .A2(new_n471), .A3(G264), .A4(new_n260), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(new_n369), .A3(new_n475), .A4(new_n463), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n506), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n507), .A2(new_n510), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n471), .A2(G257), .A3(new_n260), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n475), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n386), .A2(new_n388), .A3(G250), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n326), .A2(G244), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n403), .B2(new_n404), .ZN(new_n525));
  AND2_X1   g0325(.A1(KEYINPUT4), .A2(G244), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n386), .A2(new_n388), .A3(new_n526), .A4(new_n326), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n527), .A2(KEYINPUT78), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(KEYINPUT78), .ZN(new_n529));
  OAI221_X1 g0329(.A(new_n523), .B1(new_n525), .B2(KEYINPUT4), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n520), .B1(new_n530), .B2(new_n251), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G190), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n229), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G97), .A2(G107), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n229), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n539), .A2(new_n214), .B1(new_n227), .B2(new_n334), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n407), .B1(G20), .B2(new_n267), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n389), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n229), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n309), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n289), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n485), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(G97), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n532), .B(new_n548), .C1(new_n365), .C2(new_n531), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n547), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n523), .B1(new_n525), .B2(KEYINPUT4), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT78), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n527), .B(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n251), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n519), .A2(new_n475), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n554), .A2(G179), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n284), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n549), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n214), .B1(new_n270), .B2(new_n560), .ZN(new_n561));
  AND4_X1   g0361(.A1(KEYINPUT80), .A2(new_n224), .A3(new_n534), .A4(new_n229), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G87), .A2(G97), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT80), .B1(new_n563), .B2(new_n229), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n489), .A2(new_n214), .A3(G68), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n560), .B1(new_n307), .B2(new_n534), .ZN(new_n569));
  OAI211_X1 g0369(.A(KEYINPUT81), .B(new_n561), .C1(new_n562), .C2(new_n564), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n309), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n335), .A2(new_n337), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n546), .A2(G87), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n223), .A2(new_n326), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n228), .A2(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n403), .B2(new_n404), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n251), .B1(new_n579), .B2(new_n496), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n261), .A2(G45), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n581), .A2(G274), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n206), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n260), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n369), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n584), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n495), .B1(new_n434), .B2(new_n578), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(new_n251), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n588), .B2(G200), .ZN(new_n589));
  INV_X1    g0389(.A(new_n335), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n546), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n572), .A2(new_n573), .A3(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n580), .A2(new_n330), .A3(new_n584), .ZN(new_n593));
  AOI21_X1  g0393(.A(G169), .B1(new_n580), .B2(new_n584), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n575), .A2(new_n589), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT82), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n595), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n571), .A2(new_n309), .B1(new_n337), .B2(new_n335), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n589), .A2(new_n599), .A3(new_n574), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT82), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n559), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n211), .A2(G1698), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(G257), .B2(G1698), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n404), .B2(new_n403), .ZN(new_n606));
  INV_X1    g0406(.A(G303), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n267), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n251), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n471), .A2(G270), .A3(new_n260), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n475), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT83), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n609), .A2(new_n613), .A3(new_n610), .A4(new_n475), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n289), .A2(G116), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n615), .B(KEYINPUT84), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n297), .A2(G116), .A3(new_n484), .ZN(new_n618));
  AOI21_X1  g0418(.A(G20), .B1(new_n259), .B2(G97), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n619), .A2(new_n522), .B1(G20), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n309), .A2(new_n621), .A3(KEYINPUT20), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT20), .B1(new_n309), .B2(new_n621), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n617), .B(new_n618), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n612), .A2(G169), .A3(new_n614), .A4(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n611), .A2(new_n330), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n625), .ZN(new_n630));
  INV_X1    g0430(.A(new_n624), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n616), .B1(new_n631), .B2(new_n622), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n284), .B1(new_n632), .B2(new_n618), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(KEYINPUT21), .A3(new_n612), .A4(new_n614), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n628), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n612), .A2(new_n614), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G200), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n625), .B1(new_n636), .B2(G190), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n603), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n453), .A2(new_n518), .A3(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n363), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n428), .B(KEYINPUT17), .ZN(new_n644));
  INV_X1    g0444(.A(new_n318), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n341), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n315), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n447), .A2(new_n441), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT90), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n381), .B1(new_n380), .B2(new_n371), .ZN(new_n651));
  AOI211_X1 g0451(.A(KEYINPUT10), .B(new_n370), .C1(new_n378), .C2(new_n379), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n377), .A2(KEYINPUT90), .A3(new_n382), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n643), .B1(new_n649), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n598), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n517), .A2(new_n596), .A3(new_n558), .A4(new_n549), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n509), .A2(new_n628), .A3(new_n630), .A4(new_n634), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n558), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n598), .A2(KEYINPUT82), .A3(new_n600), .ZN(new_n662));
  OAI211_X1 g0462(.A(KEYINPUT26), .B(new_n661), .C1(new_n662), .C2(new_n601), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n556), .B2(new_n557), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n554), .A2(G179), .A3(new_n555), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n667), .B(KEYINPUT89), .C1(new_n531), .C2(new_n284), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n550), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n598), .A2(new_n600), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n660), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n656), .B1(new_n453), .B2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n261), .A2(new_n214), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n625), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n640), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n635), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n681), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n506), .A2(new_n688), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n518), .A2(new_n689), .B1(new_n509), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n507), .A2(new_n510), .A3(new_n517), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n635), .A2(new_n688), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n481), .A2(new_n506), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n692), .A2(new_n694), .B1(new_n695), .B2(new_n688), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT91), .ZN(G399));
  OR3_X1    g0498(.A1(new_n209), .A2(KEYINPUT92), .A3(G41), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT92), .B1(new_n209), .B2(G41), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n562), .A2(new_n564), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n620), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(new_n704), .A3(G1), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n216), .B2(new_n701), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n641), .A2(new_n518), .A3(new_n681), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n531), .A2(G179), .A3(new_n588), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n479), .A3(new_n637), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n531), .A2(new_n629), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n514), .A2(new_n463), .A3(new_n588), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n514), .A2(new_n463), .A3(new_n588), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(KEYINPUT30), .A3(new_n629), .A4(new_n531), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n710), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT31), .B1(new_n717), .B2(new_n681), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n708), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n681), .B1(new_n660), .B2(new_n672), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n669), .A2(new_n664), .A3(new_n670), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT93), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT93), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n661), .B1(new_n662), .B2(new_n601), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n728), .B1(new_n729), .B2(new_n664), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n727), .B1(new_n730), .B2(new_n726), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n507), .A2(new_n510), .A3(new_n684), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n657), .B1(new_n732), .B2(new_n658), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n681), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n723), .B1(new_n725), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n707), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(new_n701), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n214), .A2(G13), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n261), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n685), .A2(G330), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n687), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT94), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n742), .B(KEYINPUT95), .Z(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n213), .B1(G20), .B2(new_n284), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n214), .A2(new_n330), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n369), .A2(new_n365), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT97), .Z(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n214), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n369), .A3(G200), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT96), .Z(new_n757));
  AOI22_X1  g0557(.A1(new_n754), .A2(G326), .B1(G283), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n750), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(new_n365), .A3(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT33), .B(G317), .Z(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n755), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(G329), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n751), .A2(new_n755), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n607), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n759), .A2(new_n369), .A3(G200), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(G322), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n750), .A2(new_n764), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n389), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n369), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n214), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n774), .B1(G294), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n758), .A2(new_n767), .A3(new_n771), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n765), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT32), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n389), .B(new_n783), .C1(G58), .C2(new_n770), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G97), .A2(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n752), .A2(new_n202), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n227), .A2(new_n772), .B1(new_n768), .B2(new_n224), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(G68), .C2(new_n760), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n757), .A2(G107), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n784), .A2(new_n785), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n749), .B1(new_n779), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n267), .A2(new_n208), .ZN(new_n792));
  INV_X1    g0592(.A(G355), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n792), .A2(new_n793), .B1(G116), .B2(new_n208), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n489), .A2(new_n209), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n253), .B2(new_n217), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n246), .A2(new_n253), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n748), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n747), .A2(new_n791), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n802), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n685), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n745), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT98), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NOR2_X1   g0611(.A1(new_n748), .A2(new_n800), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n747), .B1(new_n227), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n768), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n267), .B1(new_n814), .B2(G107), .ZN(new_n815));
  INV_X1    g0615(.A(new_n770), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n773), .B2(new_n765), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n757), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n224), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(G97), .C2(new_n777), .ZN(new_n821));
  INV_X1    g0621(.A(new_n752), .ZN(new_n822));
  INV_X1    g0622(.A(new_n772), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G303), .A2(new_n822), .B1(new_n823), .B2(G116), .ZN(new_n824));
  INV_X1    g0624(.A(G283), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n761), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT99), .Z(new_n827));
  AOI22_X1  g0627(.A1(new_n770), .A2(G143), .B1(new_n822), .B2(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n829), .B2(new_n761), .C1(new_n780), .C2(new_n772), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT34), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n819), .A2(new_n222), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n776), .A2(new_n346), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n768), .A2(new_n202), .B1(new_n765), .B2(new_n834), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n832), .A2(new_n434), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n821), .A2(new_n827), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n341), .A2(new_n681), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n340), .A2(new_n681), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n366), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n838), .B1(new_n840), .B2(new_n341), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n813), .B1(new_n749), .B2(new_n837), .C1(new_n841), .C2(new_n801), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT100), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n724), .B2(new_n841), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n663), .A2(new_n671), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n695), .A2(new_n635), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n517), .A2(new_n596), .A3(new_n549), .A4(new_n558), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n598), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n688), .B(new_n841), .C1(new_n845), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(KEYINPUT100), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n844), .A2(new_n850), .B1(new_n724), .B2(new_n841), .ZN(new_n851));
  INV_X1    g0651(.A(new_n723), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n742), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n852), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n842), .B1(new_n854), .B2(new_n855), .ZN(G384));
  INV_X1    g0656(.A(new_n539), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n857), .A2(KEYINPUT35), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(KEYINPUT35), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(G116), .A3(new_n215), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  OAI211_X1 g0661(.A(new_n217), .B(G77), .C1(new_n346), .C2(new_n222), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n202), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n261), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n411), .A2(new_n397), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n384), .B1(new_n867), .B2(new_n399), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n409), .A2(new_n413), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n427), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n679), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n428), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n871), .A2(new_n445), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n414), .A2(new_n425), .A3(new_n427), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n440), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  AOI211_X1 g0679(.A(KEYINPUT101), .B(new_n679), .C1(new_n414), .C2(new_n427), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n444), .B2(new_n872), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n878), .B(new_n879), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n451), .B2(new_n873), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n446), .B1(new_n441), .B2(new_n442), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n644), .B1(new_n887), .B2(new_n449), .ZN(new_n888));
  INV_X1    g0688(.A(new_n873), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n886), .B1(new_n876), .B2(new_n883), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n885), .A2(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n692), .A2(new_n640), .A3(new_n603), .A4(new_n688), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n718), .A2(new_n719), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n302), .A2(new_n304), .A3(new_n313), .A4(new_n312), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n681), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n322), .B2(new_n288), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n318), .A2(new_n897), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n278), .A2(new_n279), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n286), .A2(new_n285), .B1(new_n900), .B2(G179), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n282), .B1(new_n280), .B2(KEYINPUT14), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n285), .A2(KEYINPUT72), .A3(new_n286), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n899), .B1(new_n904), .B2(new_n896), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n841), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n895), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n866), .B1(new_n892), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n882), .A2(new_n880), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n444), .A2(new_n445), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n879), .A3(new_n428), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(KEYINPUT103), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n878), .B1(new_n880), .B2(new_n882), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT103), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n882), .A2(new_n880), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n917), .B1(new_n918), .B2(new_n912), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n914), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n648), .A2(new_n644), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n918), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n923), .A2(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n907), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n909), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT105), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n453), .A2(new_n721), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n722), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n849), .A2(KEYINPUT100), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n673), .A2(new_n843), .A3(new_n688), .A4(new_n841), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n838), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n898), .A2(new_n905), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n933), .A2(new_n892), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n648), .A2(new_n872), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT102), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n838), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n844), .B2(new_n850), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n890), .A2(new_n891), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n888), .A2(new_n889), .B1(new_n883), .B2(new_n876), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n940), .B1(new_n941), .B2(KEYINPUT38), .ZN(new_n942));
  INV_X1    g0742(.A(new_n934), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT102), .ZN(new_n945));
  INV_X1    g0745(.A(new_n936), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n923), .A2(new_n886), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n948), .A2(KEYINPUT104), .A3(new_n949), .A4(new_n940), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT104), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n940), .A2(new_n949), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT38), .B1(new_n920), .B2(new_n922), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n942), .A2(KEYINPUT39), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n315), .A2(new_n688), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n937), .A2(new_n947), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n735), .A2(new_n452), .A3(new_n725), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n656), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n960), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n930), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n261), .B2(new_n739), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n930), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n865), .B1(new_n965), .B2(new_n966), .ZN(G367));
  OAI22_X1  g0767(.A1(new_n829), .A2(new_n816), .B1(new_n761), .B2(new_n780), .ZN(new_n968));
  INV_X1    g0768(.A(new_n756), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n389), .B(new_n968), .C1(G77), .C2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n776), .A2(new_n222), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n754), .A2(G143), .ZN(new_n973));
  INV_X1    g0773(.A(G137), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n772), .A2(new_n202), .B1(new_n765), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G58), .B2(new_n814), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n814), .A2(G116), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT46), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT111), .Z(new_n981));
  AOI22_X1  g0781(.A1(new_n978), .A2(new_n979), .B1(new_n760), .B2(G294), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT112), .Z(new_n984));
  AOI22_X1  g0784(.A1(new_n754), .A2(G311), .B1(G303), .B2(new_n770), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(KEYINPUT110), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(KEYINPUT110), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G283), .A2(new_n823), .B1(new_n766), .B2(G317), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n534), .B2(new_n756), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n489), .B(new_n989), .C1(G107), .C2(new_n777), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n977), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT113), .Z(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT47), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n748), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n596), .B1(new_n575), .B2(new_n688), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n598), .A2(new_n575), .A3(new_n688), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n802), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n803), .B1(new_n208), .B2(new_n335), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n242), .B2(new_n795), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n747), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n996), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n669), .A2(new_n688), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n549), .B(new_n558), .C1(new_n548), .C2(new_n688), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n510), .B2(new_n507), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n688), .B1(new_n1008), .B2(new_n661), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n692), .A2(new_n1006), .A3(new_n694), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT42), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT107), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1010), .A2(KEYINPUT42), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(KEYINPUT107), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n997), .A2(new_n998), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT106), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT43), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1017), .A2(KEYINPUT43), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1022), .A3(new_n1020), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n691), .A2(new_n1007), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1021), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n701), .B(KEYINPUT41), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n690), .A2(KEYINPUT109), .A3(new_n694), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n692), .A2(new_n694), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT109), .B1(new_n690), .B2(new_n694), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(new_n687), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n736), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n696), .A2(new_n1006), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1038), .A2(KEYINPUT44), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(KEYINPUT44), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(KEYINPUT108), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT108), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n696), .A2(new_n1006), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT45), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n696), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1039), .A2(new_n1043), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n687), .A3(new_n690), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1042), .A2(new_n1048), .A3(new_n691), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1037), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1030), .B1(new_n1052), .B2(new_n736), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1053), .A2(new_n741), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1003), .B1(new_n1029), .B2(new_n1054), .ZN(G387));
  OR2_X1    g0855(.A1(new_n690), .A2(new_n807), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n704), .A2(new_n792), .B1(G107), .B2(new_n208), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n796), .B1(new_n238), .B2(G45), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n703), .A2(KEYINPUT114), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n703), .A2(KEYINPUT114), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n333), .A2(G50), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT50), .ZN(new_n1062));
  AOI21_X1  g0862(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1057), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n746), .B1(new_n1065), .B2(new_n804), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n770), .A2(G317), .B1(G303), .B2(new_n823), .ZN(new_n1067));
  XOR2_X1   g0867(.A(KEYINPUT116), .B(G322), .Z(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(new_n773), .B2(new_n761), .C1(new_n753), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n776), .A2(new_n825), .B1(new_n768), .B2(new_n817), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(KEYINPUT49), .A3(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n969), .A2(G116), .B1(new_n766), .B2(G326), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n434), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT49), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G68), .A2(new_n823), .B1(new_n814), .B2(G77), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n777), .A2(new_n590), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n489), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n822), .A2(G159), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT115), .B(G150), .Z(new_n1082));
  OAI221_X1 g0882(.A(new_n1081), .B1(new_n765), .B2(new_n1082), .C1(new_n816), .C2(new_n202), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n348), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n760), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n534), .B2(new_n819), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1076), .A2(new_n1077), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1066), .B1(new_n1087), .B2(new_n748), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1035), .A2(new_n741), .B1(new_n1056), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1036), .A2(new_n738), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1035), .A2(new_n736), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(G393));
  INV_X1    g0892(.A(KEYINPUT117), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1050), .A2(new_n1093), .A3(new_n1051), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1093), .B2(new_n1050), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n738), .B(new_n1052), .C1(new_n1095), .C2(new_n1037), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1007), .A2(new_n802), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n803), .B1(new_n534), .B2(new_n208), .C1(new_n796), .C2(new_n249), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n746), .A2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n770), .A2(G311), .B1(new_n822), .B2(G317), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT52), .Z(new_n1101));
  OAI22_X1  g0901(.A1(new_n1068), .A2(new_n765), .B1(new_n768), .B2(new_n825), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G303), .B2(new_n760), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n389), .B1(new_n772), .B2(new_n817), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G116), .B2(new_n777), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n789), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n768), .A2(new_n222), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n761), .A2(new_n202), .B1(new_n772), .B2(new_n333), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(G143), .C2(new_n766), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n820), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n777), .A2(G77), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1109), .A2(new_n489), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n770), .A2(G159), .B1(new_n822), .B2(G150), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT51), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1106), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1099), .B1(new_n1115), .B2(new_n748), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1095), .A2(new_n741), .B1(new_n1097), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1096), .A2(new_n1117), .ZN(G390));
  AOI21_X1  g0918(.A(new_n910), .B1(new_n644), .B2(new_n648), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n883), .A2(new_n917), .B1(new_n915), .B2(KEYINPUT37), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n914), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n940), .B1(new_n1121), .B2(KEYINPUT38), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n840), .A2(new_n341), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n838), .B1(new_n734), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n934), .B(KEYINPUT118), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n957), .B(new_n1122), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n958), .B1(new_n939), .B2(new_n943), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n956), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n895), .A2(G330), .A3(new_n841), .A4(new_n943), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1129), .B(new_n1126), .C1(new_n1127), .C2(new_n956), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n961), .B(new_n656), .C1(new_n852), .C2(new_n453), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n943), .B1(new_n723), .B2(new_n841), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n939), .B1(new_n1135), .B2(new_n1130), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n895), .A2(KEYINPUT119), .A3(G330), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n841), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT119), .B1(new_n895), .B2(G330), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1125), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1134), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n701), .B1(new_n1133), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1131), .A2(new_n1143), .A3(new_n1132), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n747), .B1(new_n348), .B2(new_n812), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT120), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(KEYINPUT120), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n766), .A2(G125), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n816), .B2(new_n834), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n389), .B(new_n1152), .C1(G137), .C2(new_n760), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n777), .A2(G159), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1082), .A2(new_n768), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n772), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n756), .A2(new_n202), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(G128), .C2(new_n822), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n832), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n229), .A2(new_n761), .B1(new_n816), .B2(new_n620), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G283), .B2(new_n822), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n772), .A2(new_n534), .B1(new_n765), .B2(new_n817), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n267), .B(new_n1165), .C1(G87), .C2(new_n814), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1162), .A2(new_n1164), .A3(new_n1111), .A4(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n749), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1150), .A2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1149), .B(new_n1169), .C1(new_n956), .C2(new_n801), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1133), .B2(new_n740), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1147), .A2(new_n1171), .ZN(G378));
  INV_X1    g0972(.A(KEYINPUT123), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1134), .ZN(new_n1174));
  OAI21_X1  g0974(.A(G330), .B1(new_n924), .B2(new_n925), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n906), .B1(new_n893), .B2(new_n894), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT40), .B1(new_n942), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n653), .A2(new_n654), .A3(new_n363), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n354), .A2(new_n679), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n653), .A2(new_n654), .A3(new_n363), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1175), .A2(new_n1177), .A3(new_n1188), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1184), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n866), .B(new_n906), .C1(new_n893), .C2(new_n894), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n722), .B1(new_n1122), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1192), .B1(new_n1194), .B2(new_n909), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT122), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1188), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT122), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1194), .A2(new_n909), .A3(new_n1192), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n960), .A2(new_n1196), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1202), .A2(new_n937), .A3(new_n959), .A4(new_n947), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1174), .A2(new_n1146), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1173), .B1(new_n1204), .B2(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1146), .A2(new_n1174), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(KEYINPUT123), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1146), .B2(new_n1174), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n960), .A2(new_n1199), .A3(new_n1197), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1203), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n701), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1205), .A2(new_n1210), .A3(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n761), .A2(new_n834), .B1(new_n768), .B2(new_n1157), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n770), .A2(G128), .B1(new_n822), .B2(G125), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n974), .B2(new_n772), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(G150), .C2(new_n777), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n259), .B(new_n252), .C1(new_n756), .C2(new_n780), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G124), .B2(new_n766), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n756), .A2(new_n346), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G77), .B2(new_n814), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n825), .B2(new_n765), .C1(new_n229), .C2(new_n816), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n434), .A2(new_n252), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G116), .A2(new_n822), .B1(new_n823), .B2(new_n590), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n534), .B2(new_n761), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1228), .A2(new_n971), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(KEYINPUT58), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(KEYINPUT58), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1229), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n748), .B1(new_n1225), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n812), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n742), .B1(G50), .B2(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT121), .Z(new_n1240));
  NAND2_X1  g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1192), .B2(new_n800), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1207), .B2(new_n741), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1215), .A2(new_n1243), .ZN(G375));
  AND2_X1   g1044(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT124), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n740), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1125), .A2(new_n800), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n746), .B1(G68), .B2(new_n1238), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n816), .A2(new_n974), .B1(new_n780), .B2(new_n768), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1226), .B(new_n1250), .C1(G128), .C2(new_n766), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n489), .C1(new_n202), .C2(new_n776), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n823), .A2(G150), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n834), .B2(new_n752), .C1(new_n761), .C2(new_n1157), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G294), .A2(new_n822), .B1(new_n823), .B2(G107), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n620), .B2(new_n761), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT125), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n757), .A2(G77), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n267), .B1(new_n766), .B2(G303), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n770), .A2(G283), .B1(G97), .B2(new_n814), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1258), .A2(new_n1079), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1252), .A2(new_n1254), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1249), .B1(new_n1262), .B2(new_n748), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1248), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1246), .B1(new_n1245), .B2(new_n740), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1247), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1245), .A2(new_n1134), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1030), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1144), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(G381));
  OR3_X1    g1071(.A1(G396), .A2(G384), .A3(G393), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(G387), .A2(G381), .A3(G390), .A4(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1147), .A2(new_n1171), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1215), .A4(new_n1243), .ZN(G407));
  NAND2_X1  g1075(.A1(new_n680), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G375), .C2(new_n1278), .ZN(G409));
  NAND3_X1  g1079(.A1(new_n1215), .A2(G378), .A3(new_n1243), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1242), .B1(new_n1213), .B2(new_n741), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1208), .B2(new_n1030), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1274), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1276), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1268), .B1(new_n1286), .B2(new_n1143), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1245), .A2(KEYINPUT60), .A3(new_n1134), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1287), .A2(new_n738), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G384), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n1266), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n738), .A3(new_n1288), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G384), .B1(new_n1267), .B2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G2897), .B(new_n1277), .C1(new_n1291), .C2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1290), .B1(new_n1289), .B2(new_n1266), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1267), .A2(G384), .A3(new_n1292), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1277), .A2(G2897), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT63), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1285), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1003), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1054), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1028), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1025), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1305), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(G390), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(G387), .A2(new_n1096), .A3(new_n1117), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n810), .B(G393), .ZN(new_n1313));
  AND4_X1   g1113(.A1(KEYINPUT126), .A2(new_n1311), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1310), .B2(G390), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n1316), .A2(new_n1313), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1277), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(KEYINPUT63), .A3(new_n1302), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1300), .A2(new_n1304), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1319), .A2(new_n1302), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1319), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(KEYINPUT62), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1319), .B2(new_n1302), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1323), .A2(new_n1326), .A3(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1321), .B1(new_n1330), .B2(new_n1318), .ZN(G405));
  OR2_X1    g1131(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1274), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1280), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1302), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1303), .A3(new_n1280), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1332), .B(new_n1337), .ZN(G402));
endmodule


