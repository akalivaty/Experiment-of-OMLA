//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n941, new_n942;
  INV_X1    g000(.A(G113gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G120gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT71), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  INV_X1    g005(.A(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G127gat), .A2(G134gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT1), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211));
  AND2_X1   g010(.A1(G127gat), .A2(G134gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G127gat), .A2(G134gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(KEYINPUT70), .A3(new_n209), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217));
  INV_X1    g016(.A(new_n203), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n202), .A2(G120gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n205), .A2(new_n210), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  INV_X1    g021(.A(G155gat), .ZN(new_n223));
  INV_X1    g022(.A(G162gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT77), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(G141gat), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G141gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n229), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n227), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G155gat), .B2(G162gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT76), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n237), .A2(new_n226), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n235), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n235), .A2(new_n241), .A3(KEYINPUT78), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n241), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n205), .A2(new_n210), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n216), .A2(new_n220), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT79), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n221), .B1(new_n249), .B2(new_n250), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(KEYINPUT79), .A3(new_n253), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n245), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G225gat), .A2(G233gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT80), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n256), .A2(new_n252), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(new_n243), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT5), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT81), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n243), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n264), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT81), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT5), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n262), .A2(new_n265), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n243), .B(KEYINPUT4), .ZN(new_n275));
  AND4_X1   g074(.A1(KEYINPUT79), .A2(new_n251), .A3(new_n253), .A4(new_n256), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT79), .B1(new_n260), .B2(new_n253), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n265), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT82), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G85gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G57gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  NAND2_X1  g083(.A1(new_n273), .A2(new_n269), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT82), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n289));
  INV_X1    g088(.A(new_n284), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n278), .A2(new_n285), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n259), .A2(new_n261), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n293), .A2(new_n268), .A3(new_n265), .A4(new_n275), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n290), .B1(new_n295), .B2(new_n286), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(KEYINPUT6), .B(new_n290), .C1(new_n295), .C2(new_n286), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G8gat), .B(G36gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G197gat), .B(G204gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT22), .ZN(new_n305));
  NAND2_X1  g104(.A1(G211gat), .A2(G218gat), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  INV_X1    g106(.A(G218gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n306), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n304), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  OR3_X1    g115(.A1(new_n316), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT27), .B1(new_n316), .B2(KEYINPUT69), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G169gat), .ZN(new_n322));
  INV_X1    g121(.A(G176gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(KEYINPUT26), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n315), .B(new_n321), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT27), .B(G183gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n318), .B1(new_n330), .B2(new_n319), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n315), .A2(KEYINPUT24), .ZN(new_n337));
  NOR2_X1   g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT67), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT64), .ZN(new_n342));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n343), .B2(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n345), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n341), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT67), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n348), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n340), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n328), .B1(KEYINPUT23), .B2(new_n343), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT66), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT64), .B1(new_n324), .B2(new_n345), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n343), .A2(new_n342), .A3(KEYINPUT23), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT65), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n339), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n346), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT65), .A3(new_n351), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  AOI221_X4 g161(.A(new_n334), .B1(new_n350), .B2(new_n353), .C1(new_n362), .C2(new_n341), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n341), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n350), .A2(new_n353), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT68), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n333), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G226gat), .ZN(new_n368));
  INV_X1    g167(.A(G233gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(KEYINPUT29), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n362), .A2(new_n341), .B1(new_n350), .B2(new_n353), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(new_n332), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n360), .A2(KEYINPUT65), .A3(new_n351), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT65), .B1(new_n360), .B2(new_n351), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n376), .A2(new_n377), .A3(new_n339), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n365), .B1(new_n378), .B2(KEYINPUT25), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(KEYINPUT74), .A3(new_n333), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n370), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n314), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n370), .B(new_n333), .C1(new_n363), .C2(new_n366), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n375), .A2(new_n380), .A3(new_n371), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n314), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n303), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT30), .ZN(new_n389));
  INV_X1    g188(.A(new_n314), .ZN(new_n390));
  INV_X1    g189(.A(new_n371), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n379), .A2(new_n334), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n374), .A2(KEYINPUT68), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n394), .B2(new_n333), .ZN(new_n395));
  INV_X1    g194(.A(new_n370), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n375), .B2(new_n380), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n386), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n303), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n371), .A2(new_n367), .B1(new_n381), .B2(new_n370), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n386), .B(new_n302), .C1(new_n402), .C2(new_n314), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT75), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n398), .A2(KEYINPUT75), .A3(new_n386), .A4(new_n302), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n389), .A2(new_n401), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n299), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT83), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n299), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT84), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n310), .B(KEYINPUT85), .Z(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n313), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n242), .B1(new_n419), .B2(new_n246), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n314), .B1(new_n251), .B2(new_n418), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G22gat), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT86), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n246), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n390), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n252), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n421), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n427), .A2(G228gat), .A3(G233gat), .A4(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n423), .B1(new_n422), .B2(new_n429), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n413), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT87), .A3(new_n430), .ZN(new_n435));
  XNOR2_X1  g234(.A(G78gat), .B(G106gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT31), .B(G50gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n413), .B(new_n440), .C1(new_n431), .C2(new_n432), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n221), .B(new_n333), .C1(new_n363), .C2(new_n366), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT72), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n394), .A2(KEYINPUT72), .A3(new_n221), .A4(new_n333), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n367), .A2(new_n256), .ZN(new_n447));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT34), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT73), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n449), .A2(KEYINPUT34), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(KEYINPUT73), .A3(KEYINPUT34), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT32), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n457));
  INV_X1    g256(.A(new_n448), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT33), .B1(new_n457), .B2(new_n458), .ZN(new_n460));
  XNOR2_X1  g259(.A(G15gat), .B(G43gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n461), .B(new_n462), .Z(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n459), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  AOI221_X4 g264(.A(new_n456), .B1(KEYINPUT33), .B2(new_n463), .C1(new_n457), .C2(new_n458), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n455), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n457), .A2(new_n458), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n459), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n449), .A2(KEYINPUT73), .A3(KEYINPUT34), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT73), .B1(new_n449), .B2(KEYINPUT34), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(new_n464), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n472), .A2(new_n475), .A3(new_n476), .A4(new_n453), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n442), .A2(new_n467), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT35), .B1(new_n412), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n389), .A2(new_n401), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT35), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n405), .A2(new_n406), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n299), .A2(KEYINPUT93), .ZN(new_n484));
  INV_X1    g283(.A(new_n298), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(KEYINPUT93), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n467), .A2(new_n477), .A3(KEYINPUT94), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT94), .B1(new_n467), .B2(new_n477), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n442), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n479), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT92), .B(KEYINPUT38), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT37), .B1(new_n398), .B2(new_n386), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT91), .B1(new_n402), .B2(new_n390), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(new_n314), .C1(new_n395), .C2(new_n397), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AOI211_X1 g298(.A(new_n493), .B(new_n494), .C1(new_n499), .C2(KEYINPUT37), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n302), .A2(new_n493), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n500), .A2(new_n303), .B1(new_n399), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n486), .B1(new_n299), .B2(KEYINPUT93), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n398), .A2(KEYINPUT37), .A3(new_n386), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n493), .B1(new_n504), .B2(new_n494), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n439), .A2(new_n441), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n270), .A2(new_n264), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT89), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(new_n264), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT39), .B(new_n509), .C1(new_n512), .C2(new_n508), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n264), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n284), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n516), .A2(KEYINPUT90), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n516), .B2(KEYINPUT90), .ZN(new_n519));
  INV_X1    g318(.A(new_n296), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n407), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n507), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n465), .A2(new_n455), .A3(new_n466), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n476), .A2(new_n472), .B1(new_n475), .B2(new_n453), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n467), .A2(new_n477), .A3(KEYINPUT36), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n411), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n410), .B1(new_n299), .B2(new_n407), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n507), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n524), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n492), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(G1gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT100), .ZN(new_n540));
  INV_X1    g339(.A(G8gat), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT16), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(G1gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT99), .ZN(new_n547));
  NAND2_X1  g346(.A1(KEYINPUT100), .A2(G8gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT99), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n542), .A2(new_n547), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(G8gat), .B1(new_n546), .B2(new_n539), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G71gat), .B(G78gat), .ZN(new_n554));
  AND2_X1   g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  INV_X1    g354(.A(G57gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G64gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT101), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n556), .A2(G64gat), .ZN(new_n559));
  OAI221_X1 g358(.A(new_n554), .B1(KEYINPUT9), .B2(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n556), .A2(G64gat), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n557), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n563), .A2(new_n554), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n553), .B1(KEYINPUT21), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(new_n316), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  OR3_X1    g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G211gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n571), .B1(new_n569), .B2(new_n570), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n575), .B1(new_n572), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n537), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n572), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n574), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n536), .A3(new_n577), .ZN(new_n583));
  NAND3_X1  g382(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(KEYINPUT102), .B(KEYINPUT7), .Z(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n585), .A2(new_n588), .B1(KEYINPUT8), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n587), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n590), .B(new_n591), .C1(new_n588), .C2(new_n585), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G43gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT15), .B1(new_n595), .B2(G50gat), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n595), .B2(G50gat), .ZN(new_n597));
  OR3_X1    g396(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT97), .B(G29gat), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G36gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n595), .A2(G50gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT98), .B(G50gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n603), .B1(new_n604), .B2(new_n595), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n600), .B(new_n602), .C1(KEYINPUT15), .C2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n599), .B1(new_n598), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n597), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(KEYINPUT17), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n584), .B(new_n613), .C1(new_n615), .C2(new_n594), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G134gat), .B(G162gat), .Z(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n580), .A2(new_n583), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n535), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n612), .A2(new_n553), .ZN(new_n625));
  INV_X1    g424(.A(new_n553), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n614), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT18), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n612), .B(new_n553), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n628), .B(KEYINPUT13), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G169gat), .B(G197gat), .Z(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT95), .B(KEYINPUT11), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G113gat), .B(G141gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n630), .A2(new_n642), .A3(new_n633), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  INV_X1    g445(.A(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT104), .B(G176gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n592), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n565), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n594), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n594), .A2(KEYINPUT10), .A3(new_n565), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT105), .Z(new_n661));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n654), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n650), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n660), .ZN(new_n665));
  INV_X1    g464(.A(new_n650), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n665), .B(new_n666), .C1(new_n660), .C2(new_n654), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n645), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n624), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n299), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g472(.A1(new_n670), .A2(new_n522), .ZN(new_n674));
  NAND2_X1  g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n543), .A2(new_n541), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT106), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n674), .A2(new_n541), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n680), .B(new_n681), .C1(new_n678), .C2(new_n677), .ZN(G1325gat));
  NOR2_X1   g481(.A1(new_n489), .A2(new_n490), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(G15gat), .B1(new_n670), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT107), .ZN(new_n686));
  INV_X1    g485(.A(new_n530), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(G15gat), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n670), .B2(new_n688), .ZN(G1326gat));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n507), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n423), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n622), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n535), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n695), .A2(KEYINPUT109), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n695), .B2(KEYINPUT109), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n580), .A2(new_n583), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n669), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n601), .B1(new_n702), .B2(new_n299), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n535), .A2(new_n694), .A3(new_n701), .ZN(new_n704));
  INV_X1    g503(.A(new_n601), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n671), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(G1328gat));
  OAI21_X1  g507(.A(G36gat), .B1(new_n702), .B2(new_n407), .ZN(new_n709));
  INV_X1    g508(.A(G36gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n704), .A2(new_n710), .A3(new_n522), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT46), .Z(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(G1329gat));
  NOR3_X1   g512(.A1(new_n702), .A2(new_n595), .A3(new_n530), .ZN(new_n714));
  AOI21_X1  g513(.A(G43gat), .B1(new_n704), .B2(new_n684), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g516(.A(new_n604), .B1(new_n702), .B2(new_n442), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n442), .A2(new_n604), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT110), .Z(new_n720));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT48), .Z(G1331gat));
  AND3_X1   g522(.A1(new_n624), .A2(new_n645), .A3(new_n668), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n671), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n522), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n728), .B(new_n729), .Z(G1333gat));
  AOI21_X1  g529(.A(G71gat), .B1(new_n724), .B2(new_n684), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n687), .A2(G71gat), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g533(.A1(new_n724), .A2(new_n507), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  INV_X1    g535(.A(new_n700), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n644), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n697), .A2(new_n668), .A3(new_n698), .A4(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n299), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  AOI22_X1  g540(.A1(new_n412), .A2(new_n507), .B1(new_n528), .B2(new_n529), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n524), .A2(new_n742), .B1(new_n479), .B2(new_n491), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(new_n622), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n535), .A2(KEYINPUT111), .A3(new_n694), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n738), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT51), .A4(new_n738), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n750), .A2(new_n749), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n668), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n671), .A2(new_n586), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n740), .B1(new_n753), .B2(new_n754), .ZN(G1336gat));
  NAND3_X1  g554(.A1(new_n522), .A2(new_n668), .A3(new_n587), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT113), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n751), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G92gat), .B1(new_n739), .B2(new_n407), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n748), .A2(new_n750), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n757), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(KEYINPUT52), .ZN(new_n766));
  AOI211_X1 g565(.A(KEYINPUT114), .B(new_n760), .C1(new_n759), .C2(new_n764), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n761), .B1(new_n766), .B2(new_n767), .ZN(G1337gat));
  XOR2_X1   g567(.A(KEYINPUT115), .B(G99gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n739), .B2(new_n530), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n683), .A2(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n753), .B2(new_n771), .ZN(G1338gat));
  INV_X1    g571(.A(new_n668), .ZN(new_n773));
  OR3_X1    g572(.A1(new_n442), .A2(G106gat), .A3(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT116), .Z(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n751), .A2(new_n752), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT117), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  OAI21_X1  g578(.A(G106gat), .B1(new_n739), .B2(new_n442), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n751), .A2(new_n752), .A3(new_n781), .A4(new_n776), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n780), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n775), .B1(new_n748), .B2(new_n750), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT53), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT118), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n783), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1339gat));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n666), .B1(new_n662), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n659), .A2(new_n661), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(KEYINPUT54), .A3(new_n665), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n794), .B1(new_n793), .B2(new_n796), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n644), .B(new_n667), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n627), .A2(new_n628), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n631), .A2(new_n632), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n639), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n643), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n668), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n694), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n667), .B(new_n694), .C1(new_n798), .C2(new_n799), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n804), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n700), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n623), .A2(new_n811), .A3(new_n645), .A4(new_n773), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n580), .A2(new_n583), .A3(new_n773), .A4(new_n622), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT119), .B1(new_n813), .B2(new_n644), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n522), .A2(new_n299), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n478), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n202), .A3(new_n644), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n683), .A2(new_n507), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G113gat), .B1(new_n823), .B2(new_n645), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(G1340gat));
  NOR2_X1   g624(.A1(new_n773), .A2(new_n204), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G120gat), .B1(new_n823), .B2(new_n773), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1341gat));
  AOI21_X1  g628(.A(G127gat), .B1(new_n820), .B2(new_n737), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n823), .A2(new_n206), .A3(new_n700), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(G1342gat));
  NAND3_X1  g631(.A1(new_n820), .A2(new_n207), .A3(new_n694), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT56), .Z(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n823), .B2(new_n622), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT120), .Z(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n507), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n530), .A2(new_n817), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(G141gat), .A3(new_n645), .ZN(new_n842));
  INV_X1    g641(.A(new_n839), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n816), .B2(new_n507), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  AOI211_X1 g644(.A(new_n845), .B(new_n442), .C1(new_n810), .C2(new_n815), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT121), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n849), .B(new_n843), .C1(new_n844), .C2(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n644), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n842), .B1(new_n852), .B2(G141gat), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n847), .A2(new_n645), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT58), .B(new_n842), .C1(new_n856), .C2(G141gat), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n855), .A2(new_n857), .ZN(G1344gat));
  INV_X1    g657(.A(KEYINPUT125), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n813), .A2(new_n644), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n808), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n799), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n797), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(KEYINPUT123), .A3(new_n667), .A4(new_n694), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n865), .A3(new_n805), .ZN(new_n866));
  INV_X1    g665(.A(new_n807), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n860), .B1(new_n868), .B2(new_n700), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n845), .B1(new_n869), .B2(new_n442), .ZN(new_n870));
  INV_X1    g669(.A(new_n846), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n773), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n839), .B(KEYINPUT122), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G148gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(KEYINPUT124), .A3(KEYINPUT59), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n229), .B1(new_n872), .B2(new_n873), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT59), .B1(new_n851), .B2(new_n668), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n230), .A2(new_n231), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n876), .A2(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n841), .A2(new_n883), .A3(new_n773), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n859), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n851), .A2(new_n668), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n879), .A3(new_n883), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT124), .B1(new_n875), .B2(KEYINPUT59), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n878), .A2(new_n877), .A3(new_n879), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n885), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(KEYINPUT125), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n886), .A2(new_n893), .ZN(G1345gat));
  AOI21_X1  g693(.A(G155gat), .B1(new_n840), .B2(new_n737), .ZN(new_n895));
  INV_X1    g694(.A(new_n851), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n700), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g697(.A(G162gat), .B1(new_n840), .B2(new_n694), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n896), .A2(new_n622), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(G162gat), .ZN(G1347gat));
  INV_X1    g700(.A(new_n816), .ZN(new_n902));
  INV_X1    g701(.A(new_n822), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n671), .A2(new_n407), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT126), .Z(new_n905));
  NOR3_X1   g704(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G169gat), .B1(new_n907), .B2(new_n645), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n816), .A2(new_n819), .A3(new_n904), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n322), .A3(new_n644), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1348gat));
  AOI21_X1  g710(.A(G176gat), .B1(new_n909), .B2(new_n668), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n773), .A2(new_n323), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n906), .B2(new_n913), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n907), .B2(new_n700), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n909), .A2(new_n330), .A3(new_n737), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n907), .B2(new_n622), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(KEYINPUT127), .B2(KEYINPUT61), .ZN(new_n920));
  NOR2_X1   g719(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n909), .A2(new_n319), .A3(new_n694), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1351gat));
  NAND4_X1  g723(.A1(new_n816), .A2(new_n507), .A3(new_n530), .A4(new_n904), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(G197gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(new_n644), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n905), .A2(new_n687), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n870), .B2(new_n871), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(new_n644), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(new_n927), .ZN(G1352gat));
  NOR3_X1   g731(.A1(new_n925), .A2(G204gat), .A3(new_n773), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n773), .B(new_n929), .C1(new_n870), .C2(new_n871), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n647), .B2(new_n935), .ZN(G1353gat));
  AOI21_X1  g735(.A(new_n307), .B1(new_n930), .B2(new_n737), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT63), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n926), .A2(new_n307), .A3(new_n737), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1354gat));
  AOI21_X1  g739(.A(G218gat), .B1(new_n926), .B2(new_n694), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n622), .A2(new_n308), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n930), .B2(new_n942), .ZN(G1355gat));
endmodule


