//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT64), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G125), .B(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n188), .B2(new_n193), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT75), .B(G237), .Z(new_n196));
  INV_X1    g010(.A(G953), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(G214), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT75), .B(G237), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G953), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(G143), .A3(G214), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT18), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n203), .ZN(new_n208));
  AOI21_X1  g022(.A(G143), .B1(new_n202), .B2(G214), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI221_X1 g024(.A(new_n195), .B1(new_n204), .B2(new_n207), .C1(new_n210), .C2(new_n205), .ZN(new_n211));
  XNOR2_X1  g025(.A(G113), .B(G122), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n200), .A2(new_n206), .A3(new_n203), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n206), .B1(new_n200), .B2(new_n203), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT17), .ZN(new_n217));
  INV_X1    g031(.A(G125), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n218), .A2(KEYINPUT16), .A3(G140), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT78), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n193), .B2(KEYINPUT16), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n188), .ZN(new_n224));
  OAI211_X1 g038(.A(G146), .B(new_n220), .C1(new_n222), .C2(new_n219), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n224), .B(new_n225), .C1(new_n210), .C2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n211), .B(new_n214), .C1(new_n217), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT91), .B1(new_n215), .B2(new_n216), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT91), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n200), .A2(new_n206), .A3(new_n203), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n210), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT19), .ZN(new_n233));
  OR2_X1    g047(.A1(new_n193), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n193), .A2(new_n233), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(new_n192), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT92), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n193), .B(KEYINPUT19), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT92), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(new_n192), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n237), .A2(new_n240), .A3(new_n225), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n229), .A2(new_n232), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n214), .B1(new_n242), .B2(new_n211), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n228), .B1(new_n243), .B2(KEYINPUT93), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT93), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n245), .B(new_n214), .C1(new_n242), .C2(new_n211), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n187), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT20), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(new_n187), .C1(new_n244), .C2(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n211), .B1(new_n217), .B2(new_n227), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(new_n214), .ZN(new_n253));
  OAI21_X1  g067(.A(G475), .B1(new_n253), .B2(G902), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(G234), .A2(G237), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(G952), .A3(new_n197), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT76), .B(G902), .Z(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(G953), .A3(new_n256), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT21), .B(G898), .Z(new_n260));
  OAI21_X1  g074(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G128), .B(G143), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT96), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n263), .A2(KEYINPUT96), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  INV_X1    g081(.A(G116), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n268), .A2(G122), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n269), .B2(KEYINPUT14), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(G122), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n270), .B(new_n272), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n265), .A2(new_n266), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT9), .B(G234), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G217), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n277), .A2(new_n278), .A3(G953), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT13), .ZN(new_n280));
  INV_X1    g094(.A(G128), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(G143), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n282), .A2(KEYINPUT94), .B1(new_n281), .B2(G143), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(KEYINPUT94), .B2(new_n282), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT95), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT95), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n283), .B(new_n286), .C1(KEYINPUT94), .C2(new_n282), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n199), .A2(G128), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n285), .B(new_n287), .C1(new_n280), .C2(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n289), .A2(G134), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n272), .A2(new_n267), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n269), .A2(new_n271), .A3(G107), .ZN(new_n292));
  INV_X1    g106(.A(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n262), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n275), .B(new_n279), .C1(new_n290), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n279), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n289), .B2(G134), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(new_n274), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT97), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n258), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n298), .A2(new_n274), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT97), .A3(new_n279), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G478), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n306), .A2(KEYINPUT15), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n305), .B(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n255), .A2(new_n261), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G122), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT8), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n267), .A2(KEYINPUT83), .A3(G104), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n267), .A2(G104), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G101), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n319), .A2(new_n267), .A3(KEYINPUT83), .A4(G104), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n315), .A2(new_n317), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n213), .A2(G107), .ZN(new_n322));
  OAI21_X1  g136(.A(G101), .B1(new_n322), .B2(new_n316), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT2), .B(G113), .Z(new_n326));
  AND2_X1   g140(.A1(KEYINPUT73), .A2(G119), .ZN(new_n327));
  NOR2_X1   g141(.A1(KEYINPUT73), .A2(G119), .ZN(new_n328));
  OAI21_X1  g142(.A(G116), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n268), .A2(G119), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(KEYINPUT5), .A3(new_n330), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(G113), .C1(KEYINPUT5), .C2(new_n329), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n325), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n332), .ZN(new_n335));
  OAI21_X1  g149(.A(G113), .B1(new_n329), .B2(KEYINPUT5), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(new_n324), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n313), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n315), .A2(new_n320), .A3(new_n317), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G101), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT4), .A3(new_n321), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n329), .A2(new_n330), .ZN(new_n343));
  INV_X1    g157(.A(new_n326), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n331), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n347), .A3(G101), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n325), .A2(new_n333), .A3(new_n331), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n312), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n199), .B1(new_n189), .B2(new_n191), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT1), .ZN(new_n354));
  OAI21_X1  g168(.A(G128), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n188), .A2(G143), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n192), .B2(G143), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT71), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT71), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n354), .B1(new_n192), .B2(G143), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n360), .B(new_n357), .C1(new_n361), .C2(new_n281), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n188), .A2(G143), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n192), .B2(G143), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n354), .A3(G128), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n359), .A2(new_n218), .A3(new_n362), .A4(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n362), .A2(new_n365), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(KEYINPUT88), .A3(new_n218), .A4(new_n359), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT65), .ZN(new_n371));
  INV_X1    g185(.A(new_n363), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT64), .B(G146), .ZN(new_n373));
  OAI211_X1 g187(.A(G128), .B(new_n372), .C1(new_n373), .C2(new_n199), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT0), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n364), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g192(.A(KEYINPUT0), .B(G128), .Z(new_n379));
  NAND2_X1  g193(.A1(new_n357), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n368), .A2(new_n370), .B1(G125), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n197), .A2(G224), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n383), .A2(KEYINPUT7), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n352), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n368), .A2(new_n370), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n387), .A3(G125), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n376), .A2(new_n377), .B1(new_n357), .B2(new_n379), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT87), .B1(new_n389), .B2(new_n218), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n386), .A2(new_n391), .A3(new_n384), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n311), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(KEYINPUT90), .B(new_n311), .C1(new_n385), .C2(new_n392), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n386), .A2(new_n391), .A3(new_n383), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n383), .B1(new_n386), .B2(new_n391), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n351), .A2(KEYINPUT6), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n312), .B1(new_n349), .B2(new_n350), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI211_X1 g217(.A(KEYINPUT6), .B(new_n312), .C1(new_n349), .C2(new_n350), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT89), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n405), .B(new_n408), .C1(new_n398), .C2(new_n399), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G210), .B1(G237), .B2(G902), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n397), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n397), .B2(new_n410), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n310), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G469), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n281), .B1(new_n356), .B2(KEYINPUT1), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n416), .B1(new_n364), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n417), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n419), .B(KEYINPUT84), .C1(new_n353), .C2(new_n363), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n420), .A3(new_n365), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n325), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n422), .B1(new_n423), .B2(new_n325), .ZN(new_n424));
  INV_X1    g238(.A(G137), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT66), .B1(new_n425), .B2(G134), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT66), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n293), .A3(G137), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT11), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n293), .B2(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(KEYINPUT11), .A3(G134), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n429), .A2(new_n206), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n431), .A2(new_n432), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT67), .A3(new_n206), .A4(new_n429), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n429), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G131), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n424), .A2(KEYINPUT12), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n424), .A2(KEYINPUT86), .A3(KEYINPUT12), .A4(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n424), .A2(new_n441), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n197), .A2(G227), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT82), .ZN(new_n451));
  XOR2_X1   g265(.A(G110), .B(G140), .Z(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n423), .A2(KEYINPUT10), .A3(new_n325), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT10), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n422), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n342), .A2(new_n348), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n389), .ZN(new_n458));
  INV_X1    g272(.A(new_n441), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n454), .A2(new_n456), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT85), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n455), .A2(new_n422), .B1(new_n457), .B2(new_n389), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n462), .A2(new_n463), .A3(new_n459), .A4(new_n454), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n449), .A2(new_n453), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n454), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n441), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n453), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n415), .B(new_n302), .C1(new_n466), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n465), .A2(new_n453), .A3(new_n468), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n449), .A2(new_n465), .ZN(new_n472));
  OAI211_X1 g286(.A(G469), .B(new_n471), .C1(new_n472), .C2(new_n453), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n415), .A2(new_n311), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G221), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n276), .B2(new_n311), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n309), .A2(new_n414), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n425), .A2(KEYINPUT69), .A3(G134), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT69), .B1(new_n425), .B2(G134), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n483), .B(new_n484), .C1(new_n293), .C2(G137), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n435), .A2(new_n437), .B1(G131), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n362), .A2(new_n365), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n360), .B1(new_n355), .B2(new_n357), .ZN(new_n489));
  OAI22_X1  g303(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(G131), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n438), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n482), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n438), .A2(new_n491), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n486), .A2(new_n487), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(KEYINPUT72), .A3(new_n423), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n441), .A2(new_n389), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n441), .A2(new_n389), .A3(KEYINPUT68), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n493), .A2(new_n497), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n423), .A2(new_n486), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT74), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n423), .A2(KEYINPUT74), .A3(new_n486), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n507), .A2(KEYINPUT30), .A3(new_n508), .A4(new_n498), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n346), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n508), .A3(new_n498), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n511), .A2(new_n346), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n202), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n318), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n514), .B(new_n515), .Z(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT31), .ZN(new_n518));
  INV_X1    g332(.A(new_n516), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n502), .A2(new_n346), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n520), .B1(new_n512), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n505), .A2(new_n331), .A3(new_n345), .A4(new_n498), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n520), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n519), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n510), .A2(new_n527), .A3(new_n512), .A4(new_n516), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n518), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(G472), .A2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT32), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n510), .A2(new_n512), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n519), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n511), .A2(new_n346), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n346), .B2(new_n502), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n524), .B(new_n516), .C1(new_n537), .C2(new_n520), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n511), .B(new_n346), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n525), .B1(new_n541), .B2(KEYINPUT28), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n519), .A2(new_n539), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n258), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G472), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n529), .A2(KEYINPUT32), .A3(new_n530), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n533), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n278), .B1(new_n302), .B2(G234), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT79), .ZN(new_n551));
  INV_X1    g365(.A(G110), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n281), .A2(KEYINPUT23), .A3(G119), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n327), .A2(new_n328), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(new_n281), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT23), .B1(new_n554), .B2(new_n281), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g371(.A1(KEYINPUT73), .A2(G119), .ZN(new_n558));
  NAND2_X1  g372(.A1(KEYINPUT73), .A2(G119), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n281), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT77), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT77), .B1(new_n281), .B2(G119), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n562), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G110), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n552), .A2(new_n557), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n224), .B2(new_n225), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n552), .A2(new_n557), .B1(new_n564), .B2(new_n565), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n225), .A2(new_n194), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n551), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n224), .A2(new_n225), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n555), .A2(new_n556), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G110), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n572), .B(new_n574), .C1(new_n565), .C2(new_n564), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(G110), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n564), .A2(new_n565), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n194), .B(new_n225), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n578), .A3(KEYINPUT79), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT22), .B(G137), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n197), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n571), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n575), .A2(new_n578), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n551), .A3(new_n582), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n258), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n550), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n258), .B(new_n588), .C1(new_n584), .C2(new_n586), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n549), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n584), .A2(new_n586), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n549), .A2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(KEYINPUT81), .Z(new_n597));
  NOR2_X1   g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n481), .A2(new_n548), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  OAI211_X1 g414(.A(new_n261), .B(new_n310), .C1(new_n412), .C2(new_n413), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n251), .A2(new_n254), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n301), .A2(new_n603), .A3(new_n304), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n296), .A2(new_n299), .A3(KEYINPUT33), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(G478), .A3(new_n302), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n305), .A2(new_n306), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT98), .B1(new_n601), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n310), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n397), .A2(new_n410), .ZN(new_n612));
  INV_X1    g426(.A(new_n411), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n397), .A2(new_n410), .A3(new_n411), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n609), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n261), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n529), .A2(new_n302), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G472), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(new_n531), .ZN(new_n623));
  INV_X1    g437(.A(new_n598), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n480), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n620), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  OR2_X1    g442(.A1(new_n602), .A2(new_n308), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n601), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n623), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n583), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n585), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n595), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n592), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n635), .B1(new_n623), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n641), .A2(new_n635), .A3(new_n622), .A4(new_n531), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n481), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT37), .B(G110), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  NOR2_X1   g461(.A1(new_n414), .A2(new_n480), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n257), .B(KEYINPUT102), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(G900), .B2(new_n259), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n629), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n548), .A2(new_n648), .A3(new_n641), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n529), .A2(KEYINPUT32), .A3(new_n530), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT32), .B1(new_n529), .B2(new_n530), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n519), .B1(new_n510), .B2(new_n512), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n311), .B1(new_n541), .B2(new_n516), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n657), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n533), .A2(new_n657), .A3(new_n547), .A4(new_n663), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n614), .A2(new_n615), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  INV_X1    g483(.A(new_n639), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n308), .B1(new_n251), .B2(new_n254), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n669), .A2(new_n310), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n656), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n480), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n651), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT40), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n667), .A2(new_n672), .A3(new_n656), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n199), .ZN(G45));
  NOR2_X1   g496(.A1(new_n609), .A2(new_n652), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n548), .A2(new_n648), .A3(new_n641), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  AOI21_X1  g499(.A(new_n624), .B1(new_n660), .B2(new_n546), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n466), .A2(new_n469), .ZN(new_n687));
  OAI21_X1  g501(.A(G469), .B1(new_n687), .B2(new_n258), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n479), .A3(new_n470), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n686), .A2(new_n620), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n548), .A2(new_n630), .A3(new_n598), .A4(new_n690), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  INV_X1    g511(.A(new_n309), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n414), .A2(new_n689), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n548), .A2(new_n698), .A3(new_n641), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  OAI211_X1 g515(.A(new_n671), .B(new_n310), .C1(new_n412), .C2(new_n413), .ZN(new_n702));
  INV_X1    g516(.A(new_n261), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT107), .B(G472), .Z(new_n705));
  OAI211_X1 g519(.A(new_n518), .B(new_n528), .C1(new_n516), .C2(new_n542), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n621), .A2(new_n705), .B1(new_n530), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n704), .A2(new_n598), .A3(new_n690), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  NAND4_X1  g523(.A1(new_n699), .A2(new_n707), .A3(new_n639), .A4(new_n683), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT108), .B(G125), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G27));
  NAND3_X1  g526(.A1(new_n614), .A2(new_n310), .A3(new_n615), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n480), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n548), .A2(new_n598), .A3(new_n683), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT42), .B1(new_n715), .B2(KEYINPUT109), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT110), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n716), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G131), .ZN(G33));
  AND4_X1   g540(.A1(new_n548), .A2(new_n598), .A3(new_n653), .A4(new_n714), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n293), .ZN(G36));
  NAND2_X1  g542(.A1(new_n255), .A2(new_n608), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT43), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n623), .A3(new_n670), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n729), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n639), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n733), .B1(new_n736), .B2(new_n623), .ZN(new_n737));
  INV_X1    g551(.A(new_n713), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n471), .B1(new_n472), .B2(new_n453), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n415), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n740), .B2(new_n739), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(KEYINPUT46), .A3(new_n475), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n470), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT46), .B1(new_n742), .B2(new_n475), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n479), .B(new_n676), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n732), .A2(new_n737), .A3(new_n738), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G137), .ZN(G39));
  OAI21_X1  g563(.A(new_n479), .B1(new_n744), .B2(new_n745), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT47), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n752), .B(new_n479), .C1(new_n744), .C2(new_n745), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n683), .A2(new_n624), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n548), .A2(new_n754), .A3(new_n713), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  NAND3_X1  g571(.A1(new_n533), .A2(new_n547), .A3(new_n663), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT103), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n665), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n624), .A2(new_n729), .A3(new_n611), .A4(new_n478), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n688), .A2(new_n470), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT49), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(KEYINPUT49), .ZN(new_n765));
  OR4_X1    g579(.A1(new_n760), .A2(new_n764), .A3(new_n669), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n255), .A2(new_n308), .A3(new_n651), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT112), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n255), .A2(new_n770), .A3(new_n308), .A4(new_n651), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n548), .A2(new_n641), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n707), .A2(new_n639), .A3(new_n683), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n727), .B1(new_n774), .B2(new_n714), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n719), .B2(new_n724), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n601), .B1(new_n609), .B2(new_n629), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n623), .A3(new_n625), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n599), .B(new_n779), .C1(new_n642), .C2(new_n644), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n708), .A2(new_n700), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n694), .A2(new_n695), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n694), .A2(new_n695), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n691), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n780), .B1(new_n784), .B2(KEYINPUT111), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n696), .A2(new_n786), .A3(new_n691), .A4(new_n781), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n777), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n639), .A2(new_n652), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n674), .A2(new_n616), .A3(new_n671), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n664), .B2(new_n666), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n760), .A2(KEYINPUT113), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n654), .A2(new_n684), .A3(new_n710), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n760), .B2(new_n791), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n793), .B(new_n790), .C1(new_n759), .C2(new_n665), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT52), .B(new_n798), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n788), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(KEYINPUT114), .A3(new_n802), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n799), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n805), .B1(new_n813), .B2(new_n788), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(KEYINPUT115), .B(new_n805), .C1(new_n813), .C2(new_n788), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n767), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n707), .A2(new_n598), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n649), .A2(new_n819), .A3(new_n735), .A4(new_n690), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n669), .A2(new_n310), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(KEYINPUT50), .A3(new_n821), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n730), .A2(new_n650), .A3(new_n689), .A4(new_n713), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n639), .A3(new_n707), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n738), .A2(new_n690), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n760), .A2(new_n257), .A3(new_n624), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n255), .A3(new_n607), .A4(new_n606), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n762), .A2(new_n479), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n751), .A2(new_n753), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(KEYINPUT117), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(KEYINPUT117), .B2(new_n835), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n649), .A2(new_n819), .A3(new_n738), .A4(new_n735), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT51), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n830), .A2(new_n617), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n820), .A2(new_n616), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(G952), .A3(new_n197), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n827), .A2(new_n686), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n835), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n838), .B1(new_n848), .B2(new_n834), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT51), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n841), .B(new_n847), .C1(new_n832), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n840), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n805), .B1(new_n788), .B2(new_n804), .ZN(new_n855));
  INV_X1    g669(.A(new_n780), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n775), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n722), .A2(new_n716), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n784), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT116), .B1(new_n784), .B2(new_n858), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n810), .A3(new_n812), .A4(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n855), .A2(new_n767), .A3(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n840), .A2(new_n851), .A3(KEYINPUT118), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n818), .A2(new_n854), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(G952), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n766), .B1(new_n866), .B2(new_n867), .ZN(G75));
  NAND2_X1  g682(.A1(new_n855), .A2(new_n863), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n258), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n411), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n400), .B(new_n405), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT55), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(KEYINPUT119), .B2(new_n874), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n871), .A2(KEYINPUT56), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n871), .B2(KEYINPUT56), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n197), .A2(G952), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(G51));
  XNOR2_X1  g694(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n474), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n767), .B1(new_n855), .B2(new_n863), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n882), .B1(new_n864), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n687), .B(KEYINPUT121), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n870), .A2(new_n742), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n878), .B1(new_n886), .B2(new_n887), .ZN(G54));
  INV_X1    g702(.A(new_n870), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n244), .A2(new_n246), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(KEYINPUT58), .A2(G475), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n891), .B1(new_n889), .B2(new_n892), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(new_n878), .ZN(G60));
  NAND2_X1  g709(.A1(new_n604), .A2(new_n605), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT122), .ZN(new_n897));
  NAND2_X1  g711(.A1(G478), .A2(G902), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT59), .Z(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n864), .B2(new_n883), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(KEYINPUT123), .B(new_n900), .C1(new_n864), .C2(new_n883), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n879), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n899), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n818), .B2(new_n864), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n905), .B1(new_n907), .B2(new_n897), .ZN(G63));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n909));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT60), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n855), .B2(new_n863), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n637), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n879), .B1(new_n912), .B2(new_n594), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n909), .B(KEYINPUT61), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n913), .B(new_n879), .C1(new_n594), .C2(new_n912), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT61), .B1(new_n918), .B2(new_n909), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n919), .ZN(G66));
  AOI21_X1  g734(.A(new_n197), .B1(new_n260), .B2(G224), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n785), .A2(new_n787), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n197), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n406), .B1(G898), .B2(new_n197), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n923), .B(new_n924), .Z(G69));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n713), .B1(new_n609), .B2(new_n629), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n686), .A2(new_n674), .A3(new_n676), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n748), .A2(new_n756), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n797), .B1(new_n930), .B2(KEYINPUT62), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n679), .B2(new_n680), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n933), .B(new_n931), .C1(new_n679), .C2(new_n680), .ZN(new_n936));
  AOI21_X1  g750(.A(G953), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n504), .A2(new_n509), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n238), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n926), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(G900), .B2(G953), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n624), .B(new_n702), .C1(new_n660), .C2(new_n546), .ZN(new_n943));
  AOI211_X1 g757(.A(new_n727), .B(new_n797), .C1(new_n747), .C2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n725), .A2(new_n944), .A3(new_n748), .A4(new_n756), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(G953), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n937), .A2(new_n926), .A3(new_n940), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT127), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n197), .B1(G227), .B2(G900), .ZN(new_n950));
  OR3_X1    g764(.A1(new_n937), .A2(new_n926), .A3(new_n940), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n951), .A2(new_n952), .A3(new_n946), .A4(new_n941), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n950), .B1(new_n949), .B2(new_n953), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(G72));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n935), .A2(new_n936), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n922), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n661), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n958), .B1(new_n945), .B2(new_n922), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n534), .A2(new_n516), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n878), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n816), .A2(new_n817), .ZN(new_n966));
  INV_X1    g780(.A(new_n958), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n535), .B2(new_n517), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n965), .B1(new_n966), .B2(new_n968), .ZN(G57));
endmodule


