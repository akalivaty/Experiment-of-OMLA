//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(G237), .A2(G953), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(G143), .A3(G214), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT18), .A3(G131), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT18), .A2(G131), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n194), .A2(new_n196), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n198), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n211));
  AND4_X1   g025(.A1(G143), .A2(new_n190), .A3(new_n191), .A4(G214), .ZN(new_n212));
  AOI21_X1  g026(.A(G143), .B1(new_n195), .B2(G214), .ZN(new_n213));
  OAI21_X1  g027(.A(G131), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n197), .A2(KEYINPUT84), .A3(G131), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n199), .A3(G125), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n203), .B2(new_n219), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n205), .ZN(new_n222));
  OAI211_X1 g036(.A(G146), .B(new_n220), .C1(new_n203), .C2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT85), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT84), .B1(new_n197), .B2(G131), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  AOI211_X1 g041(.A(new_n215), .B(new_n227), .C1(new_n194), .C2(new_n196), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT17), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT85), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n222), .A2(new_n223), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n226), .A2(new_n228), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT86), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n194), .A2(new_n227), .A3(new_n196), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n211), .A4(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n216), .A2(new_n217), .A3(new_n211), .A4(new_n236), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT86), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n189), .B(new_n210), .C1(new_n233), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n225), .A2(new_n232), .A3(new_n237), .A4(new_n239), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n244), .A2(KEYINPUT87), .A3(new_n189), .A4(new_n210), .ZN(new_n245));
  INV_X1    g059(.A(new_n189), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n210), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n243), .A2(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G475), .B1(new_n248), .B2(G902), .ZN(new_n249));
  INV_X1    g063(.A(G902), .ZN(new_n250));
  XOR2_X1   g064(.A(G116), .B(G122), .Z(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G107), .ZN(new_n252));
  XNOR2_X1  g066(.A(G116), .B(G122), .ZN(new_n253));
  INV_X1    g067(.A(G107), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(KEYINPUT13), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(G143), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n258), .B2(KEYINPUT13), .ZN(new_n261));
  OAI21_X1  g075(.A(G134), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n193), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G134), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n256), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT88), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G116), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT14), .A3(G122), .ZN(new_n271));
  OAI211_X1 g085(.A(G107), .B(new_n271), .C1(new_n251), .C2(KEYINPUT14), .ZN(new_n272));
  OAI21_X1  g086(.A(G134), .B1(new_n258), .B2(new_n263), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n266), .A2(new_n273), .B1(new_n254), .B2(new_n253), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n267), .A2(new_n268), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT70), .B(G217), .Z(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT9), .B(G234), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n276), .A2(G953), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n269), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n278), .B1(new_n269), .B2(new_n275), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT89), .B(new_n250), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G478), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT15), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n281), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n279), .ZN(new_n287));
  INV_X1    g101(.A(new_n284), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(KEYINPUT89), .A3(new_n250), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(G234), .A2(G237), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(G952), .A3(new_n191), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(G902), .A3(G953), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT21), .B(G898), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT20), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n243), .A2(new_n245), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n234), .A2(new_n236), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n203), .B(KEYINPUT19), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n301), .B(new_n223), .C1(G146), .C2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n303), .B2(new_n210), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G475), .A2(G902), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n304), .B1(new_n243), .B2(new_n245), .ZN(new_n309));
  INV_X1    g123(.A(new_n307), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n309), .A2(KEYINPUT20), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n249), .B(new_n298), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT90), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n306), .A2(new_n299), .A3(new_n307), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT20), .B1(new_n309), .B2(new_n310), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n249), .A4(new_n298), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n276), .B1(G234), .B2(new_n250), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n257), .B2(G119), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT71), .A3(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n257), .A2(G119), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT24), .B(G110), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(KEYINPUT73), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n324), .A2(new_n326), .B1(G119), .B2(new_n257), .ZN(new_n333));
  INV_X1    g147(.A(new_n330), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT72), .B1(new_n325), .B2(G128), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT23), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n328), .A2(KEYINPUT72), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G110), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n325), .A2(G128), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n337), .A2(new_n339), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n331), .A2(new_n335), .A3(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n223), .A2(new_n206), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n346), .A2(G110), .B1(new_n333), .B2(new_n334), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n224), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT74), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n354), .A3(KEYINPUT75), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n343), .A2(new_n344), .B1(new_n224), .B2(new_n347), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n353), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n352), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n322), .B1(new_n360), .B2(G902), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n357), .A2(new_n353), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n362), .A2(KEYINPUT75), .B1(new_n357), .B2(new_n352), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n363), .A2(KEYINPUT25), .A3(new_n250), .A4(new_n358), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n321), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n320), .A2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n363), .A2(new_n368), .A3(new_n358), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n360), .A2(KEYINPUT76), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G472), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n250), .A3(KEYINPUT67), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(G472), .B2(G902), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT0), .A2(G128), .ZN(new_n380));
  OR2_X1    g194(.A1(KEYINPUT0), .A2(G128), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n193), .A2(G146), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n205), .A2(G143), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT64), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n193), .B2(G146), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n205), .A2(KEYINPUT64), .A3(G143), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n193), .A2(G146), .ZN(new_n388));
  INV_X1    g202(.A(new_n380), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT11), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n265), .B2(G137), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n265), .A2(G137), .ZN(new_n394));
  INV_X1    g208(.A(G137), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT11), .A3(G134), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G131), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n396), .A3(new_n227), .A4(new_n394), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n391), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G116), .B(G119), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT2), .B(G113), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT2), .B(G113), .Z(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n402), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n395), .A2(G134), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n265), .A2(G137), .ZN(new_n411));
  OAI21_X1  g225(.A(G131), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n205), .A2(G143), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT1), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n414), .A2(G128), .B1(new_n413), .B2(new_n388), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n416));
  AND4_X1   g230(.A1(new_n386), .A2(new_n387), .A3(new_n416), .A4(new_n388), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n412), .B(new_n399), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n401), .A2(new_n409), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT28), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n419), .A2(KEYINPUT66), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT66), .B1(new_n419), .B2(new_n420), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n384), .A2(new_n390), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n399), .B2(new_n398), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n399), .A2(new_n412), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n386), .A2(new_n387), .A3(new_n416), .A4(new_n388), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT1), .ZN(new_n428));
  OAI21_X1  g242(.A(G128), .B1(new_n382), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n413), .A2(new_n388), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n426), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n408), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n419), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT65), .B1(new_n434), .B2(KEYINPUT28), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT65), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n436), .B(new_n420), .C1(new_n433), .C2(new_n419), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n423), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n195), .A2(G210), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT27), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT26), .B(G101), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n401), .A2(new_n445), .A3(new_n418), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n401), .B2(new_n418), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n408), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n442), .A3(new_n419), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT31), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n448), .A2(KEYINPUT31), .A3(new_n442), .A4(new_n419), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n379), .B1(new_n444), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT68), .B1(new_n454), .B2(KEYINPUT32), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT68), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n443), .A2(new_n438), .B1(new_n451), .B2(new_n452), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n379), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n434), .A2(KEYINPUT28), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n423), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n442), .A2(KEYINPUT29), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n250), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n442), .B(new_n423), .C1(new_n435), .C2(new_n437), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n448), .A2(new_n419), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT29), .B1(new_n466), .B2(new_n443), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT69), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n465), .A2(KEYINPUT69), .A3(new_n467), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n374), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n458), .A2(new_n457), .A3(new_n379), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n373), .B1(new_n460), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G210), .B1(G237), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G122), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G113), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n402), .B2(KEYINPUT5), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT5), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n325), .A3(G116), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n482), .A2(new_n325), .A3(KEYINPUT79), .A4(G116), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n481), .A2(new_n487), .A3(KEYINPUT80), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT80), .B1(new_n481), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n254), .A3(G104), .ZN(new_n492));
  INV_X1    g306(.A(G101), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n188), .A2(G107), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n188), .A2(G107), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n254), .A2(G104), .ZN(new_n497));
  OAI21_X1  g311(.A(G101), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n407), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n488), .A2(new_n489), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G101), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n504), .A3(G101), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n503), .A2(new_n408), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n479), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n481), .A2(new_n487), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT80), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n407), .A2(new_n495), .A3(new_n498), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n481), .A2(new_n487), .A3(KEYINPUT80), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n503), .A2(new_n408), .A3(new_n505), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n478), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n507), .A2(KEYINPUT6), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n517), .B(new_n479), .C1(new_n500), .C2(new_n506), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n424), .A2(G125), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n431), .A2(new_n427), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n519), .B1(G125), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G224), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(G953), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n521), .B(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n516), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n478), .B(KEYINPUT8), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n510), .A2(new_n407), .A3(new_n512), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n495), .A2(new_n498), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n511), .A2(new_n508), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT81), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n511), .A2(KEYINPUT81), .A3(new_n508), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT7), .B1(new_n522), .B2(G953), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n415), .A2(new_n417), .A3(G125), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n201), .B1(new_n384), .B2(new_n390), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT82), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n521), .A2(KEYINPUT82), .A3(new_n535), .ZN(new_n541));
  OR3_X1    g355(.A1(new_n536), .A2(new_n537), .A3(new_n535), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n540), .A2(new_n515), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n250), .B1(new_n534), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n477), .B1(new_n525), .B2(new_n544), .ZN(new_n545));
  AND4_X1   g359(.A1(new_n515), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n528), .A2(new_n529), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n530), .A2(new_n531), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n533), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n526), .ZN(new_n550));
  AOI21_X1  g364(.A(G902), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n516), .A2(new_n518), .A3(new_n524), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n476), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT83), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(KEYINPUT83), .B(new_n477), .C1(new_n525), .C2(new_n544), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G214), .B1(G237), .B2(G902), .ZN(new_n559));
  OAI21_X1  g373(.A(G221), .B1(new_n277), .B2(G902), .ZN(new_n560));
  XNOR2_X1  g374(.A(G110), .B(G140), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n191), .A2(G227), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n429), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n427), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n495), .A2(new_n498), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n400), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n503), .A2(new_n391), .A3(new_n505), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n569), .B1(new_n431), .B2(new_n427), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n567), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n568), .A2(new_n569), .B1(new_n567), .B2(new_n573), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n571), .B1(new_n577), .B2(new_n572), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n563), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n520), .A2(new_n567), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n529), .B1(new_n427), .B2(new_n565), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n400), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT12), .ZN(new_n583));
  INV_X1    g397(.A(new_n563), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n400), .C1(new_n580), .C2(new_n581), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n583), .A2(new_n575), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n579), .A2(KEYINPUT78), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(G469), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n590), .B(new_n563), .C1(new_n576), .C2(new_n578), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n588), .A2(new_n589), .A3(new_n250), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(G469), .A2(G902), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n583), .A2(new_n575), .A3(new_n586), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT77), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n583), .A2(new_n575), .A3(new_n596), .A4(new_n586), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n563), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n572), .B(new_n574), .C1(KEYINPUT10), .C2(new_n581), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n400), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n584), .A3(new_n575), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n592), .B(new_n593), .C1(new_n589), .C2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n558), .A2(new_n559), .A3(new_n560), .A4(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n319), .A2(new_n475), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  OAI21_X1  g421(.A(new_n249), .B1(new_n308), .B2(new_n311), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n287), .B(KEYINPUT33), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n283), .A2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n287), .A2(new_n250), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT92), .B(G478), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n559), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n545), .B2(new_n553), .ZN(new_n618));
  INV_X1    g432(.A(new_n297), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT91), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n458), .B2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n444), .A2(new_n453), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(KEYINPUT91), .A3(new_n250), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n625), .A3(G472), .ZN(new_n626));
  INV_X1    g440(.A(new_n454), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n603), .A2(new_n372), .A3(new_n560), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT93), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  OAI211_X1 g448(.A(new_n249), .B(new_n290), .C1(new_n308), .C2(new_n311), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n620), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(KEYINPUT36), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n353), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n349), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n357), .A2(new_n640), .A3(new_n353), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n366), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT94), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n361), .A2(new_n364), .ZN(new_n646));
  OAI211_X1 g460(.A(KEYINPUT95), .B(new_n645), .C1(new_n646), .C2(new_n321), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n644), .B(KEYINPUT94), .Z(new_n649));
  OAI21_X1  g463(.A(new_n648), .B1(new_n365), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n651), .A2(new_n626), .A3(new_n627), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n247), .A2(new_n246), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n300), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n250), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n314), .A2(new_n315), .B1(new_n655), .B2(G475), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n317), .B1(new_n656), .B2(new_n298), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n312), .A2(KEYINPUT90), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n605), .B(new_n652), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  XNOR2_X1  g475(.A(KEYINPUT96), .B(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n293), .B1(new_n295), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n635), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n468), .A2(new_n469), .ZN(new_n665));
  INV_X1    g479(.A(new_n464), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n471), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n454), .A2(KEYINPUT32), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n455), .A4(new_n459), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n603), .A2(new_n560), .A3(new_n618), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n664), .A2(new_n670), .A3(new_n651), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XOR2_X1   g487(.A(new_n663), .B(KEYINPUT39), .Z(new_n674));
  NAND3_X1  g488(.A1(new_n603), .A2(new_n560), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT40), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n466), .A2(new_n442), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n434), .A2(new_n442), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(G902), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n374), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n473), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n455), .A3(new_n459), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n647), .A2(new_n650), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n682), .A2(new_n559), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n290), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n656), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n557), .B(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n676), .A2(new_n684), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  AOI21_X1  g504(.A(new_n683), .B1(new_n460), .B2(new_n474), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n609), .A2(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n656), .A2(new_n692), .A3(new_n663), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n691), .A2(new_n671), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND3_X1  g509(.A1(new_n588), .A2(new_n250), .A3(new_n591), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n592), .ZN(new_n698));
  INV_X1    g512(.A(new_n560), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n465), .A2(KEYINPUT69), .A3(new_n467), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT69), .B1(new_n465), .B2(new_n467), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n701), .A2(new_n702), .A3(new_n464), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n669), .B1(new_n703), .B2(new_n374), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n455), .A2(new_n459), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n372), .B(new_n700), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n692), .B1(new_n316), .B2(new_n249), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n619), .A3(new_n618), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT41), .B(G113), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n636), .A2(new_n670), .A3(new_n372), .A4(new_n700), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  AND2_X1   g527(.A1(new_n697), .A2(new_n592), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT98), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n560), .A4(new_n618), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n618), .A2(new_n560), .A3(new_n592), .A4(new_n697), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT98), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n319), .A2(new_n719), .A3(new_n691), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  OAI21_X1  g535(.A(G472), .B1(new_n458), .B2(G902), .ZN(new_n722));
  INV_X1    g536(.A(new_n462), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n453), .B1(new_n442), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n378), .B(KEYINPUT99), .Z(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n372), .A3(new_n726), .A4(new_n619), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n717), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n686), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NAND2_X1  g544(.A1(new_n722), .A2(new_n726), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n650), .B2(new_n647), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n693), .A2(new_n718), .A3(new_n716), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n601), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n601), .A2(new_n735), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n598), .A2(new_n736), .A3(G469), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n592), .A3(new_n593), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n699), .A2(new_n617), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n557), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n670), .A2(new_n372), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  INV_X1    g557(.A(new_n663), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n707), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n608), .A2(new_n615), .A3(new_n744), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n557), .A2(new_n739), .A3(new_n740), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n457), .B1(new_n458), .B2(new_n379), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n669), .B(new_n750), .C1(new_n703), .C2(new_n374), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT101), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n751), .A2(new_n752), .A3(new_n372), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(new_n751), .B2(new_n372), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n746), .B1(new_n755), .B2(KEYINPUT42), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND3_X1  g571(.A1(new_n475), .A2(new_n664), .A3(new_n741), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NAND3_X1  g573(.A1(new_n316), .A2(new_n249), .A3(new_n615), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n762), .B1(new_n760), .B2(new_n761), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT104), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n761), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n683), .B1(new_n627), .B2(new_n626), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n765), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n557), .A2(new_n559), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT102), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n598), .A2(new_n736), .A3(KEYINPUT45), .A4(new_n737), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n598), .A2(new_n601), .ZN(new_n778));
  OAI211_X1 g592(.A(G469), .B(new_n777), .C1(new_n778), .C2(KEYINPUT45), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n593), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n593), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n592), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n560), .ZN(new_n785));
  INV_X1    g599(.A(new_n674), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n776), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(KEYINPUT102), .A3(new_n560), .A4(new_n674), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n775), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n765), .A2(new_n770), .A3(KEYINPUT44), .A4(new_n771), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n774), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  NOR2_X1   g606(.A1(new_n704), .A2(new_n705), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n775), .A2(new_n372), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n693), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT105), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n693), .A2(new_n793), .A3(KEYINPUT105), .A4(new_n794), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n560), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT47), .B1(new_n784), .B2(new_n560), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  NOR3_X1   g616(.A1(new_n682), .A2(new_n373), .A3(new_n292), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n775), .A2(new_n699), .A3(new_n698), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g619(.A(G952), .B(new_n191), .C1(new_n805), .C2(new_n616), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n731), .A2(new_n373), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n293), .B(new_n807), .C1(new_n763), .C2(new_n764), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n806), .B1(new_n719), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n292), .B1(new_n767), .B2(new_n769), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n804), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n293), .B(new_n804), .C1(new_n763), .C2(new_n764), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n751), .A2(new_n752), .A3(new_n372), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n454), .A2(KEYINPUT32), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n472), .A2(new_n473), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT101), .B1(new_n818), .B2(new_n373), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n813), .A2(new_n815), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n810), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n775), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n811), .A2(new_n807), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n785), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n560), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n698), .A2(new_n560), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n827), .B1(KEYINPUT113), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(KEYINPUT113), .B2(new_n833), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n805), .A2(new_n608), .A3(new_n615), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n700), .A2(new_n617), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n688), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n808), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n811), .A2(KEYINPUT50), .A3(new_n807), .A4(new_n839), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n836), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n813), .A2(new_n815), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n732), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n835), .A2(KEYINPUT51), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n799), .A2(new_n800), .A3(new_n831), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT111), .B1(new_n847), .B2(new_n827), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT111), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n833), .A2(new_n849), .A3(new_n826), .A4(new_n809), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n845), .A2(new_n843), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n825), .A2(new_n846), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT108), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n604), .B1(new_n313), .B2(new_n318), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n555), .A2(new_n556), .A3(new_n619), .A4(new_n559), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n628), .A2(new_n629), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n616), .A2(new_n635), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n856), .A2(new_n475), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n855), .B1(new_n860), .B2(new_n659), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n855), .A2(new_n606), .A3(new_n659), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n313), .A2(new_n318), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n670), .A2(new_n651), .A3(new_n718), .A4(new_n716), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n712), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n729), .B1(new_n706), .B2(new_n708), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n603), .A2(new_n685), .A3(new_n560), .A4(new_n744), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n608), .A2(new_n870), .A3(new_n775), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n749), .A2(new_n732), .B1(new_n691), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n756), .A3(new_n758), .A4(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n608), .A2(new_n290), .A3(new_n618), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n365), .A2(new_n649), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n663), .A2(KEYINPUT109), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT109), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n699), .B1(new_n744), .B2(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n876), .A2(new_n739), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n875), .A2(new_n682), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n694), .A2(new_n733), .A3(new_n881), .A4(new_n672), .ZN(new_n882));
  AND2_X1   g696(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n691), .B(new_n671), .C1(new_n664), .C2(new_n693), .ZN(new_n885));
  NOR2_X1   g699(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n733), .A3(new_n881), .A4(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n874), .B2(new_n889), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n656), .A2(new_n727), .A3(new_n717), .A4(new_n685), .ZN(new_n891));
  INV_X1    g705(.A(new_n706), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n621), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n872), .A3(new_n712), .A4(new_n720), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n742), .A2(new_n745), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n707), .A2(new_n741), .A3(new_n744), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n819), .B2(new_n816), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n895), .B(new_n758), .C1(new_n897), .C2(new_n743), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n606), .A2(new_n659), .A3(new_n862), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT108), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n860), .A2(new_n855), .A3(new_n659), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n882), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n733), .A4(new_n881), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n899), .A2(new_n903), .A3(new_n907), .A4(KEYINPUT53), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT54), .B1(new_n890), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n899), .A2(new_n903), .A3(new_n907), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n899), .A4(new_n903), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n854), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT115), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT115), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n854), .A2(new_n910), .A3(new_n919), .A4(new_n916), .ZN(new_n920));
  OR2_X1    g734(.A1(G952), .A2(G953), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n760), .A2(new_n373), .A3(new_n617), .A4(new_n699), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n682), .B(new_n688), .C1(KEYINPUT49), .C2(new_n698), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n698), .A2(KEYINPUT49), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT107), .Z(new_n928));
  NAND4_X1  g742(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n922), .A2(new_n929), .ZN(G75));
  AOI21_X1  g744(.A(new_n250), .B1(new_n913), .B2(new_n914), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n932), .A3(G210), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n516), .A2(new_n518), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n524), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n932), .B1(new_n931), .B2(G210), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n191), .A2(G952), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT56), .B1(new_n931), .B2(G210), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n940), .A2(new_n944), .ZN(G51));
  AND3_X1   g759(.A1(new_n913), .A2(new_n915), .A3(new_n914), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n593), .B(KEYINPUT57), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n588), .B(new_n591), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n779), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n931), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n941), .B1(new_n950), .B2(new_n952), .ZN(G54));
  AND2_X1   g767(.A1(KEYINPUT58), .A2(G475), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n931), .A2(new_n306), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n306), .B1(new_n931), .B2(new_n954), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n941), .ZN(G60));
  INV_X1    g771(.A(KEYINPUT117), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n910), .A2(new_n916), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT59), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n609), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n609), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n961), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n946), .B2(new_n947), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n942), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n958), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n899), .A2(new_n903), .A3(new_n888), .A4(new_n884), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n912), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n915), .B1(new_n970), .B2(new_n908), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n962), .B1(new_n946), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n964), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(KEYINPUT117), .A3(new_n942), .A4(new_n966), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n968), .A2(new_n974), .ZN(G63));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT60), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n913), .B2(new_n914), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n369), .A2(new_n370), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n642), .A2(new_n643), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT119), .Z(new_n982));
  AOI21_X1  g796(.A(new_n941), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT61), .B1(new_n984), .B2(KEYINPUT118), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT118), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n986), .B(new_n987), .C1(new_n980), .C2(new_n983), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n985), .A2(new_n988), .ZN(G66));
  INV_X1    g803(.A(new_n296), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n191), .B1(new_n990), .B2(G224), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n903), .A2(new_n869), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT120), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n993), .B2(new_n191), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n935), .B1(G898), .B2(new_n191), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT121), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n994), .B(new_n996), .ZN(G69));
  AOI21_X1  g811(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n446), .A2(new_n447), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(new_n302), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n775), .A2(new_n675), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n475), .A2(new_n859), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT122), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n475), .A2(new_n859), .A3(KEYINPUT122), .A4(new_n1003), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n801), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n689), .A2(new_n733), .A3(new_n885), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n885), .A2(new_n733), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(KEYINPUT62), .A3(new_n689), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1009), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n791), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1002), .B1(new_n1016), .B2(new_n191), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT124), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n801), .A2(new_n1013), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n875), .B1(new_n753), .B2(new_n754), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1020), .B1(new_n787), .B2(new_n788), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n898), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1022), .A2(new_n191), .A3(new_n791), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1001), .B1(G900), .B2(G953), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1018), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1017), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1024), .A2(new_n1018), .A3(new_n1025), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n999), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT123), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1017), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(G953), .B1(new_n1015), .B2(new_n791), .ZN(new_n1032));
  OAI21_X1  g846(.A(KEYINPUT123), .B1(new_n1032), .B2(new_n1002), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n998), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(KEYINPUT125), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT125), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1028), .ZN(new_n1039));
  NOR3_X1   g853(.A1(new_n1039), .A2(new_n1017), .A3(new_n1026), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n1037), .B(new_n1038), .C1(new_n1040), .C2(new_n999), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1036), .A2(new_n1041), .ZN(G72));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  NAND3_X1  g858(.A1(new_n1022), .A2(new_n791), .A3(new_n1023), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1044), .B1(new_n993), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1046), .A2(new_n443), .A3(new_n419), .A4(new_n448), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n993), .A2(new_n1016), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1044), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g864(.A(new_n1047), .B(new_n942), .C1(new_n1050), .C2(new_n677), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n466), .A2(new_n443), .ZN(new_n1052));
  XOR2_X1   g866(.A(new_n1052), .B(KEYINPUT126), .Z(new_n1053));
  INV_X1    g867(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1049), .B1(new_n1054), .B2(new_n449), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1055), .B1(new_n890), .B2(new_n909), .ZN(new_n1056));
  XOR2_X1   g870(.A(new_n1056), .B(KEYINPUT127), .Z(new_n1057));
  NOR2_X1   g871(.A1(new_n1051), .A2(new_n1057), .ZN(G57));
endmodule


