//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027;
  XOR2_X1   g000(.A(KEYINPUT71), .B(KEYINPUT2), .Z(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(G148gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G127gat), .ZN(new_n214));
  INV_X1    g013(.A(G127gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G134gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G113gat), .B(G120gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT64), .A2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G120gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G113gat), .ZN(new_n223));
  INV_X1    g022(.A(G113gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G120gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G127gat), .B(G134gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(new_n219), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n208), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(KEYINPUT72), .A2(G148gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(KEYINPUT72), .A2(G148gat), .ZN(new_n234));
  OAI21_X1  g033(.A(G141gat), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI221_X4 g034(.A(new_n230), .B1(new_n232), .B2(new_n210), .C1(new_n235), .C2(new_n204), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n204), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n210), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT73), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n212), .B(new_n229), .C1(new_n236), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT4), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT75), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT72), .B(G148gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n205), .B1(new_n243), .B2(G141gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n238), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n230), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n237), .A2(KEYINPUT73), .A3(new_n238), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n248), .A2(new_n249), .A3(new_n212), .A4(new_n229), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n242), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n212), .B(new_n254), .C1(new_n236), .C2(new_n239), .ZN(new_n255));
  INV_X1    g054(.A(new_n229), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n246), .A2(new_n247), .B1(new_n207), .B2(new_n211), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n255), .B(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n257), .A2(KEYINPUT75), .A3(new_n249), .A4(new_n229), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n251), .A2(new_n252), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  OR3_X1    g060(.A1(new_n257), .A2(KEYINPUT76), .A3(new_n229), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n212), .B1(new_n236), .B2(new_n239), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n256), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(KEYINPUT76), .A3(new_n240), .ZN(new_n265));
  INV_X1    g064(.A(new_n252), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(KEYINPUT5), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G1gat), .B(G29gat), .ZN(new_n269));
  INV_X1    g068(.A(G85gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT0), .B(G57gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n241), .A2(new_n250), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n259), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n268), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n274), .B1(new_n268), .B2(new_n277), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI211_X1 g081(.A(new_n279), .B(new_n274), .C1(new_n268), .C2(new_n277), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT24), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(G183gat), .A3(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G169gat), .ZN(new_n297));
  INV_X1    g096(.A(G176gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n293), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT25), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n291), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n299), .A2(KEYINPUT26), .A3(new_n294), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n294), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(new_n308), .A3(new_n291), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n305), .A2(new_n306), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n299), .B1(new_n289), .B2(new_n292), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n296), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n302), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G226gat), .ZN(new_n317));
  INV_X1    g116(.A(G233gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n319), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT69), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326));
  AND2_X1   g125(.A1(G197gat), .A2(G204gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(G197gat), .A2(G204gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G197gat), .ZN(new_n330));
  INV_X1    g129(.A(G204gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G197gat), .A2(G204gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT68), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G211gat), .B(G218gat), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n325), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n337), .B1(new_n325), .B2(new_n335), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n323), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n329), .A2(new_n334), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n324), .B(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n336), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n335), .A3(new_n337), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(KEYINPUT70), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n321), .A2(new_n322), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n319), .B1(new_n314), .B2(new_n315), .ZN(new_n350));
  AND4_X1   g149(.A1(new_n312), .A2(new_n293), .A3(new_n296), .A4(new_n300), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n312), .B1(new_n311), .B2(new_n296), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n320), .B1(new_n353), .B2(new_n310), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n347), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n349), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n355), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n350), .A2(new_n354), .A3(new_n347), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n349), .A2(new_n355), .A3(KEYINPUT30), .A4(new_n359), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n362), .A2(new_n365), .A3(new_n369), .A4(new_n366), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT80), .B1(new_n284), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT35), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n314), .A2(new_n256), .ZN(new_n374));
  INV_X1    g173(.A(G227gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(new_n318), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n302), .A2(new_n310), .A3(new_n229), .A4(new_n313), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT34), .ZN(new_n380));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT65), .ZN(new_n382));
  XOR2_X1   g181(.A(G15gat), .B(G43gat), .Z(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n377), .B1(new_n374), .B2(new_n378), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(KEYINPUT33), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT32), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n378), .ZN(new_n390));
  AOI221_X4 g189(.A(new_n387), .B1(KEYINPUT33), .B2(new_n384), .C1(new_n390), .C2(new_n376), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n380), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n229), .B1(new_n353), .B2(new_n310), .ZN(new_n393));
  INV_X1    g192(.A(new_n378), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n376), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT32), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n398), .A3(new_n384), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT34), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n379), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n388), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT67), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n392), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n402), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT67), .A3(new_n380), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G22gat), .B(G50gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n346), .A2(new_n340), .B1(new_n255), .B2(new_n315), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n344), .A2(new_n345), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n263), .A2(new_n414), .A3(new_n315), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n412), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n255), .A2(new_n315), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n347), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n263), .A2(new_n253), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n420), .A2(new_n411), .A3(new_n415), .A4(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT77), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n418), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n418), .B2(new_n422), .ZN(new_n426));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT31), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n418), .A2(new_n422), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n430), .B1(new_n432), .B2(new_n424), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n410), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n428), .B1(new_n425), .B2(new_n426), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n430), .A3(new_n424), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n409), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n408), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n371), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n268), .A2(new_n277), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n273), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n279), .A3(new_n278), .ZN(new_n442));
  INV_X1    g241(.A(new_n283), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT80), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n439), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n372), .A2(new_n373), .A3(new_n438), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n367), .B1(new_n442), .B2(new_n443), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n392), .A2(new_n403), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n406), .A2(KEYINPUT66), .A3(new_n380), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n448), .A2(new_n437), .A3(new_n434), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT35), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n434), .A2(new_n437), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n349), .A2(new_n355), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT79), .B(new_n347), .C1(new_n350), .C2(new_n354), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n458), .A2(KEYINPUT37), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n349), .A2(new_n355), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n358), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n456), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT37), .B1(new_n363), .B2(new_n364), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n465), .A2(KEYINPUT38), .A3(new_n358), .A4(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n467), .A2(new_n443), .A3(new_n442), .A4(new_n360), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n266), .B1(new_n262), .B2(new_n265), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n252), .B1(new_n275), .B2(new_n259), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n470), .A2(new_n471), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n472), .A2(new_n473), .A3(new_n273), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(KEYINPUT40), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n281), .B1(new_n474), .B2(KEYINPUT40), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n371), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n468), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n367), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n444), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n434), .A2(new_n437), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n405), .A2(new_n407), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n447), .A2(new_n454), .B1(new_n478), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G190gat), .B(G218gat), .Z(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT99), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G92gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n270), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT97), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n494), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G99gat), .ZN(new_n501));
  INV_X1    g300(.A(G106gat), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT8), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(G99gat), .B(G106gat), .Z(new_n506));
  INV_X1    g305(.A(KEYINPUT97), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT7), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n494), .A2(new_n499), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(KEYINPUT96), .B2(KEYINPUT7), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT98), .B(G85gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n493), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n503), .B(new_n509), .C1(new_n513), .C2(new_n494), .ZN(new_n514));
  INV_X1    g313(.A(new_n506), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G50gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT15), .B1(new_n518), .B2(G43gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(G43gat), .B2(new_n518), .ZN(new_n520));
  NOR2_X1   g319(.A1(G29gat), .A2(G36gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT14), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527));
  AND2_X1   g326(.A1(KEYINPUT83), .A2(G43gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(KEYINPUT83), .A2(G43gat), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n528), .A2(new_n529), .A3(G50gat), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT84), .B1(new_n518), .B2(G43gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT84), .ZN(new_n532));
  INV_X1    g331(.A(G43gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(G50gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n527), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT85), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(KEYINPUT85), .B(new_n527), .C1(new_n530), .C2(new_n535), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n526), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT14), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n521), .B(new_n541), .ZN(new_n542));
  OAI22_X1  g341(.A1(new_n542), .A2(KEYINPUT82), .B1(new_n523), .B2(new_n524), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n520), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT17), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n517), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n517), .ZN(new_n551));
  AND2_X1   g350(.A1(G232gat), .A2(G233gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT41), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n492), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n517), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n540), .A2(new_n545), .A3(new_n548), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n548), .B1(new_n540), .B2(new_n545), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(new_n553), .A3(new_n551), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n492), .A3(new_n556), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n488), .B1(new_n558), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n490), .A2(KEYINPUT99), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT41), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  NAND3_X1  g368(.A1(new_n558), .A2(new_n564), .A3(new_n488), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n569), .ZN(new_n572));
  INV_X1    g371(.A(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(new_n565), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT101), .ZN(new_n577));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(G211gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT91), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  INV_X1    g386(.A(G71gat), .ZN(new_n588));
  INV_X1    g387(.A(G78gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G57gat), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n591), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n585), .A2(new_n586), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n586), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n587), .B2(new_n584), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n593), .A2(KEYINPUT92), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n601));
  XNOR2_X1  g400(.A(G15gat), .B(G22gat), .ZN(new_n602));
  INV_X1    g401(.A(G1gat), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n603), .A2(KEYINPUT16), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n602), .A2(new_n603), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT86), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT87), .ZN(new_n608));
  XOR2_X1   g407(.A(G15gat), .B(G22gat), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G1gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n602), .A2(new_n604), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n607), .B(G8gat), .C1(new_n612), .C2(KEYINPUT86), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT87), .B1(new_n605), .B2(new_n606), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT86), .ZN(new_n615));
  INV_X1    g414(.A(G8gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n290), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n290), .B1(new_n601), .B2(new_n618), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n583), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(new_n619), .A3(new_n582), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n581), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n627));
  NAND3_X1  g426(.A1(new_n598), .A2(new_n599), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  NAND3_X1  g429(.A1(new_n622), .A2(new_n624), .A3(new_n581), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n625), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n514), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n515), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n514), .A2(new_n641), .A3(new_n506), .ZN(new_n644));
  INV_X1    g443(.A(new_n596), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n598), .A2(new_n510), .A3(new_n516), .A4(new_n599), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G230gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n318), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n647), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n600), .A2(new_n517), .A3(KEYINPUT10), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n640), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n652), .A2(new_n657), .A3(new_n639), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n576), .A2(new_n577), .A3(new_n636), .A4(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n636), .A2(new_n574), .A3(new_n571), .A4(new_n662), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT101), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n486), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n618), .B1(new_n560), .B2(new_n561), .ZN(new_n668));
  NAND2_X1  g467(.A1(G229gat), .A2(G233gat), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n613), .A2(new_n617), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n546), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT89), .B1(new_n670), .B2(new_n546), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT89), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n618), .A2(new_n676), .A3(new_n545), .A4(new_n540), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n677), .A3(new_n671), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n669), .B(KEYINPUT13), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n673), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n668), .A2(new_n669), .A3(new_n671), .A4(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G113gat), .B(G141gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n330), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT11), .B(G169gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT12), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT81), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT81), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n684), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n674), .A2(new_n681), .A3(new_n683), .A4(new_n689), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n667), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n444), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(new_n603), .ZN(G1324gat));
  INV_X1    g499(.A(new_n698), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n616), .B1(new_n701), .B2(new_n371), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT16), .B(G8gat), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n698), .A2(new_n439), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(KEYINPUT42), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n704), .A2(new_n706), .A3(KEYINPUT42), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n704), .B2(KEYINPUT42), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(G1325gat));
  NAND2_X1  g508(.A1(new_n482), .A2(new_n484), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n701), .A2(G15gat), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(G15gat), .B1(new_n701), .B2(new_n408), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1326gat));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n455), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT43), .B(G22gat), .Z(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  NAND2_X1  g516(.A1(new_n447), .A2(new_n454), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n485), .A2(new_n478), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n576), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n636), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n697), .A3(new_n662), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n724), .A2(G29gat), .A3(new_n444), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT45), .Z(new_n726));
  OAI21_X1  g525(.A(KEYINPUT44), .B1(new_n486), .B2(new_n576), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n408), .A2(new_n434), .A3(new_n437), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n439), .A2(new_n444), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(KEYINPUT80), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n371), .B1(new_n443), .B2(new_n442), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT35), .B1(new_n732), .B2(new_n445), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n731), .A2(new_n733), .B1(KEYINPUT35), .B2(new_n453), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n485), .A2(new_n478), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n728), .B(new_n575), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n727), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n723), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n444), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n726), .A2(new_n739), .ZN(G1328gat));
  NOR3_X1   g539(.A1(new_n724), .A2(G36gat), .A3(new_n439), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT46), .ZN(new_n742));
  OAI21_X1  g541(.A(G36gat), .B1(new_n738), .B2(new_n439), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1329gat));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n738), .A2(new_n710), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n528), .A2(new_n529), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n408), .A2(new_n748), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n724), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n745), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  OAI221_X1 g551(.A(KEYINPUT47), .B1(new_n724), .B2(new_n750), .C1(new_n746), .C2(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1330gat));
  OAI21_X1  g553(.A(G50gat), .B1(new_n738), .B2(new_n455), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n720), .A2(new_n518), .A3(new_n481), .A4(new_n723), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n757), .A2(KEYINPUT103), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(KEYINPUT103), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n722), .B1(new_n727), .B2(new_n736), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n518), .B1(new_n763), .B2(new_n481), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n761), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT104), .B1(new_n765), .B2(new_n756), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n767));
  NOR4_X1   g566(.A1(new_n764), .A2(new_n767), .A3(new_n757), .A4(new_n761), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n766), .B2(new_n768), .ZN(G1331gat));
  NOR2_X1   g568(.A1(new_n721), .A2(new_n575), .ZN(new_n770));
  INV_X1    g569(.A(new_n697), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n661), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n770), .B(new_n773), .C1(new_n734), .C2(new_n735), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT105), .ZN(new_n775));
  INV_X1    g574(.A(new_n486), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n770), .A4(new_n773), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n778), .A3(new_n284), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G57gat), .ZN(G1332gat));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n781));
  INV_X1    g580(.A(new_n770), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n486), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n777), .B1(new_n783), .B2(new_n773), .ZN(new_n784));
  NOR4_X1   g583(.A1(new_n486), .A2(KEYINPUT105), .A3(new_n782), .A4(new_n772), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n775), .A2(new_n778), .A3(KEYINPUT106), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n371), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n791));
  XOR2_X1   g590(.A(KEYINPUT49), .B(G64gat), .Z(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(G1333gat));
  NAND4_X1  g592(.A1(new_n786), .A2(G71gat), .A3(new_n711), .A4(new_n787), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n775), .A2(new_n778), .A3(new_n408), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n588), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT50), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n799), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1334gat));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n481), .A3(new_n787), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g602(.A1(new_n697), .A2(new_n636), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n661), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n737), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(new_n444), .A3(new_n512), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n720), .A2(new_n804), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n720), .A2(new_n811), .A3(new_n804), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n661), .A3(new_n812), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n813), .A2(new_n444), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n808), .B1(new_n814), .B2(new_n512), .ZN(G1336gat));
  INV_X1    g614(.A(new_n789), .ZN(new_n816));
  OAI21_X1  g615(.A(G92gat), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n816), .A2(G92gat), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n817), .B(new_n818), .C1(new_n813), .C2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n737), .A2(new_n371), .A3(new_n806), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G92gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n811), .A2(KEYINPUT108), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n720), .B2(new_n804), .ZN(new_n826));
  INV_X1    g625(.A(new_n804), .ZN(new_n827));
  INV_X1    g626(.A(new_n825), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n486), .A2(new_n576), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n661), .B(new_n819), .C1(new_n826), .C2(new_n829), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n822), .B(new_n818), .C1(new_n824), .C2(new_n830), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n439), .B(new_n805), .C1(new_n727), .C2(new_n736), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n832), .B2(new_n493), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT109), .B1(new_n833), .B2(KEYINPUT52), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n821), .B1(new_n831), .B2(new_n834), .ZN(G1337gat));
  OAI21_X1  g634(.A(G99gat), .B1(new_n807), .B2(new_n710), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n408), .A2(new_n501), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n813), .B2(new_n837), .ZN(G1338gat));
  NAND3_X1  g637(.A1(new_n737), .A2(new_n481), .A3(new_n806), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G106gat), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n455), .A2(G106gat), .A3(new_n662), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n810), .A2(new_n812), .A3(new_n841), .ZN(new_n842));
  XOR2_X1   g641(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n826), .A2(new_n829), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n845), .A2(new_n841), .B1(new_n839), .B2(G106gat), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(G1339gat));
  NAND2_X1  g647(.A1(new_n816), .A2(new_n284), .ZN(new_n849));
  INV_X1    g648(.A(new_n660), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n655), .A2(new_n656), .A3(new_n650), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT54), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n657), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n655), .A2(new_n656), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n651), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n639), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n851), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n640), .B1(new_n657), .B2(new_n856), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(KEYINPUT55), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n697), .A2(new_n850), .A3(new_n863), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n679), .A2(new_n675), .A3(new_n671), .A4(new_n677), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n669), .B1(new_n668), .B2(new_n671), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n688), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT111), .B(new_n688), .C1(new_n865), .C2(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n661), .C1(new_n695), .C2(new_n696), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n575), .B1(new_n864), .B2(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n874), .A2(new_n875), .B1(new_n869), .B2(new_n870), .ZN(new_n876));
  AND4_X1   g675(.A1(new_n575), .A2(new_n876), .A3(new_n850), .A4(new_n863), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n721), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n664), .A2(new_n697), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n849), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n438), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n224), .B1(new_n883), .B2(new_n697), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n455), .A2(new_n452), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(G113gat), .A3(new_n771), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n884), .A2(new_n888), .ZN(G1340gat));
  OAI21_X1  g688(.A(G120gat), .B1(new_n882), .B2(new_n662), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n661), .A2(new_n222), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT112), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT113), .Z(G1341gat));
  OR3_X1    g693(.A1(new_n887), .A2(KEYINPUT114), .A3(new_n721), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT114), .B1(new_n887), .B2(new_n721), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n215), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n883), .A2(G127gat), .A3(new_n636), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1342gat));
  AOI21_X1  g698(.A(new_n213), .B1(new_n883), .B2(new_n575), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n444), .B1(new_n878), .B2(new_n880), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n576), .A2(new_n371), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n901), .A2(new_n213), .A3(new_n886), .A4(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n900), .B1(KEYINPUT56), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT115), .B1(new_n903), .B2(KEYINPUT56), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n903), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G1343gat));
  NAND2_X1  g706(.A1(new_n878), .A2(new_n880), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n481), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n849), .A2(new_n711), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT116), .B1(new_n860), .B2(new_n861), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n697), .A3(new_n850), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n575), .B1(new_n914), .B2(new_n872), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n721), .B1(new_n915), .B2(new_n877), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n455), .B1(new_n916), .B2(new_n880), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n910), .B(new_n911), .C1(new_n917), .C2(new_n909), .ZN(new_n918));
  OAI21_X1  g717(.A(G141gat), .B1(new_n918), .B2(new_n771), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n711), .A2(new_n455), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n901), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n921), .A2(new_n203), .A3(new_n697), .A4(new_n816), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT58), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT58), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1344gat));
  INV_X1    g726(.A(new_n918), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT59), .B(new_n243), .C1(new_n928), .C2(new_n661), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n930));
  INV_X1    g729(.A(new_n872), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n859), .A2(new_n862), .A3(new_n850), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n694), .B(KEYINPUT90), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n693), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n576), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n575), .A2(new_n876), .A3(new_n850), .A4(new_n863), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n636), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g736(.A(KEYINPUT57), .B(new_n481), .C1(new_n937), .C2(new_n879), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT118), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n908), .A2(new_n940), .A3(KEYINPUT57), .A4(new_n481), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n663), .A2(new_n665), .A3(new_n771), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT119), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT119), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n663), .A2(new_n665), .A3(new_n945), .A4(new_n771), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n916), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n947), .B2(new_n481), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n661), .B(new_n911), .C1(new_n942), .C2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n930), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n921), .A2(new_n243), .A3(new_n816), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n662), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT117), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n951), .A2(KEYINPUT117), .A3(new_n662), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n929), .A2(new_n950), .B1(new_n954), .B2(new_n955), .ZN(G1345gat));
  NAND2_X1  g755(.A1(new_n636), .A2(G155gat), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT120), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n921), .A2(new_n636), .A3(new_n816), .ZN(new_n959));
  INV_X1    g758(.A(G155gat), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n928), .A2(new_n958), .B1(new_n959), .B2(new_n960), .ZN(G1346gat));
  OAI21_X1  g760(.A(G162gat), .B1(new_n918), .B2(new_n576), .ZN(new_n962));
  INV_X1    g761(.A(G162gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n921), .A2(new_n963), .A3(new_n902), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n962), .A2(KEYINPUT121), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1347gat));
  NAND3_X1  g768(.A1(new_n444), .A2(new_n408), .A3(new_n371), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n970), .A2(KEYINPUT123), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(KEYINPUT123), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n908), .A2(new_n455), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(G169gat), .B1(new_n973), .B2(new_n771), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n284), .B1(new_n878), .B2(new_n880), .ZN(new_n975));
  AND4_X1   g774(.A1(new_n297), .A2(new_n975), .A3(new_n886), .A4(new_n789), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT122), .B1(new_n976), .B2(new_n697), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n975), .A2(new_n886), .A3(new_n789), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n979));
  NOR4_X1   g778(.A1(new_n978), .A2(new_n979), .A3(G169gat), .A4(new_n771), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n974), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g782(.A(KEYINPUT124), .B(new_n974), .C1(new_n977), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1348gat));
  NOR3_X1   g784(.A1(new_n973), .A2(new_n298), .A3(new_n662), .ZN(new_n986));
  INV_X1    g785(.A(new_n978), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(new_n661), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n986), .B1(new_n988), .B2(new_n298), .ZN(G1349gat));
  OAI21_X1  g788(.A(G183gat), .B1(new_n973), .B2(new_n721), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n636), .A2(new_n303), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n990), .B1(new_n978), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g792(.A(G190gat), .B1(new_n973), .B2(new_n576), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT61), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n987), .A2(new_n291), .A3(new_n575), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1351gat));
  AND2_X1   g796(.A1(new_n975), .A2(new_n789), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(new_n920), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n330), .B1(new_n999), .B2(new_n771), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n711), .A2(new_n284), .A3(new_n439), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n771), .A2(new_n330), .ZN(new_n1002));
  OAI211_X1 g801(.A(new_n1001), .B(new_n1002), .C1(new_n942), .C2(new_n948), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1000), .A2(new_n1003), .A3(KEYINPUT125), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT125), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1352gat));
  OAI211_X1 g805(.A(new_n661), .B(new_n1001), .C1(new_n942), .C2(new_n948), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(G204gat), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n998), .A2(new_n331), .A3(new_n661), .A4(new_n920), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g812(.A(new_n1008), .B(new_n1013), .C1(new_n1011), .C2(new_n1009), .ZN(G1353gat));
  NAND4_X1  g813(.A1(new_n998), .A2(new_n579), .A3(new_n636), .A4(new_n920), .ZN(new_n1015));
  OAI211_X1 g814(.A(new_n636), .B(new_n1001), .C1(new_n942), .C2(new_n948), .ZN(new_n1016));
  AND3_X1   g815(.A1(new_n1016), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1017));
  AOI21_X1  g816(.A(KEYINPUT63), .B1(new_n1016), .B2(G211gat), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(G1354gat));
  INV_X1    g818(.A(G218gat), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1020), .B1(new_n999), .B2(new_n576), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1022));
  AND2_X1   g821(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  NOR2_X1   g823(.A1(new_n576), .A2(new_n1020), .ZN(new_n1025));
  OAI211_X1 g824(.A(new_n1001), .B(new_n1025), .C1(new_n942), .C2(new_n948), .ZN(new_n1026));
  INV_X1    g825(.A(new_n1026), .ZN(new_n1027));
  NOR3_X1   g826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1027), .ZN(G1355gat));
endmodule


