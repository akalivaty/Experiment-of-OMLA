//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT86), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT80), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT80), .A3(new_n206), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n206), .A2(KEYINPUT2), .ZN(new_n214));
  AND2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n209), .A2(new_n213), .A3(new_n214), .A4(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n214), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(new_n206), .A3(new_n212), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G211gat), .A2(G218gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n230), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n225), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n224), .A3(new_n236), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n233), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n204), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT87), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT87), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(new_n204), .C1(new_n237), .C2(new_n239), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n230), .B(new_n231), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n236), .B1(new_n244), .B2(KEYINPUT29), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n218), .A2(new_n224), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n238), .A2(new_n234), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n244), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n247), .A2(new_n249), .A3(G228gat), .A4(G233gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n243), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G22gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(G78gat), .B(G106gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT31), .B(G50gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n243), .A2(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n249), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n242), .B1(new_n257), .B2(new_n204), .ZN(new_n258));
  OAI21_X1  g057(.A(G22gat), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n255), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI211_X1 g062(.A(KEYINPUT89), .B(new_n255), .C1(new_n259), .C2(new_n260), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n252), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n252), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT88), .B1(new_n251), .B2(G22gat), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT89), .B1(new_n267), .B2(new_n255), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n261), .A2(new_n262), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT26), .ZN(new_n274));
  NOR2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n275), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT70), .A3(KEYINPUT26), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n275), .B2(new_n274), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n283), .A2(KEYINPUT28), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT28), .B1(new_n283), .B2(new_n284), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n281), .B(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT25), .B1(new_n277), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n288), .A2(KEYINPUT68), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(KEYINPUT68), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n272), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n289), .B1(new_n292), .B2(new_n277), .ZN(new_n293));
  NAND3_X1  g092(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G183gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n284), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n295), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n296), .A2(new_n298), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT67), .B(G176gat), .Z(new_n304));
  NOR2_X1   g103(.A1(new_n288), .A2(G169gat), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n292), .A2(new_n277), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT65), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n294), .A2(new_n308), .B1(new_n297), .B2(new_n284), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n310), .A3(new_n299), .ZN(new_n311));
  NAND4_X1  g110(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n307), .A2(new_n309), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT25), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n287), .B1(new_n303), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT79), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n305), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT68), .B(KEYINPUT23), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n277), .B1(new_n321), .B2(new_n273), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(new_n324), .B1(new_n302), .B2(new_n293), .ZN(new_n325));
  INV_X1    g124(.A(new_n287), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT79), .B(new_n287), .C1(new_n303), .C2(new_n314), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n316), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n233), .B(new_n318), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n316), .B1(new_n327), .B2(new_n328), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n317), .B1(new_n315), .B2(new_n234), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n244), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n335));
  XNOR2_X1  g134(.A(G8gat), .B(G36gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n331), .A2(new_n334), .A3(new_n335), .A4(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n331), .A2(new_n334), .A3(new_n339), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT30), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n339), .B1(new_n331), .B2(new_n334), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G15gat), .B(G43gat), .Z(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT73), .ZN(new_n346));
  XOR2_X1   g145(.A(G71gat), .B(G99gat), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  INV_X1    g149(.A(G113gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G120gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT1), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G127gat), .ZN(new_n357));
  INV_X1    g156(.A(G127gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G134gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n353), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G127gat), .B(G134gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT72), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n351), .A2(G120gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n349), .A2(G113gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n369));
  INV_X1    g168(.A(new_n359), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n362), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n364), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n374), .B(new_n287), .C1(new_n314), .C2(new_n303), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n364), .B(new_n373), .C1(new_n325), .C2(new_n326), .ZN(new_n376));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT64), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT33), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n348), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(KEYINPUT32), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n379), .B(KEYINPUT32), .C1(new_n380), .C2(new_n348), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT75), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n376), .ZN(new_n387));
  INV_X1    g186(.A(new_n378), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n389), .B2(KEYINPUT34), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT34), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n387), .A2(KEYINPUT75), .A3(new_n391), .A4(new_n388), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(KEYINPUT34), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n385), .B(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  XOR2_X1   g195(.A(KEYINPUT95), .B(KEYINPUT35), .Z(new_n397));
  NAND3_X1  g196(.A1(new_n364), .A2(new_n373), .A3(new_n225), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n371), .A2(new_n218), .A3(new_n224), .A4(new_n362), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n400), .A2(KEYINPUT4), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n371), .A2(new_n362), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n238), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n246), .A2(new_n405), .A3(KEYINPUT3), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n404), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n402), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(new_n246), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n400), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n415), .B2(new_n404), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT84), .ZN(new_n419));
  XOR2_X1   g218(.A(G1gat), .B(G29gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n400), .A2(KEYINPUT4), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n364), .A2(new_n373), .A3(new_n225), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n428), .A3(KEYINPUT4), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n425), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT81), .B1(new_n225), .B2(new_n236), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n431), .A2(new_n407), .A3(new_n410), .A4(new_n238), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n430), .A2(new_n432), .A3(new_n403), .A4(new_n413), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n423), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n423), .ZN(new_n437));
  INV_X1    g236(.A(new_n416), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n411), .B2(new_n402), .ZN(new_n439));
  INV_X1    g238(.A(new_n433), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT93), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n423), .B1(new_n417), .B2(new_n433), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT93), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n436), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(KEYINPUT6), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n397), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n271), .A2(new_n344), .A3(new_n396), .A4(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT96), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n417), .A2(new_n433), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT93), .B1(new_n452), .B2(new_n437), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n442), .B(new_n423), .C1(new_n417), .C2(new_n433), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n455), .A2(new_n436), .B1(KEYINPUT6), .B2(new_n444), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n456), .A2(new_n395), .A3(new_n397), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(KEYINPUT96), .A3(new_n344), .A4(new_n271), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT74), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT76), .B1(new_n385), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n394), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT74), .B1(new_n394), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n385), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n441), .A2(new_n435), .A3(new_n434), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n447), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n271), .A2(new_n465), .A3(new_n467), .A4(new_n344), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n451), .A2(new_n458), .B1(KEYINPUT35), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n271), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(new_n467), .A3(new_n344), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n331), .A2(new_n334), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n339), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n244), .B(new_n318), .C1(new_n329), .C2(new_n330), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n233), .B1(new_n332), .B2(new_n333), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(KEYINPUT37), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(new_n446), .A3(new_n447), .A4(new_n341), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(KEYINPUT37), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n476), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT40), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT39), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n430), .A2(new_n432), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT90), .B1(new_n487), .B2(new_n404), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n489));
  AOI211_X1 g288(.A(new_n489), .B(new_n403), .C1(new_n430), .C2(new_n432), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(KEYINPUT91), .A3(new_n423), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n488), .A2(new_n490), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n414), .A2(new_n400), .A3(new_n403), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n486), .B1(new_n494), .B2(new_n495), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT91), .B1(new_n491), .B2(new_n423), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n485), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n443), .A2(new_n445), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n344), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n491), .A2(new_n423), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(KEYINPUT40), .A3(new_n492), .A4(new_n498), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n501), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT94), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n501), .A2(new_n503), .A3(new_n507), .A4(KEYINPUT94), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n484), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n471), .B1(new_n512), .B2(new_n470), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n465), .A2(KEYINPUT36), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n395), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n469), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G113gat), .B(G141gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT97), .B(KEYINPUT11), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT12), .ZN(new_n524));
  NOR2_X1   g323(.A1(KEYINPUT101), .A2(G8gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(G1gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(KEYINPUT101), .A2(G8gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  INV_X1    g331(.A(KEYINPUT100), .ZN(new_n533));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(KEYINPUT99), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(KEYINPUT99), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR3_X1   g339(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n537), .B(new_n538), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n533), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n542), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n544), .A2(KEYINPUT100), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(G29gat), .A2(G36gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n551), .A2(new_n539), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n546), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT98), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT98), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n552), .A2(new_n546), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n532), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n532), .A2(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n562), .B(KEYINPUT13), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n532), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n548), .A2(new_n557), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n566), .B1(new_n548), .B2(new_n557), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n569), .A2(KEYINPUT18), .A3(new_n562), .A4(new_n560), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n562), .A3(new_n560), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n524), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n574), .A3(new_n524), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT102), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT102), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n571), .A2(new_n574), .A3(new_n524), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n575), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G134gat), .B(G162gat), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G99gat), .ZN(new_n586));
  INV_X1    g385(.A(G106gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(KEYINPUT105), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT104), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT104), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(G85gat), .A3(G92gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n595), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT7), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n588), .A2(KEYINPUT105), .A3(new_n589), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n589), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n591), .A2(new_n596), .A3(new_n599), .A4(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n599), .A2(new_n596), .A3(new_n600), .A4(new_n603), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n590), .A2(KEYINPUT105), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n567), .B2(new_n568), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n558), .A2(new_n609), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT106), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT106), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n611), .A2(new_n613), .A3(new_n618), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n615), .B1(new_n611), .B2(new_n613), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n626), .A3(new_n622), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n585), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n626), .B1(new_n620), .B2(new_n622), .ZN(new_n629));
  AOI211_X1 g428(.A(new_n624), .B(new_n621), .C1(new_n617), .C2(new_n619), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n629), .A2(new_n630), .A3(new_n584), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  OR2_X1    g432(.A1(G57gat), .A2(G64gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(G57gat), .A2(G64gat), .ZN(new_n635));
  AND2_X1   g434(.A1(G71gat), .A2(G78gat), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(KEYINPUT9), .ZN(new_n637));
  NOR2_X1   g436(.A1(G71gat), .A2(G78gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n637), .B(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n565), .B1(new_n633), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT103), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n633), .ZN(new_n644));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G127gat), .B(G155gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(G183gat), .B(G211gat), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n643), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n642), .A3(new_n652), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n640), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n609), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n605), .A2(new_n608), .A3(new_n640), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n660), .A2(KEYINPUT107), .A3(new_n661), .A4(new_n663), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G230gat), .A2(G233gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n660), .A2(new_n663), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n669), .ZN(new_n673));
  XOR2_X1   g472(.A(G120gat), .B(G148gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT108), .ZN(new_n675));
  XOR2_X1   g474(.A(G176gat), .B(G204gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n673), .A2(new_n677), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n632), .A2(new_n658), .A3(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n518), .A2(new_n583), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n467), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g485(.A1(new_n518), .A2(new_n583), .ZN(new_n687));
  INV_X1    g486(.A(new_n682), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(KEYINPUT109), .A3(new_n344), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691));
  INV_X1    g490(.A(new_n344), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n683), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694));
  OAI22_X1  g493(.A1(new_n690), .A2(new_n693), .B1(new_n694), .B2(G8gat), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT16), .B(G8gat), .Z(new_n696));
  NAND4_X1  g495(.A1(new_n683), .A2(KEYINPUT42), .A3(new_n692), .A4(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n695), .B(new_n697), .C1(KEYINPUT42), .C2(new_n696), .ZN(G1325gat));
  OR3_X1    g497(.A1(new_n689), .A2(G15gat), .A3(new_n395), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n517), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n514), .A2(KEYINPUT110), .A3(new_n516), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G15gat), .B1(new_n689), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n705), .ZN(G1326gat));
  OAI21_X1  g505(.A(KEYINPUT111), .B1(new_n689), .B2(new_n271), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n683), .A2(new_n708), .A3(new_n470), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT43), .B(G22gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  XNOR2_X1  g511(.A(new_n658), .B(KEYINPUT112), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n580), .A2(new_n575), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n715), .A3(new_n681), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n513), .A2(new_n704), .ZN(new_n717));
  INV_X1    g516(.A(new_n469), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n632), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT44), .B1(new_n518), .B2(new_n632), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n716), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n726), .B2(new_n467), .ZN(new_n727));
  INV_X1    g526(.A(new_n658), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n720), .A2(new_n728), .A3(new_n681), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n467), .A2(G29gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n687), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n733), .ZN(G1328gat));
  INV_X1    g533(.A(G36gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n687), .A2(new_n735), .A3(new_n692), .A4(new_n730), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT46), .Z(new_n737));
  OAI21_X1  g536(.A(G36gat), .B1(new_n726), .B2(new_n344), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1329gat));
  INV_X1    g538(.A(G43gat), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n725), .B2(new_n703), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n395), .A2(G43gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR4_X1   g542(.A1(new_n518), .A2(new_n583), .A3(new_n729), .A4(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n513), .A2(new_n517), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n718), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(new_n582), .A3(new_n730), .A4(new_n742), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT114), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI211_X1 g550(.A(KEYINPUT115), .B(KEYINPUT47), .C1(new_n748), .C2(KEYINPUT114), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n741), .A2(new_n744), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n716), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n747), .B2(new_n720), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n469), .B1(new_n513), .B2(new_n704), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n757), .A2(new_n632), .A3(new_n721), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n703), .B(new_n754), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G43gat), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n750), .B1(new_n744), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT115), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n749), .A2(new_n745), .A3(new_n750), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n760), .A2(new_n763), .A3(new_n748), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n753), .A2(new_n765), .ZN(G1330gat));
  INV_X1    g565(.A(G50gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n271), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n725), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n687), .A2(new_n470), .A3(new_n730), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n767), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(KEYINPUT48), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT48), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1331gat));
  NAND2_X1  g573(.A1(new_n632), .A2(new_n658), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n680), .A2(new_n714), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n757), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n684), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g578(.A(new_n344), .B(KEYINPUT116), .Z(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n783), .B(new_n784), .Z(G1333gat));
  INV_X1    g584(.A(G71gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n777), .A2(new_n786), .A3(new_n396), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n777), .A2(new_n703), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n786), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n777), .A2(new_n470), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g592(.A1(new_n658), .A2(new_n715), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n757), .A2(new_n632), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(KEYINPUT51), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NOR4_X1   g597(.A1(new_n757), .A2(new_n798), .A3(new_n632), .A4(new_n795), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n800), .A2(new_n601), .A3(new_n684), .A4(new_n680), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n795), .A2(new_n681), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n723), .B2(new_n724), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n684), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n801), .B1(new_n601), .B2(new_n805), .ZN(G1336gat));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n798), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n719), .A2(new_n720), .A3(new_n794), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n781), .A2(G92gat), .A3(new_n681), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n602), .B1(new_n804), .B2(new_n692), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n797), .B2(new_n799), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  AOI211_X1 g615(.A(new_n781), .B(new_n803), .C1(new_n723), .C2(new_n724), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n602), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n818), .ZN(G1337gat));
  NAND4_X1  g618(.A1(new_n800), .A2(new_n586), .A3(new_n396), .A4(new_n680), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n804), .A2(new_n703), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n586), .B2(new_n821), .ZN(G1338gat));
  NOR3_X1   g621(.A1(new_n681), .A2(new_n271), .A3(G106gat), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT118), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n808), .A2(new_n810), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n587), .B1(new_n804), .B2(new_n470), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT53), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n797), .B2(new_n799), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  AOI211_X1 g628(.A(new_n271), .B(new_n803), .C1(new_n723), .C2(new_n724), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n587), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(G1339gat));
  NOR2_X1   g631(.A1(new_n682), .A2(new_n715), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n561), .A2(new_n563), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n562), .B1(new_n569), .B2(new_n560), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n523), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n577), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n680), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n668), .A2(new_n670), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT54), .B1(new_n668), .B2(new_n670), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n668), .A2(new_n670), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n671), .A2(KEYINPUT119), .A3(KEYINPUT54), .A4(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n677), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n668), .A2(new_n670), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n843), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT55), .A4(new_n849), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n678), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n839), .B1(new_n854), .B2(new_n714), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n632), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n838), .B1(new_n628), .B2(new_n631), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n854), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n625), .A2(new_n627), .A3(new_n585), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n584), .B1(new_n629), .B2(new_n630), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n837), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n853), .A2(new_n678), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT120), .A4(new_n852), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n856), .A2(new_n859), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n833), .B1(new_n865), .B2(new_n713), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(new_n467), .A3(new_n780), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n271), .A3(new_n396), .ZN(new_n868));
  OAI21_X1  g667(.A(G113gat), .B1(new_n868), .B2(new_n583), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n271), .A2(new_n465), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n715), .A2(new_n351), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT121), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n869), .A2(new_n875), .ZN(G1340gat));
  AOI21_X1  g675(.A(G120gat), .B1(new_n872), .B2(new_n680), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n868), .A2(new_n349), .A3(new_n681), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1341gat));
  NAND3_X1  g678(.A1(new_n872), .A2(new_n358), .A3(new_n658), .ZN(new_n880));
  OAI21_X1  g679(.A(G127gat), .B1(new_n868), .B2(new_n713), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1342gat));
  OAI21_X1  g681(.A(G134gat), .B1(new_n868), .B2(new_n632), .ZN(new_n883));
  NOR4_X1   g682(.A1(new_n866), .A2(new_n467), .A3(new_n692), .A4(new_n632), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n870), .A2(new_n355), .A3(new_n354), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n884), .A2(KEYINPUT56), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(G1343gat));
  NOR2_X1   g687(.A1(new_n703), .A2(new_n271), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT122), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n867), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n583), .A2(G141gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n703), .A2(new_n467), .A3(new_n780), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n859), .A2(new_n864), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n863), .A2(new_n715), .A3(new_n852), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n720), .B1(new_n896), .B2(new_n839), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n713), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n833), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n470), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n470), .A2(KEYINPUT57), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n582), .A2(new_n863), .A3(new_n852), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n720), .B1(new_n903), .B2(new_n839), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n728), .B1(new_n895), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n582), .B(new_n894), .C1(new_n901), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT58), .B1(new_n907), .B2(G141gat), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(KEYINPUT123), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n893), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n894), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n866), .B2(new_n271), .ZN(new_n914));
  INV_X1    g713(.A(new_n906), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n219), .B1(new_n916), .B2(new_n715), .ZN(new_n917));
  AND4_X1   g716(.A1(KEYINPUT123), .A2(new_n867), .A3(new_n890), .A4(new_n892), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT58), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n911), .A2(new_n919), .ZN(G1344gat));
  NAND3_X1  g719(.A1(new_n891), .A2(new_n220), .A3(new_n680), .ZN(new_n921));
  AOI211_X1 g720(.A(KEYINPUT59), .B(new_n220), .C1(new_n916), .C2(new_n680), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT57), .B1(new_n866), .B2(new_n271), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n858), .A2(new_n854), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n728), .B1(new_n904), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n582), .B2(new_n682), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n913), .A3(new_n470), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n924), .A2(new_n928), .A3(new_n680), .A4(new_n894), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n923), .B1(new_n929), .B2(G148gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n921), .B1(new_n922), .B2(new_n930), .ZN(G1345gat));
  NAND3_X1  g730(.A1(new_n891), .A2(new_n210), .A3(new_n658), .ZN(new_n932));
  INV_X1    g731(.A(new_n713), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n916), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n934), .B2(new_n210), .ZN(G1346gat));
  NAND3_X1  g734(.A1(new_n884), .A2(new_n211), .A3(new_n890), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n916), .A2(new_n720), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n211), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n684), .A2(new_n344), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n271), .A2(new_n396), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n900), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(G169gat), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n941), .A2(new_n942), .A3(new_n583), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n866), .B2(new_n684), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n900), .A2(KEYINPUT124), .A3(new_n467), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n871), .A3(new_n780), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n948), .A2(new_n714), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n943), .B1(new_n949), .B2(new_n942), .ZN(G1348gat));
  NOR3_X1   g749(.A1(new_n941), .A2(new_n304), .A3(new_n681), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n948), .A2(new_n681), .ZN(new_n952));
  INV_X1    g751(.A(G176gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(G1349gat));
  AND2_X1   g753(.A1(new_n658), .A2(new_n283), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n947), .A2(new_n871), .A3(new_n780), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n900), .A2(new_n933), .A3(new_n940), .ZN(new_n957));
  AOI22_X1  g756(.A1(new_n957), .A2(G183gat), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n958));
  OR2_X1    g757(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1350gat));
  OAI21_X1  g761(.A(G190gat), .B1(new_n941), .B2(new_n632), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n720), .A2(new_n284), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n948), .B2(new_n965), .ZN(G1351gat));
  INV_X1    g765(.A(new_n889), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n781), .B(new_n967), .C1(new_n945), .C2(new_n946), .ZN(new_n968));
  AOI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n715), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n924), .A2(new_n928), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n704), .A2(new_n939), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT126), .Z(new_n972));
  AND4_X1   g771(.A1(G197gat), .A2(new_n970), .A3(new_n582), .A4(new_n972), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n969), .A2(new_n973), .ZN(G1352gat));
  XOR2_X1   g773(.A(KEYINPUT127), .B(G204gat), .Z(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n681), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT62), .B1(new_n968), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n866), .A2(new_n944), .A3(new_n684), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT124), .B1(new_n900), .B2(new_n467), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n780), .B(new_n889), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n982));
  INV_X1    g781(.A(new_n977), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n970), .A2(new_n680), .A3(new_n972), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n978), .A2(new_n984), .B1(new_n985), .B2(new_n975), .ZN(G1353gat));
  NAND4_X1  g785(.A1(new_n972), .A2(new_n924), .A3(new_n658), .A4(new_n928), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n989));
  OR2_X1    g788(.A1(new_n728), .A2(G211gat), .ZN(new_n990));
  OAI22_X1  g789(.A1(new_n988), .A2(new_n989), .B1(new_n981), .B2(new_n990), .ZN(G1354gat));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n720), .A3(new_n972), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G218gat), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n632), .A2(G218gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n981), .B2(new_n994), .ZN(G1355gat));
endmodule


