//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G237), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT70), .ZN(new_n191));
  OAI211_X1 g005(.A(G214), .B(new_n187), .C1(new_n189), .C2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(KEYINPUT70), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(G237), .ZN(new_n197));
  AOI21_X1  g011(.A(G953), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(G143), .A3(G214), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n195), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT86), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT17), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n194), .A2(new_n203), .A3(new_n199), .A4(new_n195), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n192), .A2(new_n193), .ZN(new_n205));
  AOI21_X1  g019(.A(G143), .B1(new_n198), .B2(G214), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n201), .A2(new_n202), .A3(new_n204), .A4(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT72), .B(G125), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n212));
  INV_X1    g026(.A(G140), .ZN(new_n213));
  INV_X1    g027(.A(G125), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT72), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT72), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G125), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(G125), .A2(G140), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n212), .B(KEYINPUT16), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n219), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n209), .B2(new_n213), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n212), .B1(new_n223), .B2(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n211), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n207), .A2(new_n202), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n215), .A2(new_n217), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n219), .B1(new_n229), .B2(G140), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT73), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n220), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(G146), .A3(new_n211), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n208), .A2(new_n227), .A3(new_n228), .A4(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G113), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G125), .B(G140), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(KEYINPUT74), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n226), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n226), .B2(new_n223), .ZN(new_n242));
  OAI211_X1 g056(.A(KEYINPUT18), .B(G131), .C1(new_n205), .C2(new_n206), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT18), .A2(G131), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n194), .A2(new_n199), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n235), .A2(new_n238), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n235), .A2(KEYINPUT87), .A3(new_n238), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  MUX2_X1   g065(.A(new_n240), .B(new_n230), .S(KEYINPUT19), .Z(new_n252));
  OAI21_X1  g066(.A(new_n234), .B1(new_n252), .B2(G146), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n201), .A2(new_n204), .A3(new_n207), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n246), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n238), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n259));
  NOR2_X1   g073(.A1(G475), .A2(G902), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n249), .A2(new_n250), .B1(new_n256), .B2(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(new_n260), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT20), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G902), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n249), .A2(new_n250), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n238), .B1(new_n235), .B2(new_n246), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G475), .ZN(new_n270));
  NAND2_X1  g084(.A1(G234), .A2(G237), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n271), .A2(G952), .A3(new_n187), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n271), .A2(G902), .A3(G953), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT21), .B(G898), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT14), .ZN(new_n277));
  INV_X1    g091(.A(G116), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(G122), .ZN(new_n279));
  INV_X1    g093(.A(G122), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G116), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(KEYINPUT90), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n277), .B1(new_n278), .B2(G122), .ZN(new_n283));
  OAI221_X1 g097(.A(G107), .B1(KEYINPUT90), .B2(new_n279), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G107), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(G122), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n281), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n281), .B2(new_n286), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(G128), .B(G143), .ZN(new_n292));
  INV_X1    g106(.A(G134), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n284), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n293), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n289), .A2(new_n285), .A3(new_n290), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n281), .A2(new_n286), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT88), .ZN(new_n299));
  AOI21_X1  g113(.A(G107), .B1(new_n299), .B2(new_n288), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n296), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT13), .B1(new_n193), .B2(G128), .ZN(new_n302));
  INV_X1    g116(.A(G128), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(G143), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n304), .A2(KEYINPUT89), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n303), .A2(G143), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n304), .A2(KEYINPUT89), .B1(KEYINPUT13), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n293), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n295), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  INV_X1    g124(.A(G217), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n310), .A2(new_n311), .A3(G953), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n295), .B(new_n312), .C1(new_n301), .C2(new_n308), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n266), .ZN(new_n317));
  INV_X1    g131(.A(G478), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT15), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n317), .B(new_n319), .Z(new_n320));
  NAND4_X1  g134(.A1(new_n265), .A2(new_n270), .A3(new_n276), .A4(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G140), .ZN(new_n322));
  INV_X1    g136(.A(G227), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G953), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n226), .A2(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n193), .A2(G146), .ZN(new_n329));
  AND4_X1   g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(G128), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n331), .A2(G128), .B1(new_n328), .B2(new_n329), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n285), .A3(G104), .ZN(new_n336));
  INV_X1    g150(.A(G101), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n237), .A2(G107), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n334), .A2(new_n336), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n237), .A2(G107), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n285), .A2(G104), .ZN(new_n341));
  OAI21_X1  g155(.A(G101), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT79), .B1(new_n333), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n339), .A2(new_n342), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n331), .A2(G128), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n328), .A2(new_n329), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G143), .B(G146), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(G128), .A3(new_n331), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n333), .A2(new_n343), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n344), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT11), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n293), .B2(G137), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n293), .A2(G137), .ZN(new_n358));
  INV_X1    g172(.A(G137), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT11), .A3(G134), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n195), .A2(KEYINPUT67), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(new_n357), .A3(new_n358), .A4(new_n360), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n355), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT12), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n355), .A2(KEYINPUT12), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT77), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n334), .A2(new_n336), .A3(new_n374), .A4(new_n338), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(G101), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n373), .A2(G101), .A3(new_n375), .A4(new_n378), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n339), .A2(new_n377), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(KEYINPUT0), .A2(G128), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n328), .A2(new_n329), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT66), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT66), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n328), .A2(new_n329), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT0), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n303), .A3(KEYINPUT65), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT65), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(KEYINPUT0), .B2(G128), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n385), .B1(new_n328), .B2(new_n329), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n387), .A2(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n384), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n363), .A2(new_n365), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT10), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n344), .A2(new_n399), .A3(new_n353), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n345), .A2(new_n351), .A3(KEYINPUT10), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n397), .A2(new_n398), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n326), .B1(new_n371), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n395), .A2(new_n394), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n388), .B1(new_n349), .B2(new_n385), .ZN(new_n406));
  INV_X1    g220(.A(new_n389), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n382), .B1(new_n376), .B2(new_n379), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(new_n381), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n366), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n411), .A2(new_n402), .A3(new_n326), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT80), .B1(new_n403), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT80), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n402), .A3(new_n326), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n404), .A2(new_n410), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n398), .A2(new_n416), .B1(new_n369), .B2(new_n370), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n414), .B(new_n415), .C1(new_n417), .C2(new_n326), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(G469), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n371), .A2(new_n326), .A3(new_n402), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n326), .B1(new_n411), .B2(new_n402), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(KEYINPUT81), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n424));
  AOI211_X1 g238(.A(new_n424), .B(new_n326), .C1(new_n411), .C2(new_n402), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n420), .B(new_n266), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(G469), .A2(G902), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G221), .B1(new_n310), .B2(G902), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n429), .B(KEYINPUT76), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n321), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G122), .ZN(new_n434));
  XOR2_X1   g248(.A(G116), .B(G119), .Z(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT2), .B(G113), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G119), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n440), .A3(G116), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G113), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n345), .B(new_n437), .C1(new_n439), .C2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n435), .B(new_n436), .Z(new_n445));
  OAI211_X1 g259(.A(new_n434), .B(new_n443), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n434), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n409), .B2(new_n381), .ZN(new_n448));
  INV_X1    g262(.A(new_n443), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n446), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  OAI221_X1 g268(.A(new_n447), .B1(new_n451), .B2(new_n452), .C1(new_n448), .C2(new_n449), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n351), .A2(new_n209), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n408), .B2(new_n209), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n187), .A2(G224), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT83), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT83), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n454), .A2(new_n462), .A3(new_n455), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(new_n446), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n458), .A2(KEYINPUT7), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n457), .B(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n434), .B(KEYINPUT8), .Z(new_n469));
  OAI21_X1  g283(.A(new_n437), .B1(new_n439), .B2(new_n442), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n343), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n471), .B2(new_n443), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(KEYINPUT84), .B(new_n469), .C1(new_n471), .C2(new_n443), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n466), .B1(new_n476), .B2(KEYINPUT85), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n468), .B(new_n478), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n464), .A2(new_n465), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n465), .B1(new_n464), .B2(new_n480), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G214), .B1(G237), .B2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n311), .B1(G234), .B2(new_n266), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT75), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT22), .B(G137), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT23), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n440), .B2(G128), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n303), .A2(KEYINPUT23), .A3(G119), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n494), .B(new_n495), .C1(G119), .C2(new_n303), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G110), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT24), .B(G110), .Z(new_n498));
  XNOR2_X1  g312(.A(G119), .B(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n227), .B2(new_n234), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n226), .B(new_n210), .C1(new_n232), .C2(new_n220), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n496), .A2(G110), .B1(new_n499), .B2(new_n498), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n241), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n492), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n501), .ZN(new_n508));
  AOI21_X1  g322(.A(G146), .B1(new_n233), .B2(new_n211), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(new_n503), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n234), .A2(new_n504), .A3(new_n241), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n491), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT25), .B1(new_n513), .B2(new_n266), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT25), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n515), .B(G902), .C1(new_n507), .C2(new_n512), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n487), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n513), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n487), .A2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n357), .A2(new_n360), .A3(new_n195), .A4(new_n358), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n359), .A2(G134), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n293), .A2(G137), .ZN(new_n524));
  OAI21_X1  g338(.A(G131), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT69), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT69), .B1(new_n522), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n351), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n396), .A2(new_n529), .A3(new_n366), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n529), .B1(new_n396), .B2(new_n366), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n445), .B(new_n528), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n198), .A2(G210), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT27), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT27), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n198), .A2(new_n535), .A3(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT26), .B(G101), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n534), .B2(new_n536), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n532), .A2(KEYINPUT71), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT71), .B1(new_n532), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n445), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n351), .A2(new_n525), .A3(new_n522), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n398), .B2(new_n408), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n544), .B(new_n548), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT31), .B1(new_n543), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n532), .A2(new_n540), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT71), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n532), .A2(KEYINPUT71), .A3(new_n540), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n555), .A2(KEYINPUT31), .A3(new_n551), .A4(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT28), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n546), .A2(new_n544), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n532), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n544), .B1(new_n396), .B2(new_n366), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT28), .B1(new_n562), .B2(new_n528), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n552), .A2(new_n558), .B1(new_n564), .B2(new_n540), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n564), .A2(new_n540), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n555), .A2(new_n551), .A3(new_n556), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n569), .B1(new_n572), .B2(new_n557), .ZN(new_n573));
  INV_X1    g387(.A(new_n567), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT32), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n564), .A2(new_n540), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT29), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n551), .A2(new_n532), .ZN(new_n580));
  INV_X1    g394(.A(new_n540), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n549), .A2(new_n544), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n559), .B1(new_n584), .B2(new_n532), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(new_n563), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n581), .A2(new_n579), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n577), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n521), .B1(new_n576), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n433), .A2(new_n486), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  AND2_X1   g407(.A1(new_n428), .A2(new_n431), .ZN(new_n594));
  OAI21_X1  g408(.A(G472), .B1(new_n573), .B2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n565), .A2(new_n567), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n487), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n502), .A2(new_n506), .A3(new_n492), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n491), .B1(new_n510), .B2(new_n511), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n266), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n515), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n513), .A2(KEYINPUT25), .A3(new_n266), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n518), .A2(new_n520), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n594), .A2(new_n597), .A3(KEYINPUT91), .A4(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT91), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n596), .A3(new_n595), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(new_n432), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n611), .B(KEYINPUT92), .Z(new_n612));
  NAND2_X1  g426(.A1(new_n464), .A2(new_n480), .ZN(new_n613));
  INV_X1    g427(.A(new_n465), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n464), .A2(new_n465), .A3(new_n480), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(KEYINPUT93), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n485), .B1(new_n482), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n261), .A2(new_n264), .B1(new_n269), .B2(G475), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n318), .A2(G902), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n314), .A2(new_n624), .A3(new_n315), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n624), .B1(new_n314), .B2(new_n315), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n622), .B(new_n623), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n623), .ZN(new_n629));
  INV_X1    g443(.A(new_n627), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n625), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT94), .B1(new_n317), .B2(new_n318), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n621), .A2(new_n634), .A3(new_n275), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n612), .A2(new_n620), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G104), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  INV_X1    g453(.A(new_n320), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n621), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n612), .A2(new_n276), .A3(new_n620), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NAND2_X1  g459(.A1(new_n595), .A2(new_n596), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT97), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n510), .A2(new_n647), .A3(new_n511), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n647), .B1(new_n510), .B2(new_n511), .ZN(new_n650));
  OAI22_X1  g464(.A1(new_n649), .A2(new_n650), .B1(KEYINPUT36), .B2(new_n491), .ZN(new_n651));
  INV_X1    g465(.A(new_n650), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n491), .A2(KEYINPUT36), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n648), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n519), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n517), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n517), .A2(new_n656), .A3(KEYINPUT98), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n646), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n433), .A2(new_n661), .A3(new_n486), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  AOI21_X1  g478(.A(new_n520), .B1(new_n651), .B2(new_n654), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n604), .A2(new_n658), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT98), .B1(new_n517), .B2(new_n656), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n589), .B1(new_n568), .B2(new_n575), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n668), .A2(new_n669), .A3(new_n432), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n620), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n273), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n272), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n641), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XOR2_X1   g493(.A(new_n483), .B(KEYINPUT38), .Z(new_n680));
  INV_X1    g494(.A(new_n532), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT68), .B1(new_n398), .B2(new_n408), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n396), .A2(new_n529), .A3(new_n366), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n445), .B1(new_n684), .B2(new_n528), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n581), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n570), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n687), .B2(G902), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n576), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n320), .B1(new_n265), .B2(new_n270), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n484), .A2(new_n689), .A3(new_n668), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n675), .B(KEYINPUT39), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n428), .A2(new_n431), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n680), .A2(new_n691), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  NAND2_X1  g511(.A1(new_n265), .A2(new_n270), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT95), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n633), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n700), .A3(new_n675), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n671), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  OAI21_X1  g518(.A(new_n266), .B1(new_n423), .B2(new_n425), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n706), .A2(new_n426), .A3(new_n429), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n620), .A2(new_n635), .A3(new_n591), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND4_X1  g524(.A1(new_n706), .A2(new_n276), .A3(new_n426), .A4(new_n429), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n620), .A2(new_n591), .A3(new_n642), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NAND3_X1  g528(.A1(new_n617), .A2(new_n707), .A3(new_n619), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n668), .A2(new_n669), .A3(new_n321), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n617), .A2(new_n707), .A3(new_n619), .A4(KEYINPUT99), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT100), .A4(new_n719), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  AND3_X1   g539(.A1(new_n690), .A2(new_n617), .A3(new_n619), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT28), .B1(new_n685), .B2(new_n681), .ZN(new_n727));
  INV_X1    g541(.A(new_n563), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n540), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n552), .B2(new_n558), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n567), .B(KEYINPUT101), .Z(new_n732));
  AOI21_X1  g546(.A(KEYINPUT102), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n729), .B1(new_n572), .B2(new_n557), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n735));
  INV_X1    g549(.A(new_n732), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n606), .B(new_n595), .C1(new_n733), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n711), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n726), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NAND3_X1  g555(.A1(new_n731), .A2(KEYINPUT102), .A3(new_n732), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n735), .B1(new_n734), .B2(new_n736), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n744), .B(new_n595), .C1(new_n667), .C2(new_n666), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n701), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n717), .A3(new_n719), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NAND2_X1  g562(.A1(new_n483), .A2(new_n484), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n749), .A2(new_n669), .A3(new_n521), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n415), .B1(new_n417), .B2(new_n326), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n426), .B(new_n427), .C1(new_n420), .C2(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(new_n429), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n750), .A2(KEYINPUT42), .A3(new_n702), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n481), .A2(new_n482), .A3(new_n485), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n591), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n755), .B1(new_n757), .B2(new_n701), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT103), .B(G131), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G33));
  INV_X1    g575(.A(new_n677), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n757), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT104), .B(G134), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G36));
  AOI22_X1  g579(.A1(new_n659), .A2(new_n660), .B1(new_n595), .B2(new_n596), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT43), .B1(new_n698), .B2(new_n634), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n621), .A2(new_n700), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n749), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n413), .B2(new_n418), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  OAI21_X1  g588(.A(G469), .B1(new_n751), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n427), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(KEYINPUT46), .B(new_n427), .C1(new_n773), .C2(new_n775), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n426), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n780), .A2(new_n429), .A3(new_n692), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT44), .A4(new_n769), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n772), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n429), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n780), .A2(KEYINPUT47), .A3(new_n429), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n702), .A2(new_n669), .A3(new_n521), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n756), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NAND3_X1  g606(.A1(new_n708), .A2(new_n713), .A3(new_n740), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n698), .A2(new_n700), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n641), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n484), .B(new_n276), .C1(new_n481), .C2(new_n482), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n607), .A2(new_n795), .A3(new_n610), .A4(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n486), .B(new_n433), .C1(new_n661), .C2(new_n591), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n793), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n746), .A2(new_n753), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n621), .A2(new_n320), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n670), .A2(new_n804), .A3(new_n675), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n756), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n763), .B1(new_n754), .B2(new_n758), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n801), .A2(new_n724), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n670), .B(new_n620), .C1(new_n702), .C2(new_n677), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n675), .B(KEYINPUT106), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n657), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n726), .A2(new_n689), .A3(new_n753), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n747), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n810), .A2(new_n747), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n809), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(KEYINPUT107), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT107), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n815), .A2(new_n823), .A3(new_n817), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n809), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n821), .B1(new_n825), .B2(KEYINPUT53), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n724), .A2(new_n801), .A3(new_n808), .A4(new_n807), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n815), .A2(new_n823), .A3(new_n817), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n823), .B1(new_n815), .B2(new_n817), .ZN(new_n830));
  OAI211_X1 g644(.A(KEYINPUT53), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  XOR2_X1   g645(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n832));
  OAI21_X1  g646(.A(new_n819), .B1(new_n809), .B2(new_n818), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT109), .ZN(new_n835));
  INV_X1    g649(.A(new_n707), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n749), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n767), .A2(new_n272), .A3(new_n769), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT110), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n767), .A2(new_n841), .A3(new_n769), .A4(new_n272), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n838), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n745), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n689), .A2(new_n521), .A3(new_n674), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n837), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n621), .A2(new_n634), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n845), .A2(KEYINPUT112), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT112), .B1(new_n845), .B2(new_n850), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT50), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n738), .B1(new_n840), .B2(new_n842), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n485), .B1(new_n854), .B2(KEYINPUT50), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n680), .A2(new_n836), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n855), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n706), .A2(new_n426), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n430), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n787), .A2(new_n788), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n787), .A2(KEYINPUT113), .A3(new_n788), .A4(new_n862), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n756), .A3(new_n856), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n856), .A2(new_n858), .A3(new_n855), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n860), .A2(new_n867), .A3(KEYINPUT51), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT48), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n843), .A2(new_n872), .A3(new_n591), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n843), .B2(new_n591), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(KEYINPUT48), .A3(new_n873), .ZN(new_n878));
  OAI211_X1 g692(.A(G952), .B(new_n187), .C1(new_n847), .C2(new_n794), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n717), .A2(new_n719), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n881), .B2(new_n856), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n868), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n859), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n856), .A2(new_n863), .A3(new_n756), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n886), .A2(new_n845), .A3(new_n850), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT51), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n870), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT109), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n831), .A2(new_n890), .A3(new_n832), .A4(new_n833), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n827), .A2(new_n835), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(G952), .A2(G953), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n606), .A2(new_n484), .A3(new_n431), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT105), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n689), .ZN(new_n897));
  INV_X1    g711(.A(new_n680), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n698), .A2(new_n634), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n861), .B(KEYINPUT49), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n897), .A2(new_n898), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n894), .A2(new_n901), .ZN(G75));
  AOI21_X1  g716(.A(new_n266), .B1(new_n831), .B2(new_n833), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(G210), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n454), .A2(new_n455), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n459), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n905), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n904), .A2(new_n905), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n187), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n904), .B2(new_n905), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(G51));
  NOR2_X1   g731(.A1(new_n773), .A2(new_n775), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n903), .A2(KEYINPUT116), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT116), .B1(new_n903), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n427), .B(KEYINPUT57), .Z(new_n922));
  AND3_X1   g736(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n832), .B1(new_n831), .B2(new_n833), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n423), .A2(new_n425), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n913), .B1(new_n921), .B2(new_n927), .ZN(G54));
  NAND2_X1  g742(.A1(new_n831), .A2(new_n833), .ZN(new_n929));
  AND2_X1   g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n929), .A2(G902), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n914), .B1(new_n931), .B2(new_n258), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n929), .A2(G902), .A3(new_n258), .A4(new_n930), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT117), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n933), .A2(KEYINPUT117), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(G60));
  NOR2_X1   g750(.A1(new_n626), .A2(new_n627), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n923), .B2(new_n924), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n914), .ZN(new_n942));
  INV_X1    g756(.A(new_n939), .ZN(new_n943));
  INV_X1    g757(.A(new_n835), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n820), .B1(new_n945), .B2(new_n819), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n891), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n943), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n942), .B1(new_n949), .B2(new_n937), .ZN(G63));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT119), .ZN(new_n953));
  XNOR2_X1  g767(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n831), .B2(new_n833), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n655), .B(KEYINPUT120), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n914), .B1(new_n957), .B2(new_n513), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n951), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n957), .A2(new_n513), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n914), .A4(new_n959), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(G66));
  INV_X1    g779(.A(G224), .ZN(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n274), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n801), .A2(new_n724), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(G953), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(KEYINPUT121), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT121), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n968), .A2(new_n971), .A3(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n967), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT122), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n187), .A2(G898), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n454), .B2(new_n455), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n977), .B(new_n967), .C1(new_n970), .C2(new_n972), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n974), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n974), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G69));
  INV_X1    g795(.A(new_n693), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n795), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n591), .A2(new_n756), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT124), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n693), .B1(new_n794), .B2(new_n641), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n750), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n989), .A2(KEYINPUT125), .A3(new_n783), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT125), .B1(new_n989), .B2(new_n783), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n791), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n696), .A2(new_n747), .A3(new_n810), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT62), .ZN(new_n994));
  OAI21_X1  g808(.A(KEYINPUT126), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n989), .A2(new_n783), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n989), .A2(KEYINPUT125), .A3(new_n783), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n993), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .A4(new_n791), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n995), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n252), .B(KEYINPUT123), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1005), .A2(new_n187), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(new_n323), .B2(G953), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n781), .A2(new_n591), .A3(new_n726), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n791), .A2(new_n783), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n808), .A2(new_n747), .A3(new_n810), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1010), .B1(new_n1014), .B2(G953), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n672), .B1(new_n1008), .B2(new_n323), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1009), .B(new_n1015), .C1(new_n187), .C2(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1020), .B1(new_n1014), .B2(new_n968), .ZN(new_n1021));
  INV_X1    g835(.A(new_n580), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n581), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n914), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n995), .A2(new_n968), .A3(new_n1004), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n1019), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1022), .A2(new_n581), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1020), .B1(new_n582), .B2(new_n570), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n826), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1030), .ZN(new_n1032));
  OAI21_X1  g846(.A(KEYINPUT127), .B1(new_n946), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n1028), .A2(new_n1034), .ZN(G57));
endmodule


