//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n441, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n463), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n463), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  AND2_X1   g056(.A1(new_n466), .A2(new_n468), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n467), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT67), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n467), .A3(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n476), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n466), .A2(G138), .A3(new_n467), .A4(new_n468), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n510), .A2(new_n511), .A3(new_n516), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n515), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n518), .A2(G51), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n525), .A2(new_n526), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n520), .A2(G89), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n514), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n518), .A2(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n521), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n510), .A2(new_n511), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(KEYINPUT70), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(KEYINPUT70), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n520), .A2(G81), .B1(new_n518), .B2(G43), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT71), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n545), .A2(new_n550), .A3(new_n546), .A4(new_n547), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n518), .A2(new_n559), .A3(G53), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n517), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n560), .A2(new_n562), .B1(G91), .B2(new_n520), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n510), .A2(G65), .A3(new_n511), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT72), .B1(new_n566), .B2(G651), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n568));
  AOI211_X1 g143(.A(new_n568), .B(new_n514), .C1(new_n564), .C2(new_n565), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n563), .B1(new_n567), .B2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  OAI221_X1 g147(.A(new_n519), .B1(new_n521), .B2(new_n522), .C1(new_n513), .C2(new_n514), .ZN(G303));
  NAND4_X1  g148(.A1(new_n510), .A2(G87), .A3(new_n511), .A4(new_n516), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(G74), .B1(new_n510), .B2(new_n511), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n514), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT73), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT73), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n541), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G48), .B2(new_n518), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n520), .A2(G86), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n520), .A2(KEYINPUT74), .A3(G86), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n514), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n520), .A2(G85), .B1(new_n518), .B2(G47), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(new_n520), .A2(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n541), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G171), .ZN(G284));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G171), .ZN(G321));
  NOR2_X1   g182(.A1(G168), .A2(new_n604), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT75), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(KEYINPUT75), .B2(new_n608), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(KEYINPUT75), .B2(new_n608), .ZN(G280));
  INV_X1    g189(.A(new_n603), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n552), .B2(G868), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n484), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n487), .A2(G135), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n624), .A2(new_n467), .A3(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n467), .B2(G111), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n622), .B(new_n623), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  INV_X1    g204(.A(new_n476), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n470), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n631), .B(new_n632), .Z(new_n633));
  XOR2_X1   g208(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n629), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT79), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2443), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT80), .ZN(new_n653));
  OR3_X1    g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n651), .B1(new_n650), .B2(new_n653), .ZN(new_n655));
  INV_X1    g230(.A(G14), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n650), .B2(new_n653), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT18), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(KEYINPUT82), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(new_n660), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n660), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n661), .B(KEYINPUT17), .Z(new_n668));
  OAI21_X1  g243(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n665), .A2(new_n661), .A3(new_n660), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT83), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n679), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n680), .A2(KEYINPUT20), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(new_n677), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n683), .B(new_n685), .C1(KEYINPUT20), .C2(new_n680), .ZN(new_n686));
  INV_X1    g261(.A(G1991), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n688), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n690), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n691), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n691), .B2(new_n695), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G4), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n615), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT93), .B(G1348), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(KEYINPUT84), .A2(G29), .ZN(new_n706));
  NOR2_X1   g281(.A1(KEYINPUT84), .A2(G29), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G35), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT100), .Z(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT29), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n705), .B1(G2090), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G29), .A2(G32), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n487), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n484), .A2(G129), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT26), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n720), .A2(new_n721), .B1(G105), .B2(new_n470), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n716), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n715), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT27), .B(G1996), .Z(new_n726));
  NOR2_X1   g301(.A1(G5), .A2(G16), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G171), .B2(G16), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n725), .A2(new_n726), .B1(G1961), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n726), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT24), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(G34), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(G34), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n709), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n480), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n730), .B1(new_n731), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G21), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G168), .B2(G16), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(G1966), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT30), .B(G28), .ZN(new_n742));
  OR2_X1    g317(.A1(KEYINPUT31), .A2(G11), .ZN(new_n743));
  NAND2_X1  g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n742), .A2(new_n736), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n628), .B2(new_n709), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n740), .A2(G1966), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n728), .A2(G1961), .B1(new_n731), .B2(new_n737), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR4_X1   g325(.A1(new_n714), .A2(new_n729), .A3(new_n738), .A4(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n736), .A2(G33), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n487), .A2(G139), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT97), .Z(new_n754));
  AOI22_X1  g329(.A1(new_n630), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT98), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n467), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n756), .B2(new_n755), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n470), .A2(G103), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n754), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n752), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G2072), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n709), .A2(G26), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT28), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n484), .A2(G128), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n487), .A2(G140), .ZN(new_n768));
  OR2_X1    g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT95), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n766), .B1(new_n772), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n764), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n700), .A2(G19), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n552), .B2(new_n700), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT94), .B(G1341), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n709), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n709), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT99), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2078), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n751), .A2(new_n776), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT103), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n713), .A2(G2090), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT101), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT23), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n700), .A2(G20), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n789), .B(new_n790), .C1(G299), .C2(G16), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT102), .B(G1956), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n786), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n788), .A2(new_n786), .A3(new_n794), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n785), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n700), .A2(G22), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT89), .Z(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G166), .B2(new_n700), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1971), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G23), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT87), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n577), .B2(new_n700), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT33), .B(G1976), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT88), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  MUX2_X1   g383(.A(G6), .B(G305), .S(G16), .Z(new_n809));
  XOR2_X1   g384(.A(KEYINPUT32), .B(G1981), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT90), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n808), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT34), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n816), .A2(new_n817), .B1(KEYINPUT92), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(new_n817), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n487), .A2(KEYINPUT85), .A3(G131), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n484), .A2(G119), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT85), .ZN(new_n824));
  INV_X1    g399(.A(G131), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n486), .B2(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(G95), .A2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n827), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT86), .Z(new_n829));
  NAND4_X1  g404(.A1(new_n822), .A2(new_n823), .A3(new_n826), .A4(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G25), .B(new_n830), .S(new_n708), .Z(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n700), .A2(G24), .ZN(new_n834));
  INV_X1    g409(.A(G290), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n700), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1986), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n820), .A2(new_n821), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT34), .B1(new_n813), .B2(new_n815), .ZN(new_n840));
  INV_X1    g415(.A(new_n838), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT91), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n819), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT92), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n797), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n819), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n821), .B1(new_n820), .B2(new_n838), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n840), .A2(KEYINPUT91), .A3(new_n841), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n845), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n847), .A2(new_n852), .ZN(G311));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n845), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n843), .A2(new_n846), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n855), .A3(new_n797), .ZN(G150));
  AOI22_X1  g431(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(new_n514), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n520), .A2(G93), .B1(new_n518), .B2(G55), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n860), .B1(new_n549), .B2(new_n551), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n860), .A2(new_n548), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT39), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n603), .A2(new_n616), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n861), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n868), .A2(new_n870), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n864), .B1(new_n872), .B2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n628), .B(new_n480), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n487), .A2(G142), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT107), .ZN(new_n877));
  INV_X1    g452(.A(G130), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n467), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI22_X1  g455(.A1(new_n483), .A2(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(new_n830), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n830), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n885));
  INV_X1    g460(.A(new_n496), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n499), .A2(new_n888), .A3(new_n501), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n499), .B2(new_n501), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n883), .A2(new_n884), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n883), .B2(new_n884), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n893), .A2(new_n772), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n772), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n883), .A2(new_n884), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n502), .A2(KEYINPUT105), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n499), .A2(new_n888), .A3(new_n501), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n498), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n896), .B1(new_n901), .B2(new_n892), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n875), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n772), .B1(new_n893), .B2(new_n894), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n896), .A3(new_n892), .ZN(new_n905));
  INV_X1    g480(.A(new_n875), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n762), .A2(KEYINPUT106), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(new_n633), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n633), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n492), .B(new_n723), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n903), .A2(new_n907), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n903), .B2(new_n907), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n919), .A2(KEYINPUT40), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT40), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(G395));
  NAND2_X1  g498(.A1(new_n615), .A2(G299), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n603), .A2(new_n610), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n867), .A2(new_n618), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n867), .A2(new_n618), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n928), .A2(new_n929), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n931), .B(new_n932), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n835), .A2(new_n577), .ZN(new_n940));
  NAND2_X1  g515(.A1(G290), .A2(new_n578), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT108), .ZN(new_n943));
  XNOR2_X1  g518(.A(G166), .B(G305), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n940), .A2(new_n946), .A3(new_n941), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n938), .A2(new_n937), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT42), .B1(new_n950), .B2(new_n930), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n939), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n939), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g528(.A(G868), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G868), .B2(new_n860), .ZN(G295));
  OAI21_X1  g530(.A(new_n954), .B1(G868), .B2(new_n860), .ZN(G331));
  NAND2_X1  g531(.A1(new_n945), .A2(new_n948), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  NAND2_X1  g533(.A1(G171), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT110), .B1(new_n535), .B2(new_n538), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(G286), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(G171), .A2(G168), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n867), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n865), .B2(new_n866), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n965), .A2(new_n936), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n927), .B1(new_n965), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n957), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n926), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n936), .A3(new_n966), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n949), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n973), .A3(new_n918), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n969), .A2(new_n973), .A3(new_n976), .A4(new_n918), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n978), .B2(KEYINPUT109), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n980), .B(new_n981), .C1(new_n975), .C2(new_n977), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n979), .A2(new_n982), .ZN(G397));
  XNOR2_X1  g558(.A(new_n772), .B(G2067), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n891), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n479), .A2(G40), .A3(new_n471), .A4(new_n469), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT112), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n989), .A2(new_n692), .A3(new_n724), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT111), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n989), .A2(G1996), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n724), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n992), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n830), .A2(new_n832), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n830), .A2(new_n832), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(G290), .B(G1986), .Z(new_n1001));
  OAI211_X1 g576(.A(new_n997), .B(new_n1000), .C1(new_n989), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n891), .A2(new_n1005), .A3(new_n985), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n985), .B1(new_n498), .B2(new_n502), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n987), .B1(new_n1007), .B2(KEYINPUT50), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n704), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n891), .A2(new_n985), .A3(new_n988), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(G2067), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1013), .A3(KEYINPUT117), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n703), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n1012), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n603), .B1(new_n1018), .B2(KEYINPUT60), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n1020), .B(new_n615), .C1(new_n1014), .C2(new_n1017), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n1019), .A2(new_n1021), .B1(KEYINPUT60), .B2(new_n1018), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT61), .ZN(new_n1023));
  INV_X1    g598(.A(G1956), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1005), .B1(new_n891), .B2(new_n985), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n988), .B1(new_n1007), .B2(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G299), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n563), .B(KEYINPUT57), .C1(new_n567), .C2(new_n569), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n891), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n987), .B1(new_n1007), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT56), .B(G2072), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1027), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1031), .B1(new_n1027), .B2(new_n1036), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1023), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1031), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT61), .A3(new_n1037), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1032), .A2(new_n1034), .A3(new_n692), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1032), .A2(new_n1034), .A3(KEYINPUT118), .A4(new_n692), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT58), .B(G1341), .Z(new_n1051));
  NAND2_X1  g626(.A1(new_n1011), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  AOI211_X1 g628(.A(new_n1046), .B(KEYINPUT59), .C1(new_n1053), .C2(new_n552), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1045), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n552), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT119), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1046), .A3(new_n552), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT59), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1022), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1018), .A2(new_n603), .A3(new_n1038), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(new_n1039), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1006), .A2(new_n1008), .A3(new_n731), .ZN(new_n1064));
  INV_X1    g639(.A(G1966), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1033), .B1(new_n900), .B2(G1384), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n503), .A2(KEYINPUT116), .A3(KEYINPUT45), .A4(new_n985), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1007), .B2(new_n1033), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n988), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1064), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G286), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(KEYINPUT120), .A2(G8), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1075), .B(new_n1076), .C1(new_n1071), .C2(G168), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1070), .A2(new_n1065), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1064), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(G168), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1076), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT51), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1074), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT121), .B(new_n1074), .C1(new_n1077), .C2(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n467), .B1(new_n478), .B2(KEYINPUT122), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(KEYINPUT122), .B2(new_n478), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n472), .A2(G40), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1066), .A2(new_n1088), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT123), .B1(new_n986), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(G2078), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1032), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1092), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1099), .B2(G2078), .ZN(new_n1100));
  INV_X1    g675(.A(G1961), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1009), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(G301), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1096), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1102), .B1(new_n1070), .B2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1108), .A3(KEYINPUT54), .ZN(new_n1109));
  NAND3_X1  g684(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1112));
  OAI21_X1  g687(.A(G8), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1971), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1009), .A2(G2090), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1025), .A2(new_n1026), .A3(G2090), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n1118), .B2(new_n1114), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n586), .A2(new_n587), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G1981), .ZN(new_n1126));
  INV_X1    g701(.A(G1981), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n586), .A2(new_n589), .A3(new_n1127), .A4(new_n590), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT49), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1011), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(new_n1072), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(KEYINPUT49), .A3(new_n1128), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1011), .A2(G288), .A3(G8), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT114), .B1(new_n578), .B2(G1976), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1011), .A2(G8), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT52), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1124), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1109), .A2(new_n1123), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1100), .ZN(new_n1147));
  OAI21_X1  g722(.A(G171), .B1(new_n1107), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1098), .A2(G301), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g727(.A(KEYINPUT124), .B(KEYINPUT54), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1145), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1063), .A2(new_n1087), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1123), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1144), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1073), .A2(G168), .ZN(new_n1158));
  NOR4_X1   g733(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT63), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1116), .A2(new_n1120), .A3(new_n1115), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1160), .B(new_n1135), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT63), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1135), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n579), .A2(new_n1136), .A3(new_n581), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1128), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1133), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1117), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1162), .B(new_n1166), .C1(new_n1167), .C2(new_n1143), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1159), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1155), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1085), .A2(new_n1171), .A3(new_n1086), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1156), .A2(new_n1157), .A3(new_n1148), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1004), .B1(new_n1170), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n997), .A2(new_n999), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n896), .A2(new_n774), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n989), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n997), .A2(new_n1000), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT126), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT48), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n995), .A2(KEYINPUT46), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n995), .A2(KEYINPUT46), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n990), .B1(new_n984), .B2(new_n723), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1192));
  XNOR2_X1  g767(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1181), .A2(new_n1186), .A3(new_n1187), .A4(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1193), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT127), .B1(new_n1195), .B2(new_n1180), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1177), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g773(.A1(G227), .A2(new_n461), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n658), .A2(new_n1200), .ZN(new_n1201));
  NOR3_X1   g775(.A1(new_n697), .A2(new_n698), .A3(new_n1201), .ZN(new_n1202));
  OAI211_X1 g776(.A(new_n978), .B(new_n1202), .C1(new_n920), .C2(new_n919), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


