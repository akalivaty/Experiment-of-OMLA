

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(n534), .B(KEYINPUT0), .ZN(n631) );
  NOR2_X1 U555 ( .A1(G651), .A2(n631), .ZN(n651) );
  NOR2_X2 U556 ( .A1(n598), .A2(n597), .ZN(n1013) );
  BUF_X1 U557 ( .A(n601), .Z(n571) );
  BUF_X1 U558 ( .A(n559), .Z(n560) );
  XNOR2_X1 U559 ( .A(KEYINPUT67), .B(G543), .ZN(n534) );
  XNOR2_X1 U560 ( .A(n777), .B(n776), .ZN(n778) );
  AND2_X1 U561 ( .A1(n784), .A2(n790), .ZN(n785) );
  INV_X1 U562 ( .A(KEYINPUT106), .ZN(n829) );
  AND2_X1 U563 ( .A1(n826), .A2(n521), .ZN(n827) );
  NOR2_X2 U564 ( .A1(n533), .A2(n532), .ZN(G160) );
  OR2_X1 U565 ( .A1(n825), .A2(n824), .ZN(n521) );
  AND2_X1 U566 ( .A1(n828), .A2(n827), .ZN(n522) );
  AND2_X1 U567 ( .A1(n836), .A2(n835), .ZN(n523) );
  XNOR2_X1 U568 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n776) );
  INV_X1 U569 ( .A(KEYINPUT29), .ZN(n764) );
  AND2_X1 U570 ( .A1(n799), .A2(n798), .ZN(n801) );
  NOR2_X2 U571 ( .A1(n730), .A2(n729), .ZN(n766) );
  INV_X1 U572 ( .A(n832), .ZN(n833) );
  NOR2_X1 U573 ( .A1(n834), .A2(n833), .ZN(n836) );
  INV_X1 U574 ( .A(KEYINPUT78), .ZN(n540) );
  NOR2_X1 U575 ( .A1(n526), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U576 ( .A(n540), .B(KEYINPUT5), .ZN(n541) );
  XNOR2_X1 U577 ( .A(n542), .B(n541), .ZN(n550) );
  XNOR2_X1 U578 ( .A(n551), .B(KEYINPUT7), .ZN(G168) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n995) );
  NAND2_X1 U580 ( .A1(G113), .A2(n995), .ZN(n525) );
  INV_X1 U581 ( .A(G2104), .ZN(n526) );
  AND2_X1 U582 ( .A1(n526), .A2(G2105), .ZN(n996) );
  NAND2_X1 U583 ( .A1(G125), .A2(n996), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n525), .A2(n524), .ZN(n533) );
  XNOR2_X2 U585 ( .A(n527), .B(KEYINPUT66), .ZN(n999) );
  NAND2_X1 U586 ( .A1(n999), .A2(G101), .ZN(n528) );
  XOR2_X1 U587 ( .A(KEYINPUT23), .B(n528), .Z(n531) );
  NOR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X1 U589 ( .A(KEYINPUT17), .B(n529), .Z(n559) );
  NAND2_X1 U590 ( .A1(n559), .A2(G137), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U592 ( .A(G651), .ZN(n543) );
  OR2_X1 U593 ( .A1(n543), .A2(n631), .ZN(n535) );
  XOR2_X1 U594 ( .A(KEYINPUT68), .B(n535), .Z(n601) );
  NAND2_X1 U595 ( .A1(G76), .A2(n601), .ZN(n536) );
  XNOR2_X1 U596 ( .A(KEYINPUT77), .B(n536), .ZN(n539) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U598 ( .A1(n650), .A2(G89), .ZN(n537) );
  XOR2_X1 U599 ( .A(n537), .B(KEYINPUT4), .Z(n538) );
  NOR2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n542) );
  NOR2_X1 U601 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n544), .Z(n657) );
  NAND2_X1 U603 ( .A1(n657), .A2(G63), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT79), .B(n545), .Z(n547) );
  NAND2_X1 U605 ( .A1(n651), .A2(G51), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n548), .Z(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U609 ( .A1(G138), .A2(n559), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G102), .A2(n999), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U612 ( .A(n554), .B(KEYINPUT86), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G114), .A2(n995), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G126), .A2(n996), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(G164) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U618 ( .A1(G135), .A2(n560), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G111), .A2(n995), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n996), .A2(G123), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT18), .B(n563), .Z(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U624 ( .A1(G99), .A2(n999), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n1005) );
  XNOR2_X1 U626 ( .A(G2096), .B(n1005), .ZN(n568) );
  OR2_X1 U627 ( .A1(G2100), .A2(n568), .ZN(G156) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  NAND2_X1 U631 ( .A1(G64), .A2(n657), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G52), .A2(n651), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n576) );
  NAND2_X1 U634 ( .A1(G90), .A2(n650), .ZN(n573) );
  NAND2_X1 U635 ( .A1(G77), .A2(n571), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT9), .B(n574), .Z(n575) );
  NOR2_X1 U638 ( .A1(n576), .A2(n575), .ZN(G171) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G65), .A2(n657), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G91), .A2(n650), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n651), .A2(G53), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT70), .B(n579), .Z(n580) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G78), .A2(n571), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(G299) );
  XOR2_X1 U648 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n587) );
  XOR2_X1 U649 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n585) );
  NAND2_X1 U650 ( .A1(G7), .A2(G661), .ZN(n584) );
  XOR2_X1 U651 ( .A(n585), .B(n584), .Z(n1035) );
  NAND2_X1 U652 ( .A1(G567), .A2(n1035), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(G234) );
  NAND2_X1 U654 ( .A1(G56), .A2(n657), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n588), .B(KEYINPUT14), .ZN(n595) );
  NAND2_X1 U656 ( .A1(n650), .A2(G81), .ZN(n589) );
  XNOR2_X1 U657 ( .A(n589), .B(KEYINPUT12), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G68), .A2(n601), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n593) );
  XOR2_X1 U660 ( .A(KEYINPUT13), .B(KEYINPUT73), .Z(n592) );
  XNOR2_X1 U661 ( .A(n593), .B(n592), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n651), .A2(G43), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT74), .B(n596), .Z(n597) );
  NAND2_X1 U665 ( .A1(n1013), .A2(G860), .ZN(G153) );
  INV_X1 U666 ( .A(G171), .ZN(G301) );
  NAND2_X1 U667 ( .A1(n651), .A2(G54), .ZN(n606) );
  NAND2_X1 U668 ( .A1(G66), .A2(n657), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G92), .A2(n650), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U671 ( .A1(G79), .A2(n601), .ZN(n602) );
  XNOR2_X1 U672 ( .A(KEYINPUT75), .B(n602), .ZN(n603) );
  NOR2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U675 ( .A(KEYINPUT15), .B(n607), .ZN(n608) );
  INV_X1 U676 ( .A(n608), .ZN(n755) );
  INV_X1 U677 ( .A(G868), .ZN(n667) );
  NAND2_X1 U678 ( .A1(n755), .A2(n667), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n609), .B(KEYINPUT76), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G868), .A2(G301), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(G284) );
  NOR2_X1 U682 ( .A1(G286), .A2(n667), .ZN(n613) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U684 ( .A1(n613), .A2(n612), .ZN(G297) );
  INV_X1 U685 ( .A(G860), .ZN(n621) );
  NAND2_X1 U686 ( .A1(n621), .A2(G559), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n614), .A2(n608), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U689 ( .A1(n1013), .A2(n667), .ZN(n616) );
  XOR2_X1 U690 ( .A(KEYINPUT80), .B(n616), .Z(n619) );
  NAND2_X1 U691 ( .A1(G868), .A2(n608), .ZN(n617) );
  NOR2_X1 U692 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U694 ( .A1(G559), .A2(n608), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n620), .B(n1013), .ZN(n665) );
  NAND2_X1 U696 ( .A1(n621), .A2(n665), .ZN(n629) );
  NAND2_X1 U697 ( .A1(G67), .A2(n657), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G93), .A2(n650), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G80), .A2(n571), .ZN(n624) );
  XNOR2_X1 U701 ( .A(KEYINPUT81), .B(n624), .ZN(n625) );
  NOR2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n651), .A2(G55), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n668) );
  XNOR2_X1 U705 ( .A(n629), .B(n668), .ZN(G145) );
  NAND2_X1 U706 ( .A1(G49), .A2(n651), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n630), .B(KEYINPUT82), .ZN(n636) );
  NAND2_X1 U708 ( .A1(G87), .A2(n631), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n657), .A2(n634), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G88), .A2(n650), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G75), .A2(n571), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G62), .A2(n657), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G50), .A2(n651), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U719 ( .A1(n642), .A2(n641), .ZN(G166) );
  INV_X1 U720 ( .A(G166), .ZN(G303) );
  NAND2_X1 U721 ( .A1(n650), .A2(G85), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n657), .A2(G60), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n651), .A2(G47), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G72), .A2(n571), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(KEYINPUT69), .B(n649), .ZN(G290) );
  NAND2_X1 U729 ( .A1(G86), .A2(n650), .ZN(n653) );
  NAND2_X1 U730 ( .A1(G48), .A2(n651), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n571), .A2(G73), .ZN(n654) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U734 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n657), .A2(G61), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(G305) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(G288), .ZN(n664) );
  XOR2_X1 U738 ( .A(G290), .B(G305), .Z(n660) );
  XNOR2_X1 U739 ( .A(n668), .B(n660), .ZN(n661) );
  XOR2_X1 U740 ( .A(G303), .B(n661), .Z(n662) );
  XNOR2_X1 U741 ( .A(n662), .B(G299), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n664), .B(n663), .ZN(n1012) );
  XNOR2_X1 U743 ( .A(n665), .B(n1012), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n666), .A2(G868), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XNOR2_X1 U748 ( .A(n671), .B(KEYINPUT20), .ZN(n672) );
  XNOR2_X1 U749 ( .A(n672), .B(KEYINPUT83), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n673), .A2(G2090), .ZN(n674) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U752 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U756 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U757 ( .A1(G96), .A2(n678), .ZN(n963) );
  NAND2_X1 U758 ( .A1(G2106), .A2(n963), .ZN(n682) );
  NAND2_X1 U759 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U760 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U761 ( .A1(G108), .A2(n680), .ZN(n964) );
  NAND2_X1 U762 ( .A1(G567), .A2(n964), .ZN(n681) );
  NAND2_X1 U763 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U764 ( .A(KEYINPUT84), .B(n683), .ZN(n965) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U766 ( .A1(n965), .A2(n684), .ZN(n843) );
  NAND2_X1 U767 ( .A1(n843), .A2(G36), .ZN(n685) );
  XOR2_X1 U768 ( .A(KEYINPUT85), .B(n685), .Z(G176) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n728) );
  NAND2_X1 U770 ( .A1(G160), .A2(G40), .ZN(n729) );
  NOR2_X1 U771 ( .A1(n728), .A2(n729), .ZN(n830) );
  NAND2_X1 U772 ( .A1(G105), .A2(n999), .ZN(n688) );
  XOR2_X1 U773 ( .A(KEYINPUT38), .B(KEYINPUT92), .Z(n686) );
  XNOR2_X1 U774 ( .A(KEYINPUT91), .B(n686), .ZN(n687) );
  XNOR2_X1 U775 ( .A(n688), .B(n687), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G117), .A2(n995), .ZN(n690) );
  NAND2_X1 U777 ( .A1(G129), .A2(n996), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U779 ( .A1(G141), .A2(n560), .ZN(n691) );
  XNOR2_X1 U780 ( .A(KEYINPUT93), .B(n691), .ZN(n692) );
  NOR2_X1 U781 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n994) );
  NOR2_X1 U783 ( .A1(G1996), .A2(n994), .ZN(n696) );
  XOR2_X1 U784 ( .A(KEYINPUT107), .B(n696), .Z(n873) );
  NAND2_X1 U785 ( .A1(G131), .A2(n560), .ZN(n698) );
  NAND2_X1 U786 ( .A1(G107), .A2(n995), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n996), .A2(G119), .ZN(n700) );
  NAND2_X1 U789 ( .A1(G95), .A2(n999), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n1008) );
  NAND2_X1 U792 ( .A1(G1991), .A2(n1008), .ZN(n704) );
  NAND2_X1 U793 ( .A1(G1996), .A2(n994), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n879) );
  NAND2_X1 U795 ( .A1(n879), .A2(n830), .ZN(n705) );
  XNOR2_X1 U796 ( .A(KEYINPUT94), .B(n705), .ZN(n835) );
  INV_X1 U797 ( .A(n835), .ZN(n709) );
  NOR2_X1 U798 ( .A1(G1986), .A2(G290), .ZN(n707) );
  NOR2_X1 U799 ( .A1(G1991), .A2(n1008), .ZN(n706) );
  XNOR2_X1 U800 ( .A(KEYINPUT108), .B(n706), .ZN(n876) );
  NOR2_X1 U801 ( .A1(n707), .A2(n876), .ZN(n708) );
  NOR2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n873), .A2(n710), .ZN(n711) );
  XNOR2_X1 U804 ( .A(n711), .B(KEYINPUT39), .ZN(n724) );
  XNOR2_X1 U805 ( .A(G2067), .B(KEYINPUT37), .ZN(n712) );
  XNOR2_X1 U806 ( .A(n712), .B(KEYINPUT88), .ZN(n725) );
  NAND2_X1 U807 ( .A1(n560), .A2(G140), .ZN(n713) );
  XOR2_X1 U808 ( .A(KEYINPUT89), .B(n713), .Z(n715) );
  NAND2_X1 U809 ( .A1(G104), .A2(n999), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n717) );
  XNOR2_X1 U811 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n716) );
  XNOR2_X1 U812 ( .A(n717), .B(n716), .ZN(n722) );
  NAND2_X1 U813 ( .A1(G116), .A2(n995), .ZN(n719) );
  NAND2_X1 U814 ( .A1(G128), .A2(n996), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U816 ( .A(KEYINPUT35), .B(n720), .Z(n721) );
  NOR2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U818 ( .A(KEYINPUT36), .B(n723), .ZN(n988) );
  NOR2_X1 U819 ( .A1(n725), .A2(n988), .ZN(n883) );
  NAND2_X1 U820 ( .A1(n830), .A2(n883), .ZN(n832) );
  NAND2_X1 U821 ( .A1(n724), .A2(n832), .ZN(n726) );
  NAND2_X1 U822 ( .A1(n725), .A2(n988), .ZN(n899) );
  NAND2_X1 U823 ( .A1(n726), .A2(n899), .ZN(n727) );
  NAND2_X1 U824 ( .A1(n830), .A2(n727), .ZN(n839) );
  INV_X1 U825 ( .A(n728), .ZN(n730) );
  INV_X1 U826 ( .A(n766), .ZN(n743) );
  NAND2_X1 U827 ( .A1(G8), .A2(n743), .ZN(n825) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n825), .ZN(n774) );
  INV_X1 U829 ( .A(n774), .ZN(n784) );
  INV_X1 U830 ( .A(KEYINPUT65), .ZN(n741) );
  XOR2_X1 U831 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n734) );
  XOR2_X1 U832 ( .A(G1996), .B(n734), .Z(n731) );
  NOR2_X1 U833 ( .A1(n743), .A2(n731), .ZN(n732) );
  INV_X1 U834 ( .A(KEYINPUT95), .ZN(n733) );
  NAND2_X1 U835 ( .A1(n732), .A2(n733), .ZN(n738) );
  XOR2_X1 U836 ( .A(n733), .B(G1341), .Z(n736) );
  NOR2_X1 U837 ( .A1(n766), .A2(n734), .ZN(n735) );
  NAND2_X1 U838 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U839 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U840 ( .A1(n739), .A2(n1013), .ZN(n740) );
  XNOR2_X1 U841 ( .A(n741), .B(n740), .ZN(n754) );
  NOR2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n742) );
  XNOR2_X1 U843 ( .A(n742), .B(KEYINPUT96), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n766), .A2(G1348), .ZN(n745) );
  BUF_X1 U845 ( .A(n743), .Z(n773) );
  NOR2_X1 U846 ( .A1(G2067), .A2(n773), .ZN(n744) );
  NOR2_X1 U847 ( .A1(n745), .A2(n744), .ZN(n750) );
  NAND2_X1 U848 ( .A1(n766), .A2(G2072), .ZN(n746) );
  XOR2_X1 U849 ( .A(KEYINPUT27), .B(n746), .Z(n748) );
  NAND2_X1 U850 ( .A1(G1956), .A2(n773), .ZN(n747) );
  NAND2_X1 U851 ( .A1(n748), .A2(n747), .ZN(n758) );
  NOR2_X1 U852 ( .A1(n758), .A2(G299), .ZN(n749) );
  XNOR2_X1 U853 ( .A(n749), .B(KEYINPUT97), .ZN(n753) );
  NAND2_X1 U854 ( .A1(n750), .A2(n753), .ZN(n751) );
  OR2_X1 U855 ( .A1(n752), .A2(n751), .ZN(n763) );
  INV_X1 U856 ( .A(n753), .ZN(n757) );
  NAND2_X1 U857 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U858 ( .A1(n757), .A2(n756), .ZN(n761) );
  NAND2_X1 U859 ( .A1(G299), .A2(n758), .ZN(n759) );
  XOR2_X1 U860 ( .A(n759), .B(KEYINPUT28), .Z(n760) );
  NOR2_X1 U861 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U862 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U863 ( .A(n765), .B(n764), .ZN(n770) );
  NAND2_X1 U864 ( .A1(G1961), .A2(n773), .ZN(n768) );
  XOR2_X1 U865 ( .A(G2078), .B(KEYINPUT25), .Z(n855) );
  NAND2_X1 U866 ( .A1(n766), .A2(n855), .ZN(n767) );
  NAND2_X1 U867 ( .A1(n768), .A2(n767), .ZN(n771) );
  OR2_X1 U868 ( .A1(G301), .A2(n771), .ZN(n769) );
  NAND2_X1 U869 ( .A1(n770), .A2(n769), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G301), .A2(n771), .ZN(n772) );
  XNOR2_X1 U871 ( .A(n772), .B(KEYINPUT99), .ZN(n780) );
  NOR2_X1 U872 ( .A1(G2084), .A2(n773), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n786), .A2(n774), .ZN(n775) );
  NAND2_X1 U874 ( .A1(n775), .A2(G8), .ZN(n777) );
  NOR2_X1 U875 ( .A1(n778), .A2(G168), .ZN(n779) );
  NOR2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U877 ( .A(KEYINPUT31), .B(n781), .Z(n782) );
  NAND2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n790) );
  XNOR2_X1 U879 ( .A(n785), .B(KEYINPUT100), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n786), .A2(G8), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n803) );
  AND2_X1 U882 ( .A1(G286), .A2(G8), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n799) );
  INV_X1 U884 ( .A(G8), .ZN(n797) );
  NOR2_X1 U885 ( .A1(G1971), .A2(n825), .ZN(n791) );
  XOR2_X1 U886 ( .A(KEYINPUT101), .B(n791), .Z(n793) );
  NOR2_X1 U887 ( .A1(G2090), .A2(n773), .ZN(n792) );
  NOR2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U889 ( .A(n794), .B(KEYINPUT102), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n795), .A2(G303), .ZN(n796) );
  OR2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U892 ( .A(KEYINPUT103), .B(KEYINPUT32), .Z(n800) );
  XNOR2_X1 U893 ( .A(n801), .B(n800), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n820) );
  NOR2_X1 U895 ( .A1(G1976), .A2(G288), .ZN(n810) );
  NOR2_X1 U896 ( .A1(G1971), .A2(G303), .ZN(n804) );
  NOR2_X1 U897 ( .A1(n810), .A2(n804), .ZN(n916) );
  NAND2_X1 U898 ( .A1(n820), .A2(n916), .ZN(n805) );
  NAND2_X1 U899 ( .A1(G1976), .A2(G288), .ZN(n912) );
  NAND2_X1 U900 ( .A1(n805), .A2(n912), .ZN(n807) );
  INV_X1 U901 ( .A(KEYINPUT104), .ZN(n809) );
  OR2_X1 U902 ( .A1(n825), .A2(n809), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U904 ( .A1(KEYINPUT33), .A2(n808), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n809), .A2(n810), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n810), .A2(KEYINPUT33), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n811), .A2(KEYINPUT104), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n825), .A2(n814), .ZN(n815) );
  NOR2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U911 ( .A(G1981), .B(G305), .Z(n923) );
  NAND2_X1 U912 ( .A1(n817), .A2(n923), .ZN(n828) );
  NAND2_X1 U913 ( .A1(G8), .A2(G166), .ZN(n818) );
  NOR2_X1 U914 ( .A1(G2090), .A2(n818), .ZN(n819) );
  XNOR2_X1 U915 ( .A(n819), .B(KEYINPUT105), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n822), .A2(n825), .ZN(n826) );
  NOR2_X1 U918 ( .A1(G1981), .A2(G305), .ZN(n823) );
  XOR2_X1 U919 ( .A(n823), .B(KEYINPUT24), .Z(n824) );
  XNOR2_X1 U920 ( .A(n522), .B(n829), .ZN(n837) );
  XNOR2_X1 U921 ( .A(G1986), .B(G290), .ZN(n918) );
  NAND2_X1 U922 ( .A1(n830), .A2(n918), .ZN(n831) );
  XNOR2_X1 U923 ( .A(KEYINPUT87), .B(n831), .ZN(n834) );
  NAND2_X1 U924 ( .A1(n837), .A2(n523), .ZN(n838) );
  NAND2_X1 U925 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(n840), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n1035), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U929 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U931 ( .A1(n843), .A2(n842), .ZN(G188) );
  NAND2_X1 U933 ( .A1(G124), .A2(n996), .ZN(n844) );
  XNOR2_X1 U934 ( .A(n844), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U935 ( .A1(n995), .A2(G112), .ZN(n845) );
  NAND2_X1 U936 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U937 ( .A1(G136), .A2(n560), .ZN(n848) );
  NAND2_X1 U938 ( .A1(G100), .A2(n999), .ZN(n847) );
  NAND2_X1 U939 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U940 ( .A1(n850), .A2(n849), .ZN(G162) );
  XOR2_X1 U941 ( .A(G2072), .B(G33), .Z(n851) );
  NAND2_X1 U942 ( .A1(n851), .A2(G28), .ZN(n853) );
  XNOR2_X1 U943 ( .A(G26), .B(G2067), .ZN(n852) );
  NOR2_X1 U944 ( .A1(n853), .A2(n852), .ZN(n862) );
  XNOR2_X1 U945 ( .A(G1991), .B(G25), .ZN(n854) );
  XNOR2_X1 U946 ( .A(n854), .B(KEYINPUT118), .ZN(n860) );
  XNOR2_X1 U947 ( .A(G1996), .B(G32), .ZN(n857) );
  XNOR2_X1 U948 ( .A(n855), .B(G27), .ZN(n856) );
  NOR2_X1 U949 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U950 ( .A(KEYINPUT119), .B(n858), .ZN(n859) );
  NOR2_X1 U951 ( .A1(n860), .A2(n859), .ZN(n861) );
  NAND2_X1 U952 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U953 ( .A(n863), .B(KEYINPUT53), .ZN(n866) );
  XOR2_X1 U954 ( .A(G2084), .B(G34), .Z(n864) );
  XNOR2_X1 U955 ( .A(KEYINPUT54), .B(n864), .ZN(n865) );
  NAND2_X1 U956 ( .A1(n866), .A2(n865), .ZN(n868) );
  XNOR2_X1 U957 ( .A(G35), .B(G2090), .ZN(n867) );
  NOR2_X1 U958 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U959 ( .A(KEYINPUT55), .B(n869), .Z(n871) );
  INV_X1 U960 ( .A(G29), .ZN(n905) );
  XOR2_X1 U961 ( .A(n905), .B(KEYINPUT120), .Z(n870) );
  NOR2_X1 U962 ( .A1(n871), .A2(n870), .ZN(n907) );
  XOR2_X1 U963 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n902) );
  XOR2_X1 U964 ( .A(G2090), .B(G162), .Z(n872) );
  NOR2_X1 U965 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U966 ( .A(KEYINPUT51), .B(n874), .Z(n881) );
  XOR2_X1 U967 ( .A(G160), .B(G2084), .Z(n875) );
  NOR2_X1 U968 ( .A1(n876), .A2(n875), .ZN(n877) );
  NAND2_X1 U969 ( .A1(n877), .A2(n1005), .ZN(n878) );
  NOR2_X1 U970 ( .A1(n879), .A2(n878), .ZN(n880) );
  NAND2_X1 U971 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U972 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U973 ( .A(KEYINPUT116), .B(n884), .Z(n898) );
  XNOR2_X1 U974 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n888) );
  NAND2_X1 U975 ( .A1(G115), .A2(n995), .ZN(n886) );
  NAND2_X1 U976 ( .A1(G127), .A2(n996), .ZN(n885) );
  NAND2_X1 U977 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U978 ( .A(n888), .B(n887), .ZN(n893) );
  NAND2_X1 U979 ( .A1(n560), .A2(G139), .ZN(n889) );
  XNOR2_X1 U980 ( .A(n889), .B(KEYINPUT112), .ZN(n891) );
  NAND2_X1 U981 ( .A1(G103), .A2(n999), .ZN(n890) );
  NAND2_X1 U982 ( .A1(n891), .A2(n890), .ZN(n892) );
  NOR2_X1 U983 ( .A1(n893), .A2(n892), .ZN(n987) );
  XOR2_X1 U984 ( .A(G2072), .B(n987), .Z(n895) );
  XOR2_X1 U985 ( .A(G164), .B(G2078), .Z(n894) );
  NOR2_X1 U986 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U987 ( .A(KEYINPUT50), .B(n896), .Z(n897) );
  NOR2_X1 U988 ( .A1(n898), .A2(n897), .ZN(n900) );
  NAND2_X1 U989 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U990 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U991 ( .A1(KEYINPUT55), .A2(n903), .ZN(n904) );
  NOR2_X1 U992 ( .A1(n905), .A2(n904), .ZN(n906) );
  NOR2_X1 U993 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U994 ( .A1(G11), .A2(n908), .ZN(n961) );
  INV_X1 U995 ( .A(G16), .ZN(n956) );
  XOR2_X1 U996 ( .A(n956), .B(KEYINPUT56), .Z(n931) );
  XOR2_X1 U997 ( .A(n1013), .B(G1341), .Z(n910) );
  XNOR2_X1 U998 ( .A(G301), .B(G1961), .ZN(n909) );
  NOR2_X1 U999 ( .A1(n910), .A2(n909), .ZN(n921) );
  NAND2_X1 U1000 ( .A1(G1971), .A2(G303), .ZN(n911) );
  NAND2_X1 U1001 ( .A1(n912), .A2(n911), .ZN(n914) );
  XNOR2_X1 U1002 ( .A(G1956), .B(G299), .ZN(n913) );
  NOR2_X1 U1003 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1004 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1005 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1006 ( .A(n919), .B(KEYINPUT122), .ZN(n920) );
  NAND2_X1 U1007 ( .A1(n921), .A2(n920), .ZN(n927) );
  XOR2_X1 U1008 ( .A(G1966), .B(G168), .Z(n922) );
  XNOR2_X1 U1009 ( .A(KEYINPUT121), .B(n922), .ZN(n924) );
  NAND2_X1 U1010 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1011 ( .A(KEYINPUT57), .B(n925), .Z(n926) );
  NOR2_X1 U1012 ( .A1(n927), .A2(n926), .ZN(n929) );
  XNOR2_X1 U1013 ( .A(G1348), .B(n608), .ZN(n928) );
  NAND2_X1 U1014 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1015 ( .A1(n931), .A2(n930), .ZN(n958) );
  XNOR2_X1 U1016 ( .A(G1348), .B(KEYINPUT59), .ZN(n932) );
  XNOR2_X1 U1017 ( .A(n932), .B(G4), .ZN(n936) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G19), .ZN(n934) );
  XNOR2_X1 U1019 ( .A(G6), .B(G1981), .ZN(n933) );
  NOR2_X1 U1020 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1021 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1022 ( .A(KEYINPUT123), .B(G1956), .Z(n937) );
  XNOR2_X1 U1023 ( .A(G20), .B(n937), .ZN(n938) );
  NOR2_X1 U1024 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1025 ( .A(KEYINPUT60), .B(n940), .ZN(n941) );
  XNOR2_X1 U1026 ( .A(n941), .B(KEYINPUT124), .ZN(n945) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G21), .ZN(n943) );
  XNOR2_X1 U1028 ( .A(G5), .B(G1961), .ZN(n942) );
  NOR2_X1 U1029 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1030 ( .A1(n945), .A2(n944), .ZN(n953) );
  XNOR2_X1 U1031 ( .A(G1986), .B(G24), .ZN(n950) );
  XNOR2_X1 U1032 ( .A(G1971), .B(G22), .ZN(n947) );
  XNOR2_X1 U1033 ( .A(G23), .B(G1976), .ZN(n946) );
  NOR2_X1 U1034 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1035 ( .A(KEYINPUT125), .B(n948), .ZN(n949) );
  NOR2_X1 U1036 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1037 ( .A(KEYINPUT58), .B(n951), .Z(n952) );
  NOR2_X1 U1038 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1039 ( .A(KEYINPUT61), .B(n954), .ZN(n955) );
  NAND2_X1 U1040 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1041 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1042 ( .A(n959), .B(KEYINPUT126), .ZN(n960) );
  NOR2_X1 U1043 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1044 ( .A(KEYINPUT62), .B(n962), .ZN(G311) );
  XNOR2_X1 U1045 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1046 ( .A(G120), .ZN(G236) );
  INV_X1 U1047 ( .A(G96), .ZN(G221) );
  INV_X1 U1048 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1049 ( .A1(n964), .A2(n963), .ZN(G325) );
  INV_X1 U1050 ( .A(G325), .ZN(G261) );
  INV_X1 U1051 ( .A(n965), .ZN(G319) );
  XOR2_X1 U1052 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n967) );
  XNOR2_X1 U1053 ( .A(G2072), .B(G2090), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(n967), .B(n966), .ZN(n971) );
  XOR2_X1 U1055 ( .A(KEYINPUT111), .B(G2678), .Z(n969) );
  XNOR2_X1 U1056 ( .A(G2067), .B(KEYINPUT43), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1058 ( .A(n971), .B(n970), .Z(n973) );
  XNOR2_X1 U1059 ( .A(G2096), .B(G2100), .ZN(n972) );
  XNOR2_X1 U1060 ( .A(n973), .B(n972), .ZN(n975) );
  XOR2_X1 U1061 ( .A(G2084), .B(G2078), .Z(n974) );
  XNOR2_X1 U1062 ( .A(n975), .B(n974), .ZN(G227) );
  XOR2_X1 U1063 ( .A(KEYINPUT41), .B(G1971), .Z(n977) );
  XNOR2_X1 U1064 ( .A(G1986), .B(G1961), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(n977), .B(n976), .ZN(n978) );
  XOR2_X1 U1066 ( .A(n978), .B(G1981), .Z(n980) );
  XNOR2_X1 U1067 ( .A(G1991), .B(G1966), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(n980), .B(n979), .ZN(n984) );
  XOR2_X1 U1069 ( .A(G2474), .B(G1976), .Z(n982) );
  XNOR2_X1 U1070 ( .A(G1996), .B(G1956), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(n982), .B(n981), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(n984), .B(n983), .ZN(G229) );
  XOR2_X1 U1073 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n986) );
  XNOR2_X1 U1074 ( .A(G162), .B(KEYINPUT46), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n986), .B(n985), .ZN(n992) );
  XNOR2_X1 U1076 ( .A(n988), .B(n987), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(G164), .B(G160), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n990), .B(n989), .ZN(n991) );
  XOR2_X1 U1079 ( .A(n992), .B(n991), .Z(n993) );
  XNOR2_X1 U1080 ( .A(n994), .B(n993), .ZN(n1010) );
  NAND2_X1 U1081 ( .A1(G118), .A2(n995), .ZN(n998) );
  NAND2_X1 U1082 ( .A1(G130), .A2(n996), .ZN(n997) );
  NAND2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n1004) );
  NAND2_X1 U1084 ( .A1(G142), .A2(n560), .ZN(n1001) );
  NAND2_X1 U1085 ( .A1(G106), .A2(n999), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1087 ( .A(n1002), .B(KEYINPUT45), .Z(n1003) );
  NOR2_X1 U1088 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(n1008), .B(n1007), .Z(n1009) );
  XNOR2_X1 U1091 ( .A(n1010), .B(n1009), .ZN(n1011) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1011), .ZN(G395) );
  XOR2_X1 U1093 ( .A(KEYINPUT115), .B(n1012), .Z(n1015) );
  XNOR2_X1 U1094 ( .A(n1013), .B(G286), .ZN(n1014) );
  XNOR2_X1 U1095 ( .A(n1015), .B(n1014), .ZN(n1017) );
  XOR2_X1 U1096 ( .A(n608), .B(G171), .Z(n1016) );
  XNOR2_X1 U1097 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NOR2_X1 U1098 ( .A1(G37), .A2(n1018), .ZN(G397) );
  XOR2_X1 U1099 ( .A(G2438), .B(G2454), .Z(n1020) );
  XNOR2_X1 U1100 ( .A(G1341), .B(G2430), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(n1020), .B(n1019), .ZN(n1027) );
  XOR2_X1 U1102 ( .A(G2443), .B(G2427), .Z(n1022) );
  XNOR2_X1 U1103 ( .A(G1348), .B(KEYINPUT109), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(n1022), .B(n1021), .ZN(n1023) );
  XOR2_X1 U1105 ( .A(n1023), .B(G2435), .Z(n1025) );
  XNOR2_X1 U1106 ( .A(G2451), .B(G2446), .ZN(n1024) );
  XNOR2_X1 U1107 ( .A(n1025), .B(n1024), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(n1027), .B(n1026), .ZN(n1028) );
  NAND2_X1 U1109 ( .A1(n1028), .A2(G14), .ZN(n1034) );
  NAND2_X1 U1110 ( .A1(n1034), .A2(G319), .ZN(n1031) );
  NOR2_X1 U1111 ( .A1(G227), .A2(G229), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(KEYINPUT49), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  NOR2_X1 U1114 ( .A1(G395), .A2(G397), .ZN(n1032) );
  NAND2_X1 U1115 ( .A1(n1033), .A2(n1032), .ZN(G225) );
  INV_X1 U1116 ( .A(G225), .ZN(G308) );
  INV_X1 U1117 ( .A(G108), .ZN(G238) );
  INV_X1 U1118 ( .A(n1034), .ZN(G401) );
  INV_X1 U1119 ( .A(n1035), .ZN(G223) );
endmodule

