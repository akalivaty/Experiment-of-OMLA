//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT65), .Z(G220));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT68), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G236), .A3(G237), .A4(G235), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n476), .B2(new_n470), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n473), .B1(new_n477), .B2(new_n481), .ZN(G160));
  AND2_X1   g057(.A1(new_n475), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  INV_X1    g059(.A(new_n471), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(KEYINPUT71), .A3(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n471), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n484), .A2(new_n486), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G138), .B1(new_n494), .B2(KEYINPUT73), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n471), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n470), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT72), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n502), .A2(new_n504), .A3(new_n505), .A4(G2104), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n475), .A2(G126), .A3(G2105), .ZN(new_n508));
  INV_X1    g083(.A(G138), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT4), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n475), .A2(new_n511), .A3(new_n470), .A4(new_n495), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n498), .A2(new_n507), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n519), .A2(G62), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT75), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n521), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n526), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT6), .B(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT76), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n534), .A2(new_n536), .A3(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  NAND2_X1  g113(.A1(G63), .A2(G651), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT77), .B(G89), .Z(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n540), .B2(new_n525), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n519), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n538), .A2(new_n542), .A3(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(new_n537), .A2(G52), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n521), .ZN(new_n548));
  INV_X1    g123(.A(new_n518), .ZN(new_n549));
  AOI21_X1  g124(.A(G543), .B1(KEYINPUT74), .B2(KEYINPUT5), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n525), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G90), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n546), .A2(new_n548), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n521), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT78), .Z(new_n558));
  AOI22_X1  g133(.A1(new_n537), .A2(G43), .B1(G81), .B2(new_n552), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  NAND3_X1  g141(.A1(new_n537), .A2(KEYINPUT9), .A3(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n551), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(new_n552), .B2(G91), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n534), .A2(new_n536), .A3(G543), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n567), .A2(new_n571), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  NAND2_X1  g152(.A1(new_n552), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n573), .ZN(G288));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n517), .B2(new_n518), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n517), .B2(new_n518), .ZN(new_n588));
  NAND2_X1  g163(.A1(G48), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n535), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n586), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n552), .A2(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n593), .B1(new_n521), .B2(new_n594), .C1(new_n595), .C2(new_n573), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n552), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  NAND2_X1  g174(.A1(new_n537), .A2(G54), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n519), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n521), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n601), .B1(new_n600), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n599), .B(KEYINPUT80), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n597), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n597), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n622), .B(new_n623), .C1(G868), .C2(new_n560), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n485), .A2(G135), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n470), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G123), .B2(new_n483), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT82), .Z(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT83), .B(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n475), .A2(new_n465), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT15), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2435), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2435), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n651), .A3(new_n647), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2100), .Z(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  AOI21_X1  g246(.A(KEYINPUT18), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  INV_X1    g256(.A(new_n678), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n675), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n675), .A2(KEYINPUT86), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  INV_X1    g264(.A(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n688), .B(new_n693), .ZN(G229));
  NAND3_X1  g269(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT25), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n485), .A2(G139), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n696), .B(new_n697), .C1(new_n470), .C2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G29), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G29), .B2(G33), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G2072), .ZN(new_n705));
  INV_X1    g280(.A(G2072), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n706), .C1(G29), .C2(G33), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G4), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n611), .B2(new_n708), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n705), .A2(new_n707), .B1(G1348), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G27), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G164), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G2078), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(KEYINPUT30), .A2(G28), .ZN(new_n717));
  NOR2_X1   g292(.A1(KEYINPUT30), .A2(G28), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(G171), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G5), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n708), .A2(KEYINPUT23), .A3(G20), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n725));
  INV_X1    g300(.A(G20), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G16), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n724), .B(new_n727), .C1(new_n615), .C2(new_n708), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1956), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n712), .A2(G35), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G162), .B2(new_n712), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT29), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n723), .B(new_n729), .C1(G2090), .C2(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n711), .A2(new_n716), .A3(new_n719), .A4(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G11), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT31), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT28), .ZN(new_n737));
  INV_X1    g312(.A(G26), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G29), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n483), .A2(G128), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n485), .A2(G140), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n470), .A2(G116), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(G29), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n739), .B1(new_n746), .B2(new_n737), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n721), .A2(new_n722), .B1(G2067), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n631), .A2(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(G168), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G16), .B2(G21), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(KEYINPUT31), .B2(new_n735), .ZN(new_n753));
  AND4_X1   g328(.A1(new_n736), .A2(new_n748), .A3(new_n749), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT96), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n747), .A2(G2067), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n712), .B1(new_n758), .B2(G34), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT92), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(G34), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(KEYINPUT92), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G160), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n712), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT93), .B(G2084), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n754), .A2(new_n756), .A3(new_n757), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n560), .A2(G16), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G16), .B2(G19), .ZN(new_n770));
  INV_X1    g345(.A(G1341), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(KEYINPUT95), .B1(G29), .B2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n465), .A2(G105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n483), .A2(G129), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n485), .A2(G141), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(new_n712), .ZN(new_n782));
  MUX2_X1   g357(.A(new_n774), .B(KEYINPUT95), .S(new_n782), .Z(new_n783));
  XOR2_X1   g358(.A(KEYINPUT27), .B(G1996), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n785), .B1(G2090), .B2(new_n732), .C1(new_n770), .C2(new_n771), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n734), .A2(new_n768), .A3(new_n773), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n710), .A2(G1348), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(KEYINPUT97), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n787), .A2(KEYINPUT97), .A3(new_n789), .ZN(new_n792));
  MUX2_X1   g367(.A(G23), .B(G288), .S(G16), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT33), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1976), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n708), .A2(G6), .ZN(new_n796));
  INV_X1    g371(.A(G305), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n708), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G22), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G303), .B2(G16), .ZN(new_n803));
  MUX2_X1   g378(.A(new_n802), .B(new_n803), .S(KEYINPUT88), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1971), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n795), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n807));
  MUX2_X1   g382(.A(G24), .B(G290), .S(G16), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(new_n692), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n483), .A2(G119), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n485), .A2(G131), .ZN(new_n811));
  OR2_X1    g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G29), .ZN(new_n815));
  INV_X1    g390(.A(G25), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT87), .B1(new_n816), .B2(G29), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n816), .A2(KEYINPUT87), .A3(G29), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT35), .B(G1991), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n809), .B(new_n822), .C1(new_n806), .C2(KEYINPUT34), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT89), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n807), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(new_n807), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n791), .A2(new_n792), .B1(new_n828), .B2(new_n830), .ZN(G311));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  INV_X1    g407(.A(new_n792), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n790), .ZN(G150));
  NAND2_X1  g409(.A1(new_n537), .A2(G55), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(new_n521), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT98), .B(G93), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n552), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n560), .A2(KEYINPUT99), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n558), .A2(new_n559), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(KEYINPUT99), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n850), .A3(G559), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(KEYINPUT38), .B1(new_n610), .B2(new_n618), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n849), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n856), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n848), .A3(new_n854), .ZN(new_n859));
  INV_X1    g434(.A(G860), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT100), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n857), .A2(new_n859), .A3(new_n863), .A4(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n840), .A2(G860), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT101), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT102), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n865), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G145));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n507), .A2(new_n508), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n507), .A2(KEYINPUT104), .A3(new_n508), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n498), .A2(new_n879), .A3(new_n512), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n498), .B2(new_n512), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n877), .B(new_n878), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n745), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n781), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n702), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(KEYINPUT105), .A3(new_n702), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n700), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n485), .A2(G142), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n470), .A2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(G130), .B2(new_n483), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n635), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(new_n814), .Z(new_n901));
  NAND2_X1  g476(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n890), .A2(new_n893), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(G162), .B(G160), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n631), .B(new_n905), .Z(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n890), .A2(new_n893), .A3(new_n903), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n903), .B1(new_n890), .B2(new_n893), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT107), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n894), .A2(KEYINPUT107), .A3(new_n901), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n906), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n874), .B(new_n908), .C1(new_n911), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT40), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n902), .A2(new_n904), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n906), .B(new_n912), .C1(new_n916), .C2(KEYINPUT107), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n874), .A4(new_n908), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(G395));
  XNOR2_X1  g495(.A(G303), .B(G288), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(G305), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(G290), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT42), .Z(new_n924));
  XNOR2_X1  g499(.A(new_n620), .B(new_n849), .ZN(new_n925));
  INV_X1    g500(.A(new_n606), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(new_n615), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n606), .A2(G299), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT41), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n925), .A2(new_n929), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n924), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n924), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g514(.A(new_n938), .B1(G868), .B2(new_n841), .ZN(G331));
  XNOR2_X1  g515(.A(G301), .B(KEYINPUT108), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n842), .A2(G286), .A3(new_n847), .ZN(new_n942));
  AOI21_X1  g517(.A(G286), .B1(new_n842), .B2(new_n847), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n848), .A2(G168), .ZN(new_n945));
  INV_X1    g520(.A(new_n941), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n842), .A2(G286), .A3(new_n847), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n933), .A2(new_n944), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n929), .B1(new_n944), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n923), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n923), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n933), .A2(new_n944), .A3(new_n948), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n944), .A2(new_n948), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n952), .B(new_n953), .C1(new_n954), .C2(new_n929), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n955), .A3(new_n874), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(new_n955), .A3(new_n958), .A4(new_n874), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT109), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n957), .A2(KEYINPUT109), .A3(KEYINPUT44), .A4(new_n959), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(G397));
  NAND2_X1  g540(.A1(new_n498), .A2(new_n512), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT103), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n498), .A2(new_n879), .A3(new_n512), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n507), .A2(KEYINPUT104), .A3(new_n508), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT104), .B1(new_n507), .B2(new_n508), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G1384), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n473), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT70), .B1(new_n480), .B2(G2105), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n474), .B(new_n470), .C1(new_n478), .C2(new_n479), .ZN(new_n976));
  OAI211_X1 g551(.A(G40), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n973), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n745), .B(G2067), .Z(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n781), .B(G1996), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n814), .B(new_n821), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(G290), .B(G1986), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT111), .Z(new_n990));
  XOR2_X1   g565(.A(KEYINPUT122), .B(KEYINPUT63), .Z(new_n991));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n513), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  AOI211_X1 g571(.A(KEYINPUT113), .B(new_n996), .C1(new_n513), .C2(new_n993), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G2090), .ZN(new_n999));
  INV_X1    g574(.A(new_n977), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n882), .A2(new_n996), .A3(new_n993), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n993), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n977), .B1(new_n1004), .B2(new_n994), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT112), .B(G1971), .Z(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G303), .A2(G8), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT55), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(G8), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1000), .A2(new_n882), .A3(new_n993), .ZN(new_n1015));
  INV_X1    g590(.A(G1976), .ZN(new_n1016));
  OR2_X1    g591(.A1(G288), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(G8), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT52), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n586), .A2(new_n591), .A3(new_n690), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1025));
  OAI211_X1 g600(.A(G1981), .B(G305), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1025), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G305), .A2(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1023), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1026), .A2(new_n1029), .A3(G8), .A4(new_n1015), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT114), .B(G1976), .Z(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1015), .A2(G8), .A3(new_n1017), .A4(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1019), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1014), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n996), .B1(new_n882), .B2(new_n993), .ZN(new_n1037));
  OAI211_X1 g612(.A(G160), .B(G40), .C1(new_n994), .C2(KEYINPUT50), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1037), .A2(G2090), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1007), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1041), .B2(new_n1012), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1036), .A3(new_n1012), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1035), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT45), .B1(new_n882), .B2(new_n993), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n977), .ZN(new_n1048));
  INV_X1    g623(.A(new_n994), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT45), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT119), .B(new_n1000), .C1(new_n973), .C2(KEYINPUT45), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1052), .A2(new_n752), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT113), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n994), .A2(new_n992), .A3(KEYINPUT50), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1001), .A2(new_n1056), .A3(new_n1000), .A4(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1054), .B1(new_n1058), .B2(G2084), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n977), .B1(new_n973), .B2(new_n996), .ZN(new_n1060));
  INV_X1    g635(.A(G2084), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(KEYINPUT120), .A3(new_n1061), .A4(new_n998), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(G8), .B(G168), .C1(new_n1053), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT121), .B1(new_n1045), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1019), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1067));
  INV_X1    g642(.A(G8), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1013), .B2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1041), .A2(new_n1036), .A3(new_n1012), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1042), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1072), .A2(new_n1064), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n991), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT63), .B1(new_n1069), .B2(new_n1013), .ZN(new_n1076));
  OR3_X1    g651(.A1(new_n1064), .A2(new_n1035), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(G286), .B1(new_n1053), .B2(new_n1063), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1052), .A2(new_n752), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1068), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT51), .B(new_n1079), .C1(new_n1082), .C2(KEYINPUT125), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(G168), .A3(new_n1081), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1085), .B(KEYINPUT51), .C1(KEYINPUT125), .C2(new_n1082), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1003), .A2(new_n1005), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(G299), .B(KEYINPUT57), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1015), .A2(G2067), .ZN(new_n1097));
  INV_X1    g672(.A(G1348), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1058), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n610), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1095), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(KEYINPUT123), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT123), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1109), .B(new_n1097), .C1(new_n1058), .C2(new_n1098), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1107), .A2(new_n1108), .B1(new_n1110), .B2(new_n610), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT124), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1099), .A2(KEYINPUT60), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1099), .A2(KEYINPUT60), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n611), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1096), .A2(new_n1116), .A3(KEYINPUT61), .A4(new_n1102), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1111), .A2(new_n1112), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1015), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT58), .B(G1341), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1006), .A2(G1996), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n560), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1122), .B(KEYINPUT59), .Z(new_n1123));
  OAI21_X1  g698(.A(new_n1106), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1003), .A2(new_n1005), .A3(new_n715), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT126), .B(KEYINPUT53), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n722), .A2(new_n1058), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n715), .A2(KEYINPUT53), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1052), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(G301), .B(KEYINPUT54), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G40), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1047), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1128), .B1(new_n973), .B2(KEYINPUT45), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n480), .A2(G2105), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n974), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1130), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1127), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1045), .A2(new_n1131), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1089), .A2(new_n1124), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1014), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1119), .A2(new_n1068), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT116), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1030), .ZN(new_n1144));
  NOR2_X1   g719(.A1(G288), .A2(G1976), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT117), .Z(new_n1146));
  OAI21_X1  g721(.A(new_n1020), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1141), .A2(new_n1034), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1078), .A2(new_n1140), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1087), .A2(new_n1150), .A3(new_n1088), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1150), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1045), .A2(G171), .A3(new_n1129), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n990), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n981), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n745), .A2(G2067), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n814), .A2(new_n820), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n985), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT46), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1156), .B2(G1996), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n981), .B1(new_n781), .B2(new_n983), .ZN(new_n1163));
  INV_X1    g738(.A(G1996), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n981), .A2(KEYINPUT46), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT47), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n981), .A2(new_n987), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1156), .A2(G1986), .A3(G290), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT48), .Z(new_n1172));
  AOI211_X1 g747(.A(new_n1160), .B(new_n1168), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1155), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g749(.A(G401), .B1(new_n957), .B2(new_n959), .ZN(new_n1176));
  NOR2_X1   g750(.A1(G227), .A2(new_n462), .ZN(new_n1177));
  XNOR2_X1  g751(.A(new_n1177), .B(KEYINPUT127), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n1178), .A2(G229), .ZN(new_n1179));
  AND3_X1   g753(.A1(new_n1176), .A2(new_n914), .A3(new_n1179), .ZN(G308));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n914), .A3(new_n1179), .ZN(G225));
endmodule


