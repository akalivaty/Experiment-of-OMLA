

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733;

  INV_X1 U368 ( .A(n588), .ZN(n349) );
  XNOR2_X1 U369 ( .A(n348), .B(n429), .ZN(n726) );
  NAND2_X1 U370 ( .A1(n404), .A2(n405), .ZN(n348) );
  OR2_X1 U371 ( .A1(n566), .A2(n370), .ZN(n376) );
  XNOR2_X1 U372 ( .A(n532), .B(n526), .ZN(n607) );
  OR2_X1 U373 ( .A1(n686), .A2(G902), .ZN(n367) );
  NOR2_X1 U374 ( .A1(n679), .A2(n649), .ZN(n467) );
  INV_X1 U375 ( .A(n350), .ZN(n595) );
  NAND2_X1 U376 ( .A1(n590), .A2(n350), .ZN(n420) );
  XNOR2_X2 U377 ( .A(n589), .B(n349), .ZN(n350) );
  INV_X1 U378 ( .A(G953), .ZN(n719) );
  NOR2_X2 U379 ( .A1(n426), .A2(n728), .ZN(n368) );
  XNOR2_X2 U380 ( .A(n715), .B(n461), .ZN(n470) );
  XNOR2_X2 U381 ( .A(n507), .B(n506), .ZN(n611) );
  XNOR2_X2 U382 ( .A(n541), .B(KEYINPUT38), .ZN(n620) );
  NAND2_X2 U383 ( .A1(n649), .A2(n648), .ZN(n650) );
  INV_X1 U384 ( .A(n649), .ZN(n488) );
  NOR2_X1 U385 ( .A1(n624), .A2(n623), .ZN(n377) );
  XNOR2_X1 U386 ( .A(n495), .B(n383), .ZN(n569) );
  NAND2_X1 U387 ( .A1(n567), .A2(n561), .ZN(n495) );
  NAND2_X1 U388 ( .A1(n400), .A2(n398), .ZN(n589) );
  XNOR2_X1 U389 ( .A(n373), .B(n401), .ZN(n400) );
  XNOR2_X1 U390 ( .A(n360), .B(KEYINPUT99), .ZN(n728) );
  XNOR2_X1 U391 ( .A(KEYINPUT104), .B(n518), .ZN(n730) );
  NOR2_X1 U392 ( .A1(n637), .A2(n543), .ZN(n364) );
  XNOR2_X1 U393 ( .A(n377), .B(n542), .ZN(n637) );
  XNOR2_X1 U394 ( .A(n522), .B(KEYINPUT96), .ZN(n669) );
  NOR2_X1 U395 ( .A1(n700), .A2(G902), .ZN(n366) );
  XNOR2_X1 U396 ( .A(n403), .B(n402), .ZN(n700) );
  AND2_X2 U397 ( .A1(n389), .A2(G472), .ZN(n652) );
  XNOR2_X1 U398 ( .A(n580), .B(n421), .ZN(n576) );
  XOR2_X1 U399 ( .A(G146), .B(G125), .Z(n462) );
  XNOR2_X1 U400 ( .A(n470), .B(n469), .ZN(n503) );
  XNOR2_X1 U401 ( .A(n714), .B(n468), .ZN(n469) );
  INV_X1 U402 ( .A(G146), .ZN(n468) );
  XNOR2_X1 U403 ( .A(n457), .B(n456), .ZN(n499) );
  NOR2_X1 U404 ( .A1(n576), .A2(n372), .ZN(n407) );
  INV_X1 U405 ( .A(n574), .ZN(n410) );
  OR2_X1 U406 ( .A1(n665), .A2(n625), .ZN(n535) );
  INV_X1 U407 ( .A(KEYINPUT44), .ZN(n401) );
  XNOR2_X1 U408 ( .A(n472), .B(n381), .ZN(n380) );
  INV_X1 U409 ( .A(KEYINPUT77), .ZN(n381) );
  XOR2_X1 U410 ( .A(G131), .B(G140), .Z(n473) );
  XNOR2_X1 U411 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U412 ( .A(n462), .B(KEYINPUT10), .ZN(n484) );
  XNOR2_X1 U413 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n444) );
  XNOR2_X1 U414 ( .A(n391), .B(n703), .ZN(n679) );
  XNOR2_X1 U415 ( .A(n470), .B(n465), .ZN(n391) );
  INV_X1 U416 ( .A(KEYINPUT2), .ZN(n419) );
  NOR2_X1 U417 ( .A1(n636), .A2(n574), .ZN(n406) );
  NAND2_X1 U418 ( .A1(n565), .A2(n371), .ZN(n370) );
  XNOR2_X1 U419 ( .A(n564), .B(n563), .ZN(n566) );
  XNOR2_X1 U420 ( .A(n562), .B(KEYINPUT73), .ZN(n563) );
  INV_X1 U421 ( .A(KEYINPUT89), .ZN(n421) );
  BUF_X1 U422 ( .A(n611), .Z(n378) );
  NOR2_X1 U423 ( .A1(G952), .A2(n719), .ZN(n702) );
  INV_X1 U424 ( .A(KEYINPUT46), .ZN(n412) );
  NAND2_X1 U425 ( .A1(n352), .A2(n394), .ZN(n359) );
  INV_X1 U426 ( .A(n730), .ZN(n394) );
  XOR2_X1 U427 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n497) );
  XOR2_X1 U428 ( .A(G137), .B(G134), .Z(n714) );
  XNOR2_X1 U429 ( .A(G116), .B(G113), .ZN(n455) );
  NOR2_X1 U430 ( .A1(G953), .A2(G237), .ZN(n436) );
  XNOR2_X1 U431 ( .A(n484), .B(n473), .ZN(n713) );
  XNOR2_X1 U432 ( .A(G143), .B(G113), .ZN(n433) );
  XOR2_X1 U433 ( .A(G122), .B(G104), .Z(n434) );
  XNOR2_X1 U434 ( .A(n425), .B(n424), .ZN(n423) );
  XNOR2_X1 U435 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n425) );
  XNOR2_X1 U436 ( .A(KEYINPUT87), .B(KEYINPUT78), .ZN(n424) );
  INV_X1 U437 ( .A(KEYINPUT45), .ZN(n588) );
  NAND2_X1 U438 ( .A1(G234), .A2(G237), .ZN(n510) );
  BUF_X1 U439 ( .A(n636), .Z(n365) );
  OR2_X1 U440 ( .A1(G237), .A2(G902), .ZN(n508) );
  NAND2_X1 U441 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U442 ( .A1(n576), .A2(n372), .ZN(n408) );
  NOR2_X1 U443 ( .A1(n603), .A2(n623), .ZN(n384) );
  INV_X1 U444 ( .A(n519), .ZN(n417) );
  XNOR2_X1 U445 ( .A(n441), .B(n440), .ZN(n442) );
  INV_X1 U446 ( .A(KEYINPUT66), .ZN(n383) );
  XNOR2_X1 U447 ( .A(G134), .B(G116), .ZN(n446) );
  XOR2_X1 U448 ( .A(G122), .B(G107), .Z(n447) );
  XNOR2_X1 U449 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U450 ( .A(n380), .B(n471), .ZN(n475) );
  NAND2_X1 U451 ( .A1(n418), .A2(n416), .ZN(n544) );
  XNOR2_X1 U452 ( .A(n509), .B(n379), .ZN(n418) );
  NOR2_X1 U453 ( .A1(n577), .A2(n417), .ZN(n416) );
  INV_X1 U454 ( .A(KEYINPUT30), .ZN(n379) );
  XNOR2_X1 U455 ( .A(n533), .B(KEYINPUT107), .ZN(n537) );
  XNOR2_X1 U456 ( .A(n361), .B(n355), .ZN(n531) );
  XOR2_X1 U457 ( .A(KEYINPUT6), .B(n611), .Z(n584) );
  XNOR2_X1 U458 ( .A(n499), .B(n390), .ZN(n703) );
  XNOR2_X1 U459 ( .A(n471), .B(n459), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n484), .B(n485), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n487), .B(n486), .ZN(n403) );
  XNOR2_X1 U462 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n485) );
  AND2_X1 U463 ( .A1(n388), .A2(n386), .ZN(n682) );
  INV_X1 U464 ( .A(G210), .ZN(n387) );
  NOR2_X1 U465 ( .A1(n546), .A2(n541), .ZN(n525) );
  INV_X1 U466 ( .A(KEYINPUT35), .ZN(n429) );
  XNOR2_X1 U467 ( .A(n428), .B(KEYINPUT32), .ZN(n427) );
  INV_X1 U468 ( .A(KEYINPUT65), .ZN(n428) );
  NAND2_X1 U469 ( .A1(n586), .A2(n568), .ZN(n360) );
  INV_X1 U470 ( .A(n702), .ZN(n374) );
  XNOR2_X1 U471 ( .A(n695), .B(n357), .ZN(n375) );
  BUF_X1 U472 ( .A(n607), .Z(n362) );
  XOR2_X1 U473 ( .A(KEYINPUT4), .B(KEYINPUT67), .Z(n351) );
  OR2_X1 U474 ( .A1(KEYINPUT47), .A2(n535), .ZN(n352) );
  XOR2_X1 U475 ( .A(KEYINPUT69), .B(G469), .Z(n353) );
  AND2_X1 U476 ( .A1(n375), .A2(n374), .ZN(n354) );
  XOR2_X1 U477 ( .A(KEYINPUT28), .B(n530), .Z(n355) );
  INV_X1 U478 ( .A(KEYINPUT34), .ZN(n372) );
  XOR2_X1 U479 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n356) );
  XOR2_X1 U480 ( .A(n694), .B(n693), .Z(n357) );
  XOR2_X1 U481 ( .A(n688), .B(n687), .Z(n358) );
  NAND2_X1 U482 ( .A1(n524), .A2(n619), .ZN(n546) );
  NOR2_X1 U483 ( .A1(n359), .A2(n536), .ZN(n393) );
  NAND2_X1 U484 ( .A1(n593), .A2(KEYINPUT2), .ZN(n594) );
  XNOR2_X1 U485 ( .A(n594), .B(KEYINPUT85), .ZN(n596) );
  XNOR2_X1 U486 ( .A(n364), .B(KEYINPUT42), .ZN(n732) );
  NAND2_X1 U487 ( .A1(n611), .A2(n529), .ZN(n361) );
  INV_X1 U488 ( .A(n537), .ZN(n543) );
  INV_X1 U489 ( .A(n620), .ZN(n397) );
  NOR2_X1 U490 ( .A1(n583), .A2(n399), .ZN(n398) );
  NOR2_X1 U491 ( .A1(n653), .A2(n702), .ZN(n655) );
  NOR2_X2 U492 ( .A1(n607), .A2(n608), .ZN(n579) );
  NAND2_X1 U493 ( .A1(n363), .A2(n410), .ZN(n404) );
  NAND2_X1 U494 ( .A1(n409), .A2(n408), .ZN(n363) );
  NAND2_X1 U495 ( .A1(n385), .A2(n384), .ZN(n564) );
  XNOR2_X2 U496 ( .A(n366), .B(n382), .ZN(n567) );
  XNOR2_X2 U497 ( .A(n593), .B(KEYINPUT84), .ZN(n590) );
  AND2_X2 U498 ( .A1(n553), .A2(n552), .ZN(n593) );
  INV_X1 U499 ( .A(n733), .ZN(n399) );
  NAND2_X1 U500 ( .A1(n406), .A2(n407), .ZN(n405) );
  XNOR2_X2 U501 ( .A(n367), .B(n353), .ZN(n532) );
  INV_X1 U502 ( .A(n550), .ZN(n541) );
  XNOR2_X2 U503 ( .A(n467), .B(n466), .ZN(n550) );
  NAND2_X1 U504 ( .A1(n559), .A2(n560), .ZN(n422) );
  NAND2_X1 U505 ( .A1(n369), .A2(n368), .ZN(n373) );
  INV_X1 U506 ( .A(n726), .ZN(n369) );
  INV_X1 U507 ( .A(n362), .ZN(n371) );
  NOR2_X2 U508 ( .A1(n566), .A2(n371), .ZN(n586) );
  XNOR2_X2 U509 ( .A(n376), .B(n427), .ZN(n729) );
  NAND2_X1 U510 ( .A1(n493), .A2(G217), .ZN(n490) );
  XNOR2_X1 U511 ( .A(n489), .B(KEYINPUT20), .ZN(n493) );
  XNOR2_X1 U512 ( .A(n492), .B(KEYINPUT91), .ZN(n382) );
  NAND2_X1 U513 ( .A1(n569), .A2(n532), .ZN(n577) );
  XNOR2_X1 U514 ( .A(n392), .B(n356), .ZN(n553) );
  XOR2_X2 U515 ( .A(G902), .B(KEYINPUT15), .Z(n649) );
  XNOR2_X1 U516 ( .A(n354), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U517 ( .A(n580), .ZN(n385) );
  NOR2_X4 U518 ( .A1(n650), .A2(n430), .ZN(n389) );
  NOR2_X1 U519 ( .A1(n430), .A2(n387), .ZN(n386) );
  INV_X1 U520 ( .A(n650), .ZN(n388) );
  NAND2_X1 U521 ( .A1(n389), .A2(G475), .ZN(n695) );
  NAND2_X1 U522 ( .A1(n389), .A2(G478), .ZN(n696) );
  NAND2_X1 U523 ( .A1(n389), .A2(G217), .ZN(n699) );
  NAND2_X1 U524 ( .A1(n389), .A2(G469), .ZN(n690) );
  XNOR2_X2 U525 ( .A(n460), .B(n351), .ZN(n715) );
  NAND2_X1 U526 ( .A1(n395), .A2(n393), .ZN(n392) );
  XNOR2_X1 U527 ( .A(n396), .B(n412), .ZN(n395) );
  NAND2_X1 U528 ( .A1(n414), .A2(n413), .ZN(n396) );
  NOR2_X1 U529 ( .A1(n544), .A2(n397), .ZN(n415) );
  NAND2_X1 U530 ( .A1(n636), .A2(n372), .ZN(n409) );
  NOR2_X1 U531 ( .A1(n702), .A2(n684), .ZN(n685) );
  NAND2_X1 U532 ( .A1(n596), .A2(n350), .ZN(n648) );
  XNOR2_X2 U533 ( .A(n411), .B(G143), .ZN(n460) );
  XNOR2_X2 U534 ( .A(KEYINPUT64), .B(G128), .ZN(n411) );
  INV_X1 U535 ( .A(n731), .ZN(n413) );
  INV_X1 U536 ( .A(n732), .ZN(n414) );
  XNOR2_X1 U537 ( .A(n415), .B(KEYINPUT39), .ZN(n551) );
  INV_X1 U538 ( .A(n590), .ZN(n718) );
  AND2_X2 U539 ( .A1(n420), .A2(n419), .ZN(n430) );
  XNOR2_X2 U540 ( .A(n422), .B(KEYINPUT0), .ZN(n580) );
  XNOR2_X2 U541 ( .A(n528), .B(KEYINPUT19), .ZN(n559) );
  XNOR2_X1 U542 ( .A(n423), .B(n462), .ZN(n464) );
  INV_X1 U543 ( .A(n729), .ZN(n426) );
  XNOR2_X2 U544 ( .A(n573), .B(n572), .ZN(n636) );
  AND2_X1 U545 ( .A1(G214), .A2(n496), .ZN(n431) );
  XOR2_X1 U546 ( .A(n651), .B(KEYINPUT62), .Z(n432) );
  XNOR2_X1 U547 ( .A(n497), .B(G131), .ZN(n498) );
  XNOR2_X1 U548 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U549 ( .A(KEYINPUT3), .ZN(n454) );
  XNOR2_X1 U550 ( .A(n437), .B(n431), .ZN(n438) );
  INV_X1 U551 ( .A(G475), .ZN(n440) );
  XNOR2_X1 U552 ( .A(n439), .B(n438), .ZN(n692) );
  NAND2_X1 U553 ( .A1(n550), .A2(n619), .ZN(n528) );
  XNOR2_X1 U554 ( .A(n503), .B(n476), .ZN(n686) );
  XNOR2_X1 U555 ( .A(n443), .B(n442), .ZN(n521) );
  NOR2_X1 U556 ( .A1(n540), .A2(n538), .ZN(n522) );
  XNOR2_X1 U557 ( .A(n686), .B(n358), .ZN(n689) );
  XNOR2_X1 U558 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U559 ( .A(n647), .B(n646), .ZN(G75) );
  XNOR2_X1 U560 ( .A(n713), .B(KEYINPUT12), .ZN(n439) );
  XNOR2_X1 U561 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U562 ( .A(n435), .B(KEYINPUT11), .Z(n437) );
  XOR2_X1 U563 ( .A(KEYINPUT75), .B(n436), .Z(n496) );
  NOR2_X1 U564 ( .A1(G902), .A2(n692), .ZN(n443) );
  XNOR2_X1 U565 ( .A(KEYINPUT13), .B(KEYINPUT95), .ZN(n441) );
  NAND2_X1 U566 ( .A1(n719), .A2(G234), .ZN(n445) );
  XNOR2_X1 U567 ( .A(n445), .B(n444), .ZN(n477) );
  NAND2_X1 U568 ( .A1(n477), .A2(G217), .ZN(n452) );
  XNOR2_X1 U569 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U570 ( .A(n448), .B(KEYINPUT9), .Z(n450) );
  XNOR2_X1 U571 ( .A(n460), .B(KEYINPUT7), .ZN(n449) );
  XNOR2_X1 U572 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U573 ( .A(n452), .B(n451), .ZN(n697) );
  NOR2_X1 U574 ( .A1(G902), .A2(n697), .ZN(n453) );
  XOR2_X1 U575 ( .A(G478), .B(n453), .Z(n538) );
  NAND2_X1 U576 ( .A1(n521), .A2(n538), .ZN(n574) );
  XOR2_X1 U577 ( .A(G122), .B(KEYINPUT16), .Z(n459) );
  XNOR2_X1 U578 ( .A(n455), .B(n454), .ZN(n457) );
  XOR2_X1 U579 ( .A(KEYINPUT70), .B(G119), .Z(n456) );
  XNOR2_X1 U580 ( .A(G104), .B(G110), .ZN(n458) );
  XNOR2_X1 U581 ( .A(n458), .B(G107), .ZN(n471) );
  INV_X1 U582 ( .A(G101), .ZN(n461) );
  NAND2_X1 U583 ( .A1(G224), .A2(n719), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U585 ( .A1(G210), .A2(n508), .ZN(n466) );
  NAND2_X1 U586 ( .A1(G227), .A2(n719), .ZN(n472) );
  INV_X1 U587 ( .A(n473), .ZN(n474) );
  NAND2_X1 U588 ( .A1(n477), .A2(G221), .ZN(n487) );
  XOR2_X1 U589 ( .A(G110), .B(G140), .Z(n479) );
  XNOR2_X1 U590 ( .A(G128), .B(G137), .ZN(n478) );
  XNOR2_X1 U591 ( .A(n479), .B(n478), .ZN(n483) );
  XOR2_X1 U592 ( .A(KEYINPUT76), .B(KEYINPUT71), .Z(n481) );
  XNOR2_X1 U593 ( .A(G119), .B(KEYINPUT23), .ZN(n480) );
  XNOR2_X1 U594 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U595 ( .A(n483), .B(n482), .ZN(n486) );
  XOR2_X1 U596 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n491) );
  NAND2_X1 U597 ( .A1(G234), .A2(n488), .ZN(n489) );
  XNOR2_X1 U598 ( .A(n491), .B(n490), .ZN(n492) );
  NAND2_X1 U599 ( .A1(G221), .A2(n493), .ZN(n494) );
  XOR2_X1 U600 ( .A(KEYINPUT21), .B(n494), .Z(n561) );
  NAND2_X1 U601 ( .A1(n496), .A2(G210), .ZN(n501) );
  XOR2_X1 U602 ( .A(n501), .B(n500), .Z(n502) );
  XNOR2_X1 U603 ( .A(n503), .B(n502), .ZN(n651) );
  NOR2_X1 U604 ( .A1(n651), .A2(G902), .ZN(n507) );
  XNOR2_X1 U605 ( .A(KEYINPUT72), .B(KEYINPUT94), .ZN(n505) );
  INV_X1 U606 ( .A(G472), .ZN(n504) );
  NAND2_X1 U607 ( .A1(G214), .A2(n508), .ZN(n619) );
  NAND2_X1 U608 ( .A1(n611), .A2(n619), .ZN(n509) );
  XNOR2_X1 U609 ( .A(n510), .B(KEYINPUT14), .ZN(n512) );
  NAND2_X1 U610 ( .A1(G952), .A2(n512), .ZN(n511) );
  XOR2_X1 U611 ( .A(KEYINPUT88), .B(n511), .Z(n634) );
  NAND2_X1 U612 ( .A1(n719), .A2(n634), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G902), .A2(n512), .ZN(n555) );
  NOR2_X1 U614 ( .A1(G900), .A2(n555), .ZN(n513) );
  NAND2_X1 U615 ( .A1(G953), .A2(n513), .ZN(n514) );
  NAND2_X1 U616 ( .A1(n557), .A2(n514), .ZN(n515) );
  XOR2_X1 U617 ( .A(KEYINPUT79), .B(n515), .Z(n519) );
  NOR2_X1 U618 ( .A1(n541), .A2(n544), .ZN(n516) );
  XNOR2_X1 U619 ( .A(n516), .B(KEYINPUT103), .ZN(n517) );
  NOR2_X1 U620 ( .A1(n574), .A2(n517), .ZN(n518) );
  INV_X1 U621 ( .A(n584), .ZN(n554) );
  NAND2_X1 U622 ( .A1(n561), .A2(n519), .ZN(n520) );
  NOR2_X1 U623 ( .A1(n567), .A2(n520), .ZN(n529) );
  INV_X1 U624 ( .A(n521), .ZN(n540) );
  NAND2_X1 U625 ( .A1(n529), .A2(n669), .ZN(n523) );
  NOR2_X1 U626 ( .A1(n554), .A2(n523), .ZN(n524) );
  XNOR2_X1 U627 ( .A(n525), .B(KEYINPUT36), .ZN(n527) );
  INV_X1 U628 ( .A(KEYINPUT1), .ZN(n526) );
  NAND2_X1 U629 ( .A1(n527), .A2(n371), .ZN(n676) );
  XOR2_X1 U630 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n530) );
  NAND2_X1 U631 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U632 ( .A1(n559), .A2(n537), .ZN(n665) );
  NAND2_X1 U633 ( .A1(n538), .A2(n540), .ZN(n662) );
  INV_X1 U634 ( .A(n662), .ZN(n671) );
  NOR2_X1 U635 ( .A1(n669), .A2(n671), .ZN(n625) );
  NAND2_X1 U636 ( .A1(KEYINPUT47), .A2(n535), .ZN(n534) );
  NAND2_X1 U637 ( .A1(n676), .A2(n534), .ZN(n536) );
  INV_X1 U638 ( .A(n538), .ZN(n539) );
  NAND2_X1 U639 ( .A1(n540), .A2(n539), .ZN(n623) );
  XNOR2_X1 U640 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n542) );
  INV_X1 U641 ( .A(n669), .ZN(n666) );
  NOR2_X1 U642 ( .A1(n551), .A2(n666), .ZN(n545) );
  XNOR2_X1 U643 ( .A(n545), .B(KEYINPUT40), .ZN(n731) );
  XNOR2_X1 U644 ( .A(n546), .B(KEYINPUT102), .ZN(n547) );
  NOR2_X1 U645 ( .A1(n371), .A2(n547), .ZN(n548) );
  XNOR2_X1 U646 ( .A(n548), .B(KEYINPUT43), .ZN(n549) );
  NOR2_X1 U647 ( .A1(n550), .A2(n549), .ZN(n678) );
  NOR2_X1 U648 ( .A1(n662), .A2(n551), .ZN(n677) );
  NOR2_X1 U649 ( .A1(n678), .A2(n677), .ZN(n552) );
  XNOR2_X1 U650 ( .A(KEYINPUT97), .B(n567), .ZN(n602) );
  AND2_X1 U651 ( .A1(n602), .A2(n554), .ZN(n565) );
  NOR2_X1 U652 ( .A1(G898), .A2(n719), .ZN(n705) );
  INV_X1 U653 ( .A(n555), .ZN(n556) );
  NAND2_X1 U654 ( .A1(n705), .A2(n556), .ZN(n558) );
  NAND2_X1 U655 ( .A1(n558), .A2(n557), .ZN(n560) );
  INV_X1 U656 ( .A(n561), .ZN(n603) );
  XOR2_X1 U657 ( .A(KEYINPUT74), .B(KEYINPUT22), .Z(n562) );
  NOR2_X1 U658 ( .A1(n567), .A2(n378), .ZN(n568) );
  INV_X1 U659 ( .A(n569), .ZN(n608) );
  XNOR2_X1 U660 ( .A(n579), .B(KEYINPUT100), .ZN(n570) );
  NAND2_X1 U661 ( .A1(n570), .A2(n584), .ZN(n573) );
  XNOR2_X1 U662 ( .A(KEYINPUT33), .B(KEYINPUT101), .ZN(n571) );
  XNOR2_X1 U663 ( .A(n571), .B(KEYINPUT86), .ZN(n572) );
  OR2_X1 U664 ( .A1(n378), .A2(n576), .ZN(n578) );
  NOR2_X1 U665 ( .A1(n578), .A2(n577), .ZN(n657) );
  NAND2_X1 U666 ( .A1(n378), .A2(n579), .ZN(n616) );
  NOR2_X1 U667 ( .A1(n580), .A2(n616), .ZN(n581) );
  XOR2_X1 U668 ( .A(KEYINPUT31), .B(n581), .Z(n672) );
  NOR2_X1 U669 ( .A1(n657), .A2(n672), .ZN(n582) );
  NOR2_X1 U670 ( .A1(n625), .A2(n582), .ZN(n583) );
  NOR2_X1 U671 ( .A1(n602), .A2(n584), .ZN(n585) );
  NAND2_X1 U672 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U673 ( .A(KEYINPUT98), .B(n587), .ZN(n733) );
  NAND2_X1 U674 ( .A1(n430), .A2(KEYINPUT82), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n595), .A2(n590), .ZN(n591) );
  NOR2_X1 U676 ( .A1(KEYINPUT2), .A2(n591), .ZN(n592) );
  NOR2_X1 U677 ( .A1(KEYINPUT82), .A2(n592), .ZN(n598) );
  INV_X1 U678 ( .A(n648), .ZN(n597) );
  NOR2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X1 U680 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT83), .ZN(n643) );
  XOR2_X1 U682 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n605) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n605), .B(n604), .ZN(n606) );
  XOR2_X1 U685 ( .A(KEYINPUT112), .B(n606), .Z(n614) );
  XOR2_X1 U686 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n610) );
  NAND2_X1 U687 ( .A1(n608), .A2(n362), .ZN(n609) );
  XNOR2_X1 U688 ( .A(n610), .B(n609), .ZN(n612) );
  NOR2_X1 U689 ( .A1(n612), .A2(n378), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U692 ( .A(KEYINPUT51), .B(n617), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n637), .A2(n618), .ZN(n631) );
  NOR2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U695 ( .A(KEYINPUT115), .B(n621), .Z(n622) );
  NOR2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n628) );
  NOR2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n626), .B(KEYINPUT116), .ZN(n627) );
  NOR2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U700 ( .A1(n365), .A2(n629), .ZN(n630) );
  NOR2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U702 ( .A(KEYINPUT117), .B(n632), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n633), .B(KEYINPUT52), .ZN(n635) );
  AND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n640) );
  NOR2_X1 U705 ( .A1(n637), .A2(n365), .ZN(n638) );
  XNOR2_X1 U706 ( .A(KEYINPUT118), .B(n638), .ZN(n639) );
  NOR2_X1 U707 ( .A1(n640), .A2(n639), .ZN(n641) );
  AND2_X1 U708 ( .A1(n641), .A2(n719), .ZN(n642) );
  NAND2_X1 U709 ( .A1(n643), .A2(n642), .ZN(n647) );
  XOR2_X1 U710 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n645) );
  INV_X1 U711 ( .A(KEYINPUT119), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n652), .B(n432), .ZN(n653) );
  INV_X1 U714 ( .A(KEYINPUT63), .ZN(n654) );
  XNOR2_X1 U715 ( .A(n655), .B(n654), .ZN(G57) );
  NAND2_X1 U716 ( .A1(n669), .A2(n657), .ZN(n656) );
  XNOR2_X1 U717 ( .A(n656), .B(G104), .ZN(G6) );
  XOR2_X1 U718 ( .A(G107), .B(KEYINPUT27), .Z(n659) );
  NAND2_X1 U719 ( .A1(n657), .A2(n671), .ZN(n658) );
  XNOR2_X1 U720 ( .A(n659), .B(n658), .ZN(n661) );
  XOR2_X1 U721 ( .A(KEYINPUT109), .B(KEYINPUT26), .Z(n660) );
  XNOR2_X1 U722 ( .A(n661), .B(n660), .ZN(G9) );
  NOR2_X1 U723 ( .A1(n662), .A2(n665), .ZN(n663) );
  XNOR2_X1 U724 ( .A(G128), .B(n663), .ZN(n664) );
  XNOR2_X1 U725 ( .A(n664), .B(KEYINPUT29), .ZN(G30) );
  NOR2_X1 U726 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U727 ( .A(G146), .B(n667), .Z(n668) );
  XNOR2_X1 U728 ( .A(KEYINPUT110), .B(n668), .ZN(G48) );
  NAND2_X1 U729 ( .A1(n669), .A2(n672), .ZN(n670) );
  XNOR2_X1 U730 ( .A(n670), .B(G113), .ZN(G15) );
  XOR2_X1 U731 ( .A(G116), .B(KEYINPUT111), .Z(n674) );
  NAND2_X1 U732 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U733 ( .A(n674), .B(n673), .ZN(G18) );
  XOR2_X1 U734 ( .A(G125), .B(KEYINPUT37), .Z(n675) );
  XNOR2_X1 U735 ( .A(n676), .B(n675), .ZN(G27) );
  XOR2_X1 U736 ( .A(G134), .B(n677), .Z(G36) );
  XOR2_X1 U737 ( .A(G140), .B(n678), .Z(G42) );
  XNOR2_X1 U738 ( .A(KEYINPUT55), .B(KEYINPUT80), .ZN(n681) );
  XNOR2_X1 U739 ( .A(n679), .B(KEYINPUT54), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n681), .B(n680), .ZN(n683) );
  XNOR2_X1 U741 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U742 ( .A(KEYINPUT56), .B(n685), .ZN(G51) );
  XOR2_X1 U743 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n688) );
  XNOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n687) );
  NOR2_X1 U745 ( .A1(n702), .A2(n691), .ZN(G54) );
  XNOR2_X1 U746 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n694) );
  XNOR2_X1 U747 ( .A(n692), .B(KEYINPUT123), .ZN(n693) );
  XNOR2_X1 U748 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U749 ( .A1(n702), .A2(n698), .ZN(G63) );
  XNOR2_X1 U750 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U751 ( .A1(n702), .A2(n701), .ZN(G66) );
  XOR2_X1 U752 ( .A(G101), .B(n703), .Z(n704) );
  NOR2_X1 U753 ( .A1(n705), .A2(n704), .ZN(n712) );
  XOR2_X1 U754 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n707) );
  NAND2_X1 U755 ( .A1(G224), .A2(G953), .ZN(n706) );
  XNOR2_X1 U756 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U757 ( .A1(n708), .A2(G898), .ZN(n710) );
  NAND2_X1 U758 ( .A1(n350), .A2(n719), .ZN(n709) );
  NAND2_X1 U759 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U760 ( .A(n712), .B(n711), .ZN(G69) );
  XNOR2_X1 U761 ( .A(n713), .B(KEYINPUT126), .ZN(n717) );
  XNOR2_X1 U762 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U763 ( .A(n717), .B(n716), .ZN(n721) );
  XNOR2_X1 U764 ( .A(n721), .B(n718), .ZN(n720) );
  NAND2_X1 U765 ( .A1(n720), .A2(n719), .ZN(n725) );
  XNOR2_X1 U766 ( .A(G227), .B(n721), .ZN(n722) );
  NAND2_X1 U767 ( .A1(n722), .A2(G900), .ZN(n723) );
  NAND2_X1 U768 ( .A1(n723), .A2(G953), .ZN(n724) );
  NAND2_X1 U769 ( .A1(n725), .A2(n724), .ZN(G72) );
  XNOR2_X1 U770 ( .A(n726), .B(G122), .ZN(n727) );
  XNOR2_X1 U771 ( .A(n727), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U772 ( .A(n728), .B(G110), .Z(G12) );
  XNOR2_X1 U773 ( .A(n729), .B(G119), .ZN(G21) );
  XOR2_X1 U774 ( .A(n730), .B(G143), .Z(G45) );
  XOR2_X1 U775 ( .A(n731), .B(G131), .Z(G33) );
  XOR2_X1 U776 ( .A(n732), .B(G137), .Z(G39) );
  XNOR2_X1 U777 ( .A(G101), .B(n733), .ZN(G3) );
endmodule

