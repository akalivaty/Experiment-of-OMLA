//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n205), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n215), .B1(new_n216), .B2(new_n205), .C1(new_n217), .C2(new_n212), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  AND2_X1   g0020(.A1(G77), .A2(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR4_X1   g0024(.A1(new_n218), .A2(new_n220), .A3(new_n221), .A4(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT64), .B(G68), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G238), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n208), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n214), .B(new_n229), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  OAI211_X1 g0052(.A(G1), .B(G13), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n259));
  OAI21_X1  g0059(.A(G226), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n223), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n257), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G97), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n254), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n252), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n206), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n253), .ZN(new_n271));
  INV_X1    g0071(.A(G238), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n269), .A2(KEYINPUT66), .A3(new_n206), .A4(G274), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT70), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT70), .B1(new_n277), .B2(new_n278), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n267), .A2(new_n274), .A3(new_n279), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT13), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT70), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n280), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT13), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(new_n267), .A4(new_n274), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n283), .A2(KEYINPUT71), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT71), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(new_n289), .A3(KEYINPUT13), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G179), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n287), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT14), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n283), .B2(new_n287), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT14), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n292), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n209), .A2(new_n207), .A3(G1), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT12), .B1(new_n302), .B2(new_n226), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT72), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n302), .A2(KEYINPUT12), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n304), .B1(G68), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n230), .ZN(new_n308));
  INV_X1    g0108(.A(G50), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G20), .A2(G33), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n226), .A2(new_n207), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n207), .A2(G33), .ZN(new_n313));
  INV_X1    g0113(.A(G77), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n308), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT11), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n308), .B1(new_n206), .B2(G20), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n306), .B(new_n317), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n300), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT67), .B(G1698), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n262), .B1(new_n324), .B2(G226), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n265), .B1(new_n325), .B2(new_n257), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n273), .B1(new_n326), .B2(new_n254), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n286), .B1(new_n327), .B2(new_n285), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n290), .ZN(new_n330));
  OAI21_X1  g0130(.A(G190), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n321), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n293), .A2(G200), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n322), .A2(KEYINPUT73), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT69), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n277), .A2(new_n278), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n270), .A2(new_n253), .A3(G244), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(KEYINPUT68), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT68), .B1(new_n338), .B2(new_n339), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n257), .A2(new_n217), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n258), .A2(new_n259), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n345), .A2(new_n223), .B1(new_n272), .B2(new_n261), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n254), .B(new_n344), .C1(new_n346), .C2(new_n257), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n337), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n302), .A2(G77), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n310), .B1(G20), .B2(G77), .ZN(new_n352));
  XOR2_X1   g0152(.A(KEYINPUT15), .B(G87), .Z(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n313), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n349), .B1(new_n355), .B2(new_n308), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n319), .A2(G77), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n336), .B1(new_n348), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n342), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n347), .A3(new_n340), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G200), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n362), .A2(KEYINPUT69), .A3(new_n357), .A4(new_n356), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n359), .B(new_n363), .C1(new_n364), .C2(new_n361), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n343), .A2(new_n366), .A3(new_n347), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n361), .A2(new_n296), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n358), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n324), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n370));
  OR2_X1    g0170(.A1(KEYINPUT3), .A2(G33), .ZN(new_n371));
  NAND2_X1  g0171(.A1(KEYINPUT3), .A2(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n253), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(G77), .B2(new_n373), .ZN(new_n375));
  INV_X1    g0175(.A(new_n271), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G226), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n338), .A3(new_n377), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(G179), .ZN(new_n379));
  INV_X1    g0179(.A(G150), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n350), .A2(new_n313), .B1(new_n380), .B2(new_n311), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n207), .B1(new_n201), .B2(new_n309), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n308), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n319), .A2(G50), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n384), .C1(G50), .C2(new_n302), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n378), .A2(new_n296), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n335), .A2(new_n365), .A3(new_n369), .A4(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n385), .B(KEYINPUT9), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n378), .A2(G200), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n364), .C2(new_n378), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(KEYINPUT10), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(KEYINPUT10), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n311), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n201), .B1(new_n226), .B2(G58), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n207), .ZN(new_n400));
  INV_X1    g0200(.A(new_n226), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n371), .A2(new_n207), .A3(new_n372), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n371), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n372), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n395), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT75), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n318), .A2(KEYINPUT64), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT64), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G68), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n411), .A3(G58), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n207), .B1(new_n412), .B2(new_n202), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT74), .B1(new_n413), .B2(new_n397), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(new_n398), .C1(new_n399), .C2(new_n207), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT7), .B1(new_n257), .B2(new_n207), .ZN(new_n417));
  INV_X1    g0217(.A(new_n405), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n414), .A2(new_n416), .A3(new_n419), .A4(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(new_n395), .C1(new_n400), .C2(new_n406), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n408), .A2(new_n308), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT76), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n270), .A2(new_n253), .A3(G232), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n338), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n338), .B2(new_n425), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(G223), .B1(new_n258), .B2(new_n259), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G226), .A2(G1698), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n257), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n251), .A2(new_n216), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n254), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(new_n364), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n338), .A3(new_n425), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n337), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n351), .A2(new_n301), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n320), .B2(new_n351), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n423), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT17), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n226), .B1(new_n417), .B2(new_n418), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n412), .A2(new_n202), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n397), .B1(new_n445), .B2(G20), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n421), .B1(new_n447), .B2(new_n395), .ZN(new_n448));
  AOI211_X1 g0248(.A(KEYINPUT75), .B(KEYINPUT16), .C1(new_n444), .C2(new_n446), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n420), .A2(new_n308), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n439), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n428), .A2(KEYINPUT77), .A3(new_n366), .A4(new_n433), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n338), .A2(new_n425), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT76), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n338), .A2(new_n424), .A3(new_n425), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n433), .A3(new_n456), .A4(new_n366), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT77), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n435), .A2(new_n296), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n453), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n443), .B1(new_n452), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n453), .A2(new_n459), .A3(new_n460), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n423), .A2(new_n440), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT18), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n394), .A2(new_n442), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT73), .B1(new_n322), .B2(new_n334), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n388), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n302), .A2(G116), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n308), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n302), .B(new_n472), .C1(G1), .C2(new_n251), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G116), .ZN(new_n475));
  AOI21_X1  g0275(.A(G20), .B1(G33), .B2(G283), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n251), .A2(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT82), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n472), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G20), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT20), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n480), .B1(new_n476), .B2(new_n477), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n308), .B(new_n484), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n471), .B(new_n475), .C1(new_n485), .C2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n206), .B(G45), .C1(new_n252), .C2(KEYINPUT5), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT79), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G41), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT79), .A3(new_n206), .A4(G45), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(G270), .A3(new_n253), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n494), .A2(new_n498), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(G274), .A3(new_n253), .A4(new_n495), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G264), .A2(G1698), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n373), .B(new_n504), .C1(new_n345), .C2(new_n211), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n505), .B(new_n254), .C1(G303), .C2(new_n373), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT81), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n499), .A2(new_n507), .A3(G270), .A4(new_n253), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n501), .A2(new_n503), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n491), .A2(new_n509), .A3(G169), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT21), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT83), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n509), .A2(KEYINPUT21), .A3(G169), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n503), .A2(new_n506), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(G179), .A3(new_n501), .A4(new_n508), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n491), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT83), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(new_n519), .A3(new_n511), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n509), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(new_n491), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n364), .C2(new_n509), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n513), .A2(new_n518), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(G238), .B1(new_n258), .B2(new_n259), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G244), .A2(G1698), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n257), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n251), .A2(new_n483), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n254), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n253), .B(G250), .C1(G1), .C2(new_n268), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT80), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n530), .A2(KEYINPUT80), .A3(new_n531), .A4(new_n532), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n366), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n251), .A2(G20), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G97), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n207), .B1(new_n265), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n216), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n540), .A2(new_n541), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n373), .A2(new_n207), .A3(G68), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n308), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n302), .B2(new_n353), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n473), .A2(new_n354), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n535), .A2(new_n296), .A3(new_n536), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n538), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n537), .A2(G190), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n535), .A2(G200), .A3(new_n536), .ZN(new_n556));
  OAI221_X1 g0356(.A(new_n548), .B1(new_n216), .B2(new_n473), .C1(new_n302), .C2(new_n353), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  OAI21_X1  g0362(.A(G244), .B1(new_n258), .B2(new_n259), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(new_n257), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n373), .A2(new_n324), .A3(KEYINPUT4), .A4(G244), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G283), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n373), .A2(G250), .A3(G1698), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n254), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n499), .A2(G257), .A3(new_n253), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n503), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n473), .A2(new_n219), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n574));
  AND2_X1   g0374(.A1(G97), .A2(G107), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n543), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n576), .B2(KEYINPUT6), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G20), .B1(G77), .B2(new_n310), .ZN(new_n578));
  OAI21_X1  g0378(.A(G107), .B1(new_n417), .B2(new_n418), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n573), .B1(new_n580), .B2(new_n308), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n301), .A2(new_n219), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n582), .B(KEYINPUT78), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n569), .A2(G190), .A3(new_n503), .A4(new_n570), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n572), .A2(new_n581), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n583), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n571), .A2(new_n296), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n569), .A2(new_n366), .A3(new_n503), .A4(new_n570), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT86), .ZN(new_n591));
  OAI21_X1  g0391(.A(G250), .B1(new_n258), .B2(new_n259), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G257), .A2(G1698), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n257), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G294), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n251), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n254), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n499), .A2(G264), .A3(new_n253), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n503), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n591), .B1(new_n600), .B2(G200), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n499), .A2(new_n253), .ZN(new_n602));
  AOI22_X1  g0402(.A1(G264), .A2(new_n602), .B1(new_n597), .B2(KEYINPUT85), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT85), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n604), .B(new_n254), .C1(new_n594), .C2(new_n596), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n603), .A2(new_n364), .A3(new_n503), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n599), .A2(KEYINPUT86), .A3(new_n337), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n601), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n539), .A2(G116), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n207), .A2(G107), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT23), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n207), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n612), .A2(KEYINPUT22), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(KEYINPUT22), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n609), .B(new_n611), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT24), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n612), .B(KEYINPUT22), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(KEYINPUT24), .A3(new_n609), .A4(new_n611), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n619), .A3(new_n308), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n301), .A2(new_n217), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT84), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT25), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n474), .A2(G107), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n608), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n597), .A2(KEYINPUT85), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n503), .A3(new_n605), .A4(new_n598), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G169), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n600), .A2(G179), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n625), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n590), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n469), .A2(new_n525), .A3(new_n561), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(KEYINPUT92), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n291), .A2(G179), .B1(new_n298), .B2(new_n297), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n332), .B1(new_n637), .B2(new_n295), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n321), .B1(new_n291), .B2(G190), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n369), .B1(new_n639), .B2(new_n333), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT90), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n369), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n334), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n322), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n645), .A3(new_n442), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n466), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n394), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n392), .A2(KEYINPUT91), .A3(new_n393), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n636), .B1(new_n653), .B2(new_n387), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n646), .B2(new_n466), .ZN(new_n655));
  INV_X1    g0455(.A(new_n387), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n655), .A2(KEYINPUT92), .A3(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n513), .A2(new_n518), .A3(new_n520), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT87), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT87), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n513), .A2(new_n518), .A3(new_n661), .A4(new_n520), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n632), .A2(new_n663), .A3(new_n625), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n632), .B2(new_n625), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n660), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n533), .A2(new_n296), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n538), .A2(new_n552), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n533), .A2(G200), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n555), .A2(new_n558), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n590), .A2(new_n627), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n669), .ZN(new_n675));
  INV_X1    g0475(.A(new_n589), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n554), .A2(new_n559), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n675), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n581), .A2(new_n583), .B1(new_n571), .B2(new_n296), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT89), .B1(new_n679), .B2(new_n588), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT89), .A4(new_n588), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n551), .B1(new_n537), .B2(new_n366), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n557), .B1(new_n537), .B2(G190), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n685), .A2(new_n668), .B1(new_n686), .B2(new_n670), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n678), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n674), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n469), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n658), .A2(new_n691), .ZN(G369));
  NOR2_X1   g0492(.A1(new_n209), .A2(G20), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n206), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI211_X1 g0500(.A(new_n522), .B(new_n700), .C1(new_n660), .C2(new_n662), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n524), .B1(new_n491), .B2(new_n699), .ZN(new_n702));
  OAI21_X1  g0502(.A(G330), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n627), .B(new_n633), .C1(new_n626), .C2(new_n700), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT93), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n633), .B2(new_n700), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n700), .B1(new_n664), .B2(new_n665), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n659), .A2(new_n700), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(G399));
  NOR2_X1   g0512(.A1(new_n210), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n544), .A2(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n232), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT94), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n684), .B1(new_n683), .B2(new_n687), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n554), .A2(new_n559), .A3(new_n676), .A4(new_n684), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n669), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n513), .A2(new_n518), .A3(new_n633), .A4(new_n520), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n673), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n699), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI211_X1 g0528(.A(KEYINPUT29), .B(new_n699), .C1(new_n674), .C2(new_n689), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n634), .A2(new_n525), .A3(new_n561), .A4(new_n700), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n509), .A2(new_n366), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n569), .A2(new_n570), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n599), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n733), .A3(new_n537), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n731), .A2(new_n537), .A3(new_n733), .A4(KEYINPUT30), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n509), .A2(new_n571), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n366), .A3(new_n533), .A4(new_n599), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n699), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n730), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n728), .B(new_n729), .C1(G330), .C2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n719), .B1(new_n746), .B2(G1), .ZN(G364));
  NAND2_X1  g0547(.A1(new_n693), .A2(G45), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n714), .A2(G1), .A3(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n701), .A2(G330), .A3(new_n702), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n749), .B1(new_n704), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n749), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n701), .A2(new_n702), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n230), .B1(G20), .B2(new_n296), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n207), .A2(new_n364), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n366), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n207), .A2(G190), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n337), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G322), .A2(new_n762), .B1(new_n766), .B2(G283), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G329), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n767), .A2(new_n257), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n366), .A2(new_n337), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n759), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT98), .B(G326), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n763), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n760), .A2(new_n763), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n779), .A2(new_n780), .B1(new_n782), .B2(G311), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n768), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n777), .B(new_n783), .C1(new_n595), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n759), .A2(new_n764), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G303), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n373), .B1(new_n778), .B2(new_n318), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT97), .B(G159), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n770), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT32), .Z(new_n794));
  NOR2_X1   g0594(.A1(new_n786), .A2(new_n219), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G50), .B2(new_n775), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n766), .A2(G107), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G58), .A2(new_n762), .B1(new_n789), .B2(G87), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n794), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n791), .B(new_n799), .C1(G77), .C2(new_n782), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n758), .B1(new_n790), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n233), .A2(new_n268), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n210), .A2(new_n373), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n246), .C2(new_n268), .ZN(new_n804));
  INV_X1    g0604(.A(new_n210), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n373), .ZN(new_n806));
  XNOR2_X1  g0606(.A(G355), .B(KEYINPUT95), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n804), .B1(G116), .B2(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n755), .A2(new_n758), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT96), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n801), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n752), .B1(new_n757), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n751), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT99), .Z(G396));
  AND3_X1   g0615(.A1(new_n745), .A2(KEYINPUT102), .A3(G330), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT102), .B1(new_n745), .B2(G330), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT101), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n369), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n358), .A2(new_n367), .A3(new_n368), .A4(KEYINPUT101), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n365), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n690), .A2(new_n700), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n699), .B1(new_n674), .B2(new_n689), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n358), .A2(new_n699), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n822), .A2(new_n365), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n642), .A2(new_n699), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n825), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n752), .B1(new_n818), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n831), .B2(new_n817), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n828), .A2(new_n753), .A3(new_n829), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n781), .A2(new_n483), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n835), .B(new_n795), .C1(G107), .C2(new_n789), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n779), .A2(G283), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n373), .B1(new_n762), .B2(G294), .ZN(new_n838));
  INV_X1    g0638(.A(G303), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n774), .A2(new_n839), .B1(new_n765), .B2(new_n216), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G311), .B2(new_n770), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n765), .A2(new_n318), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G132), .B2(new_n770), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n844), .B(new_n373), .C1(new_n309), .C2(new_n788), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G58), .B2(new_n785), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT100), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G143), .A2(new_n762), .B1(new_n782), .B2(new_n792), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n849), .B2(new_n774), .C1(new_n380), .C2(new_n778), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT34), .Z(new_n851));
  OAI21_X1  g0651(.A(new_n842), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n758), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n758), .A2(new_n753), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n314), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n834), .A2(new_n752), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n833), .A2(new_n856), .ZN(G384));
  INV_X1    g0657(.A(new_n697), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n414), .A2(new_n416), .A3(new_n419), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n395), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n439), .B1(new_n451), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n452), .A2(new_n443), .A3(new_n461), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT18), .B1(new_n463), .B2(new_n464), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT17), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n441), .B(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n858), .B(new_n862), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n861), .B1(new_n461), .B2(new_n697), .ZN(new_n869));
  INV_X1    g0669(.A(new_n441), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n463), .A2(new_n464), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT105), .B1(new_n464), .B2(new_n858), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n874), .B(new_n697), .C1(new_n423), .C2(new_n440), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n441), .B(new_n872), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n871), .B1(new_n876), .B2(KEYINPUT37), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n868), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n873), .A2(new_n875), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n441), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n874), .B1(new_n452), .B2(new_n697), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n464), .A2(KEYINPUT105), .A3(new_n858), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n872), .A2(new_n441), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n442), .A2(new_n466), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n880), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT106), .B1(new_n879), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n321), .A2(new_n699), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n322), .A2(new_n334), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT104), .B1(new_n638), .B2(new_n699), .ZN(new_n896));
  AND4_X1   g0696(.A1(KEYINPUT104), .A2(new_n300), .A3(new_n321), .A4(new_n699), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n745), .A2(new_n898), .A3(new_n830), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT106), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n882), .A2(new_n888), .B1(new_n890), .B2(new_n880), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n878), .B(new_n900), .C1(new_n901), .C2(KEYINPUT38), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n893), .A2(KEYINPUT40), .A3(new_n899), .A4(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n868), .B2(new_n877), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n879), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n745), .A2(new_n898), .A3(new_n830), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT107), .Z(new_n910));
  NAND2_X1  g0710(.A1(new_n469), .A2(new_n745), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(G330), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n469), .B1(new_n729), .B2(new_n728), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n658), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n879), .B2(new_n892), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n322), .A2(new_n699), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n868), .A2(new_n877), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(KEYINPUT39), .A3(new_n878), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n917), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n878), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n699), .B(new_n823), .C1(new_n674), .C2(new_n689), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n822), .A2(new_n699), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n924), .B(new_n898), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n865), .A2(new_n697), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n923), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n915), .B(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n913), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n206), .B2(new_n693), .ZN(new_n932));
  OAI211_X1 g0732(.A(G116), .B(new_n231), .C1(new_n577), .C2(KEYINPUT35), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT103), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n233), .A2(G77), .A3(new_n412), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(G50), .B2(new_n318), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(G1), .A3(new_n209), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n932), .A2(new_n937), .A3(new_n940), .ZN(G367));
  NAND2_X1  g0741(.A1(new_n586), .A2(new_n699), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n590), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n676), .A2(new_n699), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n706), .A2(new_n710), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n589), .B1(new_n943), .B2(new_n633), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n700), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n687), .B1(new_n558), .B2(new_n700), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n675), .A2(new_n557), .A3(new_n699), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n952), .A2(KEYINPUT43), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n708), .A2(new_n946), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n952), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n956), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n957), .B1(new_n956), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n713), .B(KEYINPUT41), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n711), .A2(new_n709), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n966), .B1(new_n967), .B2(new_n946), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n711), .A2(KEYINPUT45), .A3(new_n709), .A4(new_n945), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT44), .B1(new_n967), .B2(new_n946), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n967), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n708), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n970), .B(new_n708), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  INV_X1    g0776(.A(new_n710), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n711), .B1(new_n707), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(new_n704), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n979), .A2(new_n746), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n975), .A2(new_n976), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n965), .B1(new_n981), .B2(new_n746), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n748), .A2(G1), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n963), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT108), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT108), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n963), .B(new_n986), .C1(new_n982), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n810), .B1(new_n805), .B2(new_n354), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n241), .A2(new_n210), .A3(new_n373), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n752), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT109), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n373), .B1(new_n785), .B2(G107), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n766), .A2(G97), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n595), .C2(new_n778), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n789), .A2(G116), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT46), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n996), .A2(new_n997), .B1(G311), .B2(new_n775), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G303), .A2(new_n762), .B1(new_n782), .B2(G283), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n997), .C2(new_n996), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n995), .B(new_n1000), .C1(G317), .C2(new_n770), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n762), .A2(G150), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n792), .A2(new_n779), .B1(new_n782), .B2(G50), .ZN(new_n1003));
  INV_X1    g0803(.A(G143), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n318), .B2(new_n786), .C1(new_n1004), .C2(new_n774), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n373), .B1(new_n769), .B2(new_n849), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n788), .A2(new_n222), .B1(new_n765), .B2(new_n314), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1001), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n758), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n992), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT110), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n756), .B2(new_n955), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n988), .A2(new_n1014), .ZN(G387));
  NOR2_X1   g0815(.A1(new_n980), .A2(new_n714), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n746), .B2(new_n979), .ZN(new_n1017));
  OR3_X1    g0817(.A1(new_n350), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT50), .B1(new_n350), .B2(G50), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1018), .A2(new_n1019), .A3(new_n268), .A4(new_n715), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n318), .A2(new_n314), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n803), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT112), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n268), .B2(new_n238), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(G107), .B2(new_n805), .C1(new_n715), .C2(new_n806), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n749), .B1(new_n1025), .B2(new_n810), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n786), .A2(new_n354), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n789), .A2(G77), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n782), .A2(G68), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n770), .A2(G150), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n994), .B1(new_n309), .B2(new_n761), .C1(new_n396), .C2(new_n774), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n778), .A2(new_n350), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n257), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G322), .A2(new_n775), .B1(new_n779), .B2(G311), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n839), .B2(new_n781), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G317), .B2(new_n762), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT48), .Z(new_n1039));
  INV_X1    g0839(.A(G283), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n786), .C1(new_n595), .C2(new_n788), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT49), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n765), .A2(new_n483), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n373), .B(new_n1043), .C1(new_n770), .C2(new_n776), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1035), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1026), .B1(new_n707), .B2(new_n756), .C1(new_n1045), .C2(new_n1011), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n979), .A2(new_n983), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT111), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1017), .A2(new_n1046), .A3(new_n1048), .ZN(G393));
  NAND3_X1  g0849(.A1(new_n975), .A2(new_n983), .A3(new_n976), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n810), .B1(new_n219), .B2(new_n805), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n249), .B2(new_n803), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n774), .A2(new_n380), .B1(new_n761), .B2(new_n396), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n257), .B1(new_n789), .B2(new_n226), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n765), .A2(new_n216), .B1(new_n769), .B2(new_n1004), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G77), .B2(new_n785), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n778), .A2(new_n309), .B1(new_n781), .B2(new_n350), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT113), .Z(new_n1060));
  AOI22_X1  g0860(.A1(G317), .A2(new_n775), .B1(new_n762), .B2(G311), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT52), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n257), .B1(new_n781), .B2(new_n595), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G303), .B2(new_n779), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n785), .A2(G116), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G283), .A2(new_n789), .B1(new_n770), .B2(G322), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1064), .A2(new_n797), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1058), .A2(new_n1060), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n749), .B(new_n1052), .C1(new_n1068), .C2(new_n758), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT114), .Z(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n756), .B2(new_n945), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n980), .B1(new_n975), .B2(new_n976), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT115), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n981), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n713), .B1(new_n1072), .B2(KEYINPUT115), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1050), .B(new_n1071), .C1(new_n1074), .C2(new_n1075), .ZN(G390));
  NAND2_X1  g0876(.A1(new_n917), .A2(new_n922), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n753), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT54), .B(G143), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT118), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1081), .A2(new_n782), .B1(G132), .B2(new_n762), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1082), .B(new_n373), .C1(new_n309), .C2(new_n765), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n778), .A2(new_n849), .ZN(new_n1084));
  INV_X1    g0884(.A(G125), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n769), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n786), .A2(new_n396), .ZN(new_n1087));
  NOR4_X1   g0887(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n788), .A2(new_n380), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT53), .ZN(new_n1090));
  INV_X1    g0890(.A(G128), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1090), .C1(new_n1091), .C2(new_n774), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT119), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n770), .A2(G294), .B1(new_n785), .B2(G77), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n216), .B2(new_n788), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n843), .B(new_n1095), .C1(G283), .C2(new_n775), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1096), .B(new_n257), .C1(new_n483), .C2(new_n761), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n778), .A2(new_n217), .B1(new_n781), .B2(new_n219), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT120), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1093), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT121), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n758), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n854), .A2(new_n350), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1078), .A2(new_n1102), .A3(new_n752), .A4(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n745), .A2(new_n898), .A3(G330), .A4(new_n830), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n898), .B1(new_n925), .B2(new_n926), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n918), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1107), .A2(new_n1108), .B1(new_n917), .B2(new_n922), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT89), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n589), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1111), .A2(new_n669), .A3(new_n671), .A4(new_n681), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT26), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n669), .A3(new_n721), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n724), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1115), .A2(new_n672), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n700), .B(new_n824), .C1(new_n1114), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n926), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n898), .ZN(new_n1120));
  AND4_X1   g0920(.A1(new_n893), .A2(new_n1120), .A3(new_n902), .A4(new_n1108), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1106), .B1(new_n1109), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n898), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n825), .B2(new_n1118), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1077), .B1(new_n1124), .B2(new_n918), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1120), .A2(new_n893), .A3(new_n902), .A4(new_n1108), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n1105), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n983), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1104), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT116), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n830), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1132), .B(new_n895), .C1(new_n896), .C2(new_n897), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n744), .A2(new_n741), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n590), .A2(new_n627), .A3(new_n633), .ZN(new_n1136));
  NOR4_X1   g0936(.A1(new_n1136), .A2(new_n524), .A3(new_n560), .A4(new_n699), .ZN(new_n1137));
  OAI211_X1 g0937(.A(G330), .B(new_n830), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n926), .B1(new_n726), .B2(new_n824), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1133), .A2(G330), .A3(new_n745), .A4(new_n830), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1123), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1143), .A2(new_n1105), .B1(new_n825), .B2(new_n1118), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n469), .A2(G330), .A3(new_n745), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n914), .B(new_n1146), .C1(new_n654), .C2(new_n657), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(KEYINPUT117), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT117), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1150), .B1(new_n1128), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1130), .B1(new_n1155), .B2(new_n713), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(new_n1147), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1149), .A2(new_n1158), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n903), .A2(G330), .A3(new_n908), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n923), .A2(new_n927), .A3(new_n928), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n903), .A2(G330), .A3(new_n908), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n929), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n651), .A2(new_n656), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n385), .A2(new_n858), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1162), .A2(new_n1164), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1173), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n929), .A2(new_n1163), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1159), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n714), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1159), .A2(KEYINPUT57), .A3(new_n1174), .A4(new_n1178), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n753), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n309), .B1(new_n255), .B2(G41), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n779), .A2(G97), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n762), .A2(G107), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1029), .A2(new_n1186), .A3(new_n1187), .A4(new_n252), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n765), .A2(new_n222), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT122), .Z(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1188), .B(new_n1191), .C1(G283), .C2(new_n770), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n782), .A2(new_n353), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n786), .A2(new_n318), .B1(new_n774), .B2(new_n483), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT123), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n257), .A3(new_n1193), .A4(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT58), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n1080), .A2(new_n788), .B1(new_n1091), .B2(new_n761), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT124), .Z(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n1085), .B2(new_n774), .C1(new_n380), .C2(new_n786), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G132), .B2(new_n779), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n849), .B2(new_n781), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1202), .B(new_n1203), .Z(new_n1204));
  AOI21_X1  g1004(.A(G33), .B1(new_n766), .B2(new_n792), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n770), .A2(G124), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n252), .A3(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1185), .B(new_n1197), .C1(new_n1204), .C2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n758), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n854), .A2(new_n309), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1184), .A2(new_n752), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT126), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1178), .A2(new_n1174), .A3(new_n983), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1183), .A2(new_n1215), .ZN(G375));
  NAND2_X1  g1016(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1154), .A2(new_n964), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1123), .A2(new_n753), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n373), .B1(new_n770), .B2(G303), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n314), .B2(new_n765), .C1(new_n483), .C2(new_n778), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1027), .B1(G294), .B2(new_n775), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n217), .B2(new_n781), .C1(new_n1040), .C2(new_n761), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(G97), .C2(new_n789), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G159), .A2(new_n789), .B1(new_n782), .B2(G150), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n257), .B1(new_n762), .B2(G137), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n309), .C2(new_n786), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n775), .A2(G132), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1190), .B(new_n1228), .C1(new_n778), .C2(new_n1080), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(G128), .C2(new_n770), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n758), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n854), .A2(new_n318), .ZN(new_n1232));
  AND4_X1   g1032(.A1(new_n752), .A2(new_n1219), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1145), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n983), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1218), .A2(new_n1235), .ZN(G381));
  AOI21_X1  g1036(.A(new_n1214), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1156), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1238), .A2(G384), .A3(G381), .ZN(new_n1239));
  INV_X1    g1039(.A(G390), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n988), .A2(new_n1014), .A3(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G393), .A2(G396), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .ZN(G407));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(G343), .C2(new_n1238), .ZN(G409));
  NAND4_X1  g1044(.A1(new_n1159), .A2(new_n964), .A3(new_n1174), .A4(new_n1178), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1245), .A2(new_n1213), .A3(new_n1212), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1156), .ZN(new_n1247));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G343), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1247), .B(new_n1250), .C1(new_n1237), .C2(new_n1156), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1145), .A2(new_n1147), .A3(KEYINPUT60), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n713), .C1(new_n1147), .C2(new_n1145), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT60), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1235), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n833), .A3(new_n856), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G384), .B(new_n1235), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1249), .A2(G2897), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1258), .B(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT61), .B1(new_n1251), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1249), .B1(new_n1246), .B2(new_n1156), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n1156), .C2(new_n1237), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT62), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G375), .A2(G378), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1263), .A4(new_n1262), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n1265), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1240), .B1(new_n988), .B2(new_n1014), .ZN(new_n1272));
  AND2_X1   g1072(.A1(G393), .A2(G396), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1241), .A2(new_n1272), .B1(new_n1242), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G387), .A2(G390), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n988), .A2(new_n1014), .A3(new_n1240), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1273), .A2(new_n1242), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1261), .A2(new_n1265), .A3(KEYINPUT127), .A4(new_n1268), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1271), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1251), .B2(new_n1260), .ZN(new_n1283));
  MUX2_X1   g1083(.A(new_n1282), .B(new_n1283), .S(new_n1264), .Z(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1274), .B2(new_n1278), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1281), .A2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(new_n1266), .A2(new_n1238), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1263), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1289), .B(new_n1290), .ZN(G402));
endmodule


