

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586;

  NAND2_X1 U319 ( .A1(n534), .A2(n503), .ZN(n463) );
  INV_X1 U320 ( .A(n525), .ZN(n503) );
  XNOR2_X2 U321 ( .A(n456), .B(n455), .ZN(n582) );
  XOR2_X2 U322 ( .A(n481), .B(KEYINPUT41), .Z(n556) );
  NOR2_X1 U323 ( .A1(n413), .A2(n500), .ZN(n453) );
  XNOR2_X1 U324 ( .A(n452), .B(KEYINPUT26), .ZN(n553) );
  XNOR2_X1 U325 ( .A(n359), .B(KEYINPUT47), .ZN(n360) );
  XNOR2_X1 U326 ( .A(n347), .B(n346), .ZN(n353) );
  INV_X1 U327 ( .A(n553), .ZN(n454) );
  XNOR2_X1 U328 ( .A(n384), .B(n383), .ZN(n386) );
  XNOR2_X1 U329 ( .A(n437), .B(n382), .ZN(n383) );
  XNOR2_X1 U330 ( .A(n379), .B(n378), .ZN(n384) );
  XOR2_X1 U331 ( .A(G113GAT), .B(G71GAT), .Z(n287) );
  XOR2_X1 U332 ( .A(G204GAT), .B(KEYINPUT70), .Z(n288) );
  AND2_X1 U333 ( .A1(n575), .A2(n556), .ZN(n355) );
  NOR2_X1 U334 ( .A1(n553), .A2(n471), .ZN(n461) );
  INV_X1 U335 ( .A(KEYINPUT114), .ZN(n359) );
  XNOR2_X1 U336 ( .A(n340), .B(KEYINPUT31), .ZN(n341) );
  XNOR2_X1 U337 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U338 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U339 ( .A(n368), .B(KEYINPUT48), .ZN(n551) );
  XNOR2_X1 U340 ( .A(n437), .B(n287), .ZN(n438) );
  XNOR2_X1 U341 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U342 ( .A(n439), .B(n438), .ZN(n447) );
  INV_X1 U343 ( .A(G204GAT), .ZN(n457) );
  XOR2_X1 U344 ( .A(n386), .B(n385), .Z(n525) );
  XNOR2_X1 U345 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U346 ( .A(n484), .B(G43GAT), .ZN(n485) );
  XNOR2_X1 U347 ( .A(n460), .B(n459), .ZN(G1353GAT) );
  XNOR2_X1 U348 ( .A(n486), .B(n485), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(G162GAT), .B(G50GAT), .Z(n427) );
  XOR2_X1 U350 ( .A(G190GAT), .B(G36GAT), .Z(n377) );
  XNOR2_X1 U351 ( .A(n427), .B(n377), .ZN(n291) );
  XOR2_X1 U352 ( .A(G43GAT), .B(KEYINPUT8), .Z(n290) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n289) );
  XNOR2_X1 U354 ( .A(n290), .B(n289), .ZN(n323) );
  XNOR2_X1 U355 ( .A(n291), .B(n323), .ZN(n295) );
  XOR2_X1 U356 ( .A(KEYINPUT11), .B(G92GAT), .Z(n293) );
  NAND2_X1 U357 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U358 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U359 ( .A(n295), .B(n294), .Z(n300) );
  XOR2_X1 U360 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n297) );
  XNOR2_X1 U361 ( .A(KEYINPUT9), .B(KEYINPUT64), .ZN(n296) );
  XNOR2_X1 U362 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U363 ( .A(G134GAT), .B(n298), .ZN(n299) );
  XNOR2_X1 U364 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U365 ( .A(G85GAT), .B(G99GAT), .Z(n349) );
  XOR2_X1 U366 ( .A(n301), .B(n349), .Z(n303) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(G106GAT), .ZN(n302) );
  XOR2_X1 U368 ( .A(n303), .B(n302), .Z(n563) );
  INV_X1 U369 ( .A(n563), .ZN(n546) );
  XOR2_X1 U370 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n305) );
  XNOR2_X1 U371 ( .A(KEYINPUT76), .B(KEYINPUT14), .ZN(n304) );
  XNOR2_X1 U372 ( .A(n305), .B(n304), .ZN(n311) );
  XOR2_X1 U373 ( .A(KEYINPUT13), .B(G71GAT), .Z(n307) );
  XNOR2_X1 U374 ( .A(G57GAT), .B(G78GAT), .ZN(n306) );
  XNOR2_X1 U375 ( .A(n307), .B(n306), .ZN(n342) );
  XOR2_X1 U376 ( .A(G155GAT), .B(G22GAT), .Z(n417) );
  XOR2_X1 U377 ( .A(n342), .B(n417), .Z(n309) );
  NAND2_X1 U378 ( .A1(G231GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U379 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U380 ( .A(n311), .B(n310), .ZN(n322) );
  XOR2_X1 U381 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n313) );
  XNOR2_X1 U382 ( .A(KEYINPUT12), .B(KEYINPUT77), .ZN(n312) );
  XNOR2_X1 U383 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U384 ( .A(n314), .B(G64GAT), .Z(n316) );
  XOR2_X1 U385 ( .A(G127GAT), .B(G15GAT), .Z(n434) );
  XNOR2_X1 U386 ( .A(G1GAT), .B(n434), .ZN(n315) );
  XNOR2_X1 U387 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U388 ( .A(n317), .B(KEYINPUT74), .Z(n320) );
  XNOR2_X1 U389 ( .A(G211GAT), .B(G183GAT), .ZN(n318) );
  XOR2_X1 U390 ( .A(n318), .B(G8GAT), .Z(n385) );
  XOR2_X1 U391 ( .A(n385), .B(KEYINPUT79), .Z(n319) );
  XNOR2_X1 U392 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U393 ( .A(n322), .B(n321), .ZN(n579) );
  XOR2_X1 U394 ( .A(n579), .B(KEYINPUT112), .Z(n573) );
  XOR2_X1 U395 ( .A(G113GAT), .B(G1GAT), .Z(n404) );
  XOR2_X1 U396 ( .A(n323), .B(n404), .Z(n325) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U398 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U399 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n327) );
  XNOR2_X1 U400 ( .A(KEYINPUT66), .B(KEYINPUT65), .ZN(n326) );
  XNOR2_X1 U401 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U402 ( .A(n329), .B(n328), .Z(n337) );
  XOR2_X1 U403 ( .A(G197GAT), .B(G36GAT), .Z(n331) );
  XNOR2_X1 U404 ( .A(G141GAT), .B(G50GAT), .ZN(n330) );
  XNOR2_X1 U405 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U406 ( .A(G169GAT), .B(G15GAT), .Z(n333) );
  XNOR2_X1 U407 ( .A(G8GAT), .B(G22GAT), .ZN(n332) );
  XNOR2_X1 U408 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U409 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U410 ( .A(n337), .B(n336), .Z(n575) );
  XNOR2_X1 U411 ( .A(G92GAT), .B(G176GAT), .ZN(n338) );
  XNOR2_X1 U412 ( .A(n288), .B(n338), .ZN(n339) );
  XNOR2_X1 U413 ( .A(n339), .B(G64GAT), .ZN(n373) );
  INV_X1 U414 ( .A(n373), .ZN(n371) );
  AND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U416 ( .A(n343), .B(G120GAT), .ZN(n347) );
  XOR2_X1 U417 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n345) );
  XNOR2_X1 U418 ( .A(KEYINPUT71), .B(KEYINPUT32), .ZN(n344) );
  XNOR2_X1 U419 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U420 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U422 ( .A(G148GAT), .B(G106GAT), .Z(n416) );
  XNOR2_X1 U423 ( .A(n350), .B(n416), .ZN(n351) );
  XOR2_X1 U424 ( .A(n351), .B(KEYINPUT67), .Z(n352) );
  XNOR2_X1 U425 ( .A(n371), .B(n354), .ZN(n481) );
  XOR2_X1 U426 ( .A(KEYINPUT46), .B(n355), .Z(n356) );
  NAND2_X1 U427 ( .A1(n573), .A2(n356), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n357), .B(KEYINPUT113), .ZN(n358) );
  NAND2_X1 U429 ( .A1(n358), .A2(n546), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n367) );
  XNOR2_X1 U431 ( .A(KEYINPUT36), .B(n563), .ZN(n583) );
  NAND2_X1 U432 ( .A1(n583), .A2(n579), .ZN(n362) );
  XNOR2_X1 U433 ( .A(KEYINPUT45), .B(n362), .ZN(n363) );
  NOR2_X1 U434 ( .A1(n481), .A2(n363), .ZN(n364) );
  XOR2_X1 U435 ( .A(KEYINPUT115), .B(n364), .Z(n365) );
  INV_X1 U436 ( .A(n575), .ZN(n566) );
  NAND2_X1 U437 ( .A1(n365), .A2(n566), .ZN(n366) );
  NAND2_X1 U438 ( .A1(n367), .A2(n366), .ZN(n368) );
  XOR2_X1 U439 ( .A(G197GAT), .B(KEYINPUT21), .Z(n370) );
  XNOR2_X1 U440 ( .A(G218GAT), .B(KEYINPUT85), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n370), .B(n369), .ZN(n414) );
  NAND2_X1 U442 ( .A1(n371), .A2(n414), .ZN(n375) );
  INV_X1 U443 ( .A(n414), .ZN(n372) );
  NAND2_X1 U444 ( .A1(n373), .A2(n372), .ZN(n374) );
  NAND2_X1 U445 ( .A1(n375), .A2(n374), .ZN(n379) );
  XOR2_X1 U446 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n376) );
  XOR2_X1 U447 ( .A(G169GAT), .B(KEYINPUT19), .Z(n381) );
  XNOR2_X1 U448 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n437) );
  AND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  NAND2_X1 U451 ( .A1(n551), .A2(n503), .ZN(n388) );
  XOR2_X1 U452 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n387) );
  XOR2_X1 U453 ( .A(n388), .B(n387), .Z(n413) );
  XOR2_X1 U454 ( .A(G141GAT), .B(KEYINPUT2), .Z(n390) );
  XNOR2_X1 U455 ( .A(KEYINPUT3), .B(KEYINPUT86), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n415) );
  XOR2_X1 U457 ( .A(G120GAT), .B(KEYINPUT0), .Z(n392) );
  XNOR2_X1 U458 ( .A(G134GAT), .B(KEYINPUT82), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n433) );
  XNOR2_X1 U460 ( .A(n415), .B(n433), .ZN(n412) );
  XOR2_X1 U461 ( .A(KEYINPUT89), .B(G57GAT), .Z(n394) );
  XNOR2_X1 U462 ( .A(G155GAT), .B(G127GAT), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U464 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n396) );
  XNOR2_X1 U465 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U467 ( .A(n398), .B(n397), .Z(n410) );
  XOR2_X1 U468 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n400) );
  XNOR2_X1 U469 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n399) );
  XNOR2_X1 U470 ( .A(n400), .B(n399), .ZN(n408) );
  XOR2_X1 U471 ( .A(G148GAT), .B(G85GAT), .Z(n402) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(G162GAT), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U474 ( .A(n404), .B(n403), .Z(n406) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U476 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U478 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U479 ( .A(n412), .B(n411), .Z(n522) );
  INV_X1 U480 ( .A(n522), .ZN(n500) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n431) );
  XOR2_X1 U482 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U485 ( .A(KEYINPUT24), .B(G204GAT), .Z(n421) );
  XNOR2_X1 U486 ( .A(G211GAT), .B(G78GAT), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U488 ( .A(n423), .B(n422), .Z(n429) );
  XOR2_X1 U489 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n425) );
  XNOR2_X1 U490 ( .A(KEYINPUT88), .B(KEYINPUT22), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U494 ( .A(n431), .B(n430), .Z(n473) );
  INV_X1 U495 ( .A(n473), .ZN(n462) );
  NAND2_X1 U496 ( .A1(n453), .A2(n462), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n432), .B(KEYINPUT55), .ZN(n448) );
  XOR2_X1 U498 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n436), .B(n435), .ZN(n439) );
  XOR2_X1 U501 ( .A(KEYINPUT20), .B(G43GAT), .Z(n441) );
  XNOR2_X1 U502 ( .A(G99GAT), .B(G190GAT), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT84), .Z(n443) );
  XNOR2_X1 U505 ( .A(G183GAT), .B(KEYINPUT83), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U507 ( .A(n445), .B(n444), .Z(n446) );
  XOR2_X1 U508 ( .A(n447), .B(n446), .Z(n527) );
  INV_X1 U509 ( .A(n527), .ZN(n534) );
  NAND2_X1 U510 ( .A1(n448), .A2(n534), .ZN(n572) );
  NOR2_X1 U511 ( .A1(n546), .A2(n572), .ZN(n451) );
  XNOR2_X1 U512 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n449), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U514 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  NAND2_X1 U515 ( .A1(n473), .A2(n527), .ZN(n452) );
  NAND2_X1 U516 ( .A1(n454), .A2(n453), .ZN(n456) );
  INV_X1 U517 ( .A(KEYINPUT124), .ZN(n455) );
  NAND2_X1 U518 ( .A1(n481), .A2(n582), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n458) );
  XOR2_X1 U520 ( .A(n503), .B(KEYINPUT27), .Z(n471) );
  XNOR2_X1 U521 ( .A(n461), .B(KEYINPUT97), .ZN(n468) );
  INV_X1 U522 ( .A(KEYINPUT98), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT25), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n522), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT99), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n522), .A2(n471), .ZN(n472) );
  XNOR2_X1 U530 ( .A(KEYINPUT96), .B(n472), .ZN(n550) );
  XOR2_X1 U531 ( .A(n473), .B(KEYINPUT28), .Z(n531) );
  NAND2_X1 U532 ( .A1(n550), .A2(n531), .ZN(n536) );
  NOR2_X1 U533 ( .A1(n534), .A2(n536), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT100), .ZN(n489) );
  NOR2_X1 U536 ( .A1(n489), .A2(n579), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(KEYINPUT102), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n478), .A2(n583), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n479), .B(KEYINPUT103), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT37), .B(n480), .Z(n521) );
  NOR2_X1 U541 ( .A1(n566), .A2(n481), .ZN(n491) );
  NAND2_X1 U542 ( .A1(n521), .A2(n491), .ZN(n483) );
  XOR2_X1 U543 ( .A(KEYINPUT38), .B(KEYINPUT104), .Z(n482) );
  XNOR2_X2 U544 ( .A(n483), .B(n482), .ZN(n508) );
  NAND2_X1 U545 ( .A1(n508), .A2(n534), .ZN(n486) );
  XOR2_X1 U546 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n484) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n488) );
  NAND2_X1 U548 ( .A1(n579), .A2(n546), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n490) );
  NOR2_X1 U550 ( .A1(n490), .A2(n489), .ZN(n512) );
  NAND2_X1 U551 ( .A1(n512), .A2(n491), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT101), .ZN(n498) );
  NAND2_X1 U553 ( .A1(n498), .A2(n500), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(KEYINPUT34), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NAND2_X1 U556 ( .A1(n503), .A2(n498), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .Z(n497) );
  NAND2_X1 U559 ( .A1(n498), .A2(n534), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(G1326GAT) );
  INV_X1 U561 ( .A(n531), .ZN(n507) );
  NAND2_X1 U562 ( .A1(n498), .A2(n507), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .Z(n502) );
  NAND2_X1 U565 ( .A1(n508), .A2(n500), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n505) );
  NAND2_X1 U568 ( .A1(n508), .A2(n503), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  INV_X1 U574 ( .A(n556), .ZN(n568) );
  NOR2_X1 U575 ( .A1(n575), .A2(n568), .ZN(n511) );
  XOR2_X1 U576 ( .A(KEYINPUT109), .B(n511), .Z(n520) );
  NAND2_X1 U577 ( .A1(n520), .A2(n512), .ZN(n517) );
  NOR2_X1 U578 ( .A1(n522), .A2(n517), .ZN(n513) );
  XOR2_X1 U579 ( .A(G57GAT), .B(n513), .Z(n514) );
  XNOR2_X1 U580 ( .A(KEYINPUT42), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n525), .A2(n517), .ZN(n515) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n527), .A2(n517), .ZN(n516) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n531), .A2(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n522), .A2(n530), .ZN(n523) );
  XOR2_X1 U590 ( .A(KEYINPUT110), .B(n523), .Z(n524) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n530), .ZN(n526) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n527), .A2(n530), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(G1338GAT) );
  NOR2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(n532), .Z(n533) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U600 ( .A1(n551), .A2(n534), .ZN(n535) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n575), .A2(n542), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT116), .Z(n539) );
  NAND2_X1 U605 ( .A1(n542), .A2(n556), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  INV_X1 U609 ( .A(n542), .ZN(n545) );
  NOR2_X1 U610 ( .A1(n573), .A2(n545), .ZN(n543) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n564), .A2(n575), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1344GAT) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n558) );
  NAND2_X1 U624 ( .A1(n564), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  XOR2_X1 U627 ( .A(G155GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U628 ( .A1(n564), .A2(n579), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(n565), .ZN(G1347GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n572), .ZN(n567) );
  XOR2_X1 U633 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  NOR2_X1 U634 ( .A1(n572), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(n571), .ZN(G1349GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  AND2_X1 U641 ( .A1(n575), .A2(n582), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  NAND2_X1 U644 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n585) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

