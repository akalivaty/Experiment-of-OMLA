//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT65), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  NAND2_X1  g0051(.A1(new_n208), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n216), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(new_n207), .A3(G1), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n206), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G68), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT12), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n255), .B2(new_n220), .ZN(new_n260));
  INV_X1    g0060(.A(new_n255), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(KEYINPUT12), .A3(G68), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT71), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n207), .A2(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n226), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n253), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT70), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n271), .A2(KEYINPUT11), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(KEYINPUT11), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n263), .A2(new_n264), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n265), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT14), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  OR2_X1    g0084(.A1(new_n284), .A2(G232), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n283), .B(new_n285), .C1(G226), .C2(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n278), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT13), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n277), .A2(KEYINPUT66), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  AOI21_X1  g0094(.A(G1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n277), .A2(KEYINPUT66), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n292), .A2(G274), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n295), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n292), .A2(G238), .A3(new_n298), .A4(new_n296), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n290), .A2(new_n291), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n291), .B1(new_n290), .B2(new_n300), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n276), .B(G169), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n303), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(G179), .A3(new_n301), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n301), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n276), .B1(new_n308), .B2(G169), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n275), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n275), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n305), .B2(new_n301), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n284), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(G223), .B1(G77), .B2(new_n321), .ZN(new_n323));
  INV_X1    g0123(.A(G222), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n283), .A2(new_n284), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n277), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n292), .A2(new_n298), .A3(new_n296), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G226), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n297), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT67), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n327), .A2(KEYINPUT67), .A3(new_n297), .A4(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(G169), .ZN(new_n335));
  INV_X1    g0135(.A(new_n216), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n208), .B2(G33), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT8), .B(G58), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n268), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n339), .A2(new_n340), .B1(G150), .B2(new_n266), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n203), .A2(G20), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n337), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT68), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n256), .A2(G50), .A3(new_n257), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(new_n345), .C1(G50), .C2(new_n261), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n343), .A2(KEYINPUT68), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(G179), .B1(new_n332), .B2(new_n333), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n335), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n334), .A2(G190), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n332), .A2(G200), .A3(new_n333), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(KEYINPUT9), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT9), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n346), .B2(new_n347), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT10), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n354), .A2(new_n356), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT10), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n351), .A4(new_n353), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n350), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n321), .A2(G1698), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G232), .B1(G107), .B2(new_n321), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n283), .A2(G1698), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n221), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n277), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n328), .A2(G244), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n297), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G200), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n256), .A2(G77), .A3(new_n257), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(G77), .B2(new_n261), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n339), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n373));
  XOR2_X1   g0173(.A(KEYINPUT15), .B(G87), .Z(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n373), .B1(new_n268), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n253), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n370), .B(new_n377), .C1(new_n313), .C2(new_n369), .ZN(new_n378));
  INV_X1    g0178(.A(G169), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n369), .B2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n369), .A2(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n318), .A2(new_n362), .A3(new_n378), .A4(new_n382), .ZN(new_n383));
  MUX2_X1   g0183(.A(G223), .B(G226), .S(G1698), .Z(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n283), .B1(G33), .B2(G87), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n385), .A2(new_n278), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n292), .A2(G232), .A3(new_n298), .A4(new_n296), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(new_n297), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n379), .ZN(new_n389));
  INV_X1    g0189(.A(G179), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n386), .A2(new_n387), .A3(new_n297), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n283), .B2(G20), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n321), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n220), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  INV_X1    g0199(.A(G58), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n220), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n201), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n266), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OR3_X1    g0204(.A1(new_n398), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n399), .B1(new_n398), .B2(new_n404), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n253), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n338), .B1(new_n206), .B2(G20), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n256), .A2(new_n408), .B1(new_n255), .B2(new_n338), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n389), .A2(KEYINPUT72), .A3(new_n391), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n394), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT73), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n392), .A2(new_n393), .B1(new_n407), .B2(new_n409), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT18), .A4(new_n411), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n413), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n388), .A2(new_n313), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n388), .A2(G200), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n420), .A2(new_n407), .A3(new_n409), .A4(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n383), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n206), .A2(G33), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n256), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n337), .A2(new_n261), .A3(new_n427), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT75), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(G107), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n255), .A2(new_n228), .ZN(new_n432));
  XOR2_X1   g0232(.A(new_n432), .B(KEYINPUT25), .Z(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n206), .A2(G45), .ZN(new_n435));
  OR2_X1    g0235(.A1(KEYINPUT5), .A2(G41), .ZN(new_n436));
  NAND2_X1  g0236(.A1(KEYINPUT5), .A2(G41), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n292), .A2(G274), .A3(new_n296), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n438), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n292), .A2(G264), .A3(new_n296), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G294), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n325), .B2(new_n223), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT87), .ZN(new_n444));
  INV_X1    g0244(.A(G257), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n365), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n322), .A2(KEYINPUT87), .A3(G257), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n439), .B(new_n441), .C1(new_n448), .C2(new_n278), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n315), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n363), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT87), .B1(new_n322), .B2(G257), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n365), .A2(new_n444), .A3(new_n445), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n277), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(new_n313), .A3(new_n439), .A4(new_n441), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n207), .A2(G87), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n281), .B2(new_n282), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT82), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n222), .A2(G20), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n319), .B2(new_n320), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT22), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n467), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n283), .A2(new_n472), .A3(KEYINPUT84), .A4(new_n462), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT85), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT85), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n466), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT23), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n207), .B2(G107), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n228), .A2(KEYINPUT23), .A3(G20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g0283(.A(KEYINPUT78), .B(G116), .Z(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G33), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(G20), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT86), .B1(new_n479), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n337), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n478), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n477), .B1(new_n466), .B2(new_n474), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT86), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(KEYINPUT86), .B(new_n487), .C1(new_n491), .C2(new_n492), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(KEYINPUT24), .A3(new_n496), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n434), .B(new_n457), .C1(new_n490), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n449), .A2(new_n379), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G179), .B2(new_n449), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n493), .A2(new_n494), .A3(new_n489), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n486), .B1(new_n476), .B2(new_n478), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT24), .B1(new_n502), .B2(KEYINPUT86), .ZN(new_n503));
  INV_X1    g0303(.A(new_n496), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n253), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n434), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n292), .A2(G257), .A3(new_n296), .A4(new_n440), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n439), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n363), .B(G244), .C1(KEYINPUT76), .C2(KEYINPUT4), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n325), .B2(new_n227), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n322), .A2(G250), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n511), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n516), .B2(new_n277), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G200), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n228), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  XOR2_X1   g0320(.A(G97), .B(G107), .Z(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(KEYINPUT6), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n396), .A2(new_n397), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n228), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n253), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n428), .A2(G97), .A3(new_n430), .ZN(new_n527));
  INV_X1    g0327(.A(G97), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n255), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g0329(.A(new_n529), .B(KEYINPUT74), .Z(new_n530));
  AND2_X1   g0330(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n517), .A2(G190), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n519), .A2(new_n526), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n526), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n517), .A2(new_n390), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n535), .C1(G169), .C2(new_n517), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n207), .B1(new_n287), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n222), .A2(new_n528), .A3(new_n228), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g0340(.A(new_n540), .B(KEYINPUT79), .Z(new_n541));
  NAND3_X1  g0341(.A1(new_n283), .A2(new_n207), .A3(G68), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n537), .B1(new_n268), .B2(new_n528), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n253), .B1(new_n255), .B2(new_n375), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n428), .A2(new_n374), .A3(new_n430), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI221_X1 g0347(.A(new_n485), .B1(new_n325), .B2(new_n221), .C1(new_n227), .C2(new_n365), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n277), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n292), .A2(new_n296), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT77), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n435), .A2(new_n551), .A3(G250), .ZN(new_n552));
  AOI21_X1  g0352(.A(G274), .B1(KEYINPUT77), .B2(G250), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n435), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n379), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n548), .A2(new_n277), .B1(new_n550), .B2(new_n554), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n390), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n547), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n556), .A2(G200), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n428), .A2(G87), .A3(new_n430), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n558), .A2(G190), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n561), .A2(new_n545), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n533), .A2(new_n536), .A3(new_n560), .A4(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n292), .A2(G270), .A3(new_n296), .A4(new_n440), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n439), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n283), .A2(G257), .A3(new_n284), .ZN(new_n568));
  XOR2_X1   g0368(.A(KEYINPUT80), .B(G303), .Z(new_n569));
  OAI221_X1 g0369(.A(new_n568), .B1(new_n569), .B2(new_n283), .C1(new_n365), .C2(new_n229), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n277), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n379), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n429), .A2(new_n573), .B1(new_n261), .B2(new_n484), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n514), .B(new_n207), .C1(G33), .C2(new_n528), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n253), .B(new_n576), .C1(new_n207), .C2(new_n484), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT20), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n572), .A2(KEYINPUT21), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT81), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT81), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n572), .A2(new_n581), .A3(new_n584), .A4(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n581), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n567), .A2(G179), .A3(new_n571), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT21), .B1(new_n572), .B2(new_n581), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n567), .A2(new_n571), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n581), .B1(G200), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n313), .B2(new_n592), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n586), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n565), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n425), .A2(new_n508), .A3(new_n596), .ZN(G372));
  XNOR2_X1  g0397(.A(new_n412), .B(KEYINPUT18), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n317), .ZN(new_n600));
  INV_X1    g0400(.A(new_n382), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n311), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n423), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n358), .A2(new_n361), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n350), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n425), .ZN(new_n607));
  INV_X1    g0407(.A(new_n507), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n586), .A2(new_n591), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT88), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(KEYINPUT88), .A3(new_n609), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n498), .A2(new_n565), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n560), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n560), .A2(new_n564), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  OR3_X1    g0418(.A1(new_n617), .A2(new_n536), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n617), .B2(new_n536), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n606), .B1(new_n607), .B2(new_n623), .ZN(G369));
  AOI21_X1  g0424(.A(new_n434), .B1(new_n490), .B2(new_n497), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G343), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT89), .B1(new_n625), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n505), .A2(new_n506), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT89), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n631), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n609), .A2(new_n631), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n508), .A2(new_n633), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT90), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n507), .A2(new_n632), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n639), .B1(new_n638), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n508), .A2(new_n633), .A3(new_n636), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n507), .A2(new_n631), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n609), .A2(new_n587), .A3(new_n632), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n587), .A2(new_n632), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n595), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G330), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n643), .A2(new_n652), .ZN(G399));
  INV_X1    g0453(.A(new_n210), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n539), .A2(G116), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n657), .B(KEYINPUT91), .Z(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n658), .A3(G1), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n214), .B2(new_n656), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT92), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT28), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n610), .A2(new_n614), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n631), .B1(new_n663), .B2(new_n621), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT29), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT95), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(KEYINPUT95), .A3(KEYINPUT29), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n631), .B1(new_n615), .B2(new_n621), .ZN(new_n669));
  XNOR2_X1  g0469(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n667), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n517), .A2(new_n441), .A3(new_n455), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n558), .A2(G179), .A3(new_n571), .A4(new_n567), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n588), .A2(new_n556), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n455), .A2(new_n441), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(KEYINPUT30), .A3(new_n677), .A4(new_n517), .ZN(new_n678));
  AOI21_X1  g0478(.A(G179), .B1(new_n567), .B2(new_n571), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n518), .A2(new_n679), .A3(new_n449), .A4(new_n556), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n675), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(KEYINPUT31), .A3(new_n631), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT93), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n631), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT31), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n508), .A2(new_n596), .A3(new_n632), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n671), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n662), .B1(new_n695), .B2(G1), .ZN(G364));
  NOR2_X1   g0496(.A1(new_n254), .A2(G20), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n206), .B1(new_n697), .B2(G45), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n655), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n650), .B2(G330), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(G330), .B2(new_n650), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n210), .A2(new_n283), .ZN(new_n703));
  INV_X1    g0503(.A(G355), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n703), .A2(new_n704), .B1(G116), .B2(new_n210), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n654), .A2(new_n283), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n294), .B2(new_n215), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n250), .A2(G45), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G13), .A2(G33), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n216), .B1(G20), .B2(new_n379), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n700), .B1(new_n710), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n207), .A2(new_n390), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G190), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n315), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n202), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT32), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n207), .A2(G190), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G179), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G159), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n724), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n729), .A2(new_n390), .A3(new_n315), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n283), .B1(new_n723), .B2(new_n728), .C1(new_n731), .C2(new_n220), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n722), .B(new_n732), .C1(new_n723), .C2(new_n728), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n390), .A2(G200), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT98), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n729), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT99), .Z(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G107), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n718), .A2(new_n313), .A3(new_n315), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT97), .Z(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n736), .A2(new_n207), .A3(new_n313), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n742), .A2(G77), .B1(new_n743), .B2(G87), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n719), .A2(G200), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT96), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n207), .B1(new_n725), .B2(G190), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT100), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n751), .A2(G58), .B1(G97), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n733), .A2(new_n739), .A3(new_n744), .A4(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n751), .A2(G322), .B1(G294), .B2(new_n756), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n738), .A2(G283), .ZN(new_n760));
  INV_X1    g0560(.A(G311), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT33), .B(G317), .Z(new_n762));
  OAI221_X1 g0562(.A(new_n321), .B1(new_n761), .B2(new_n740), .C1(new_n731), .C2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G326), .B2(new_n720), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n726), .B(KEYINPUT101), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n743), .A2(G303), .B1(new_n765), .B2(G329), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n759), .A2(new_n760), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n717), .B1(new_n768), .B2(new_n714), .ZN(new_n769));
  INV_X1    g0569(.A(new_n713), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n650), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n702), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(G396));
  NOR2_X1   g0573(.A1(new_n382), .A2(new_n631), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n378), .B1(new_n377), .B2(new_n632), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(new_n775), .B2(new_n382), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n669), .B(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n700), .B1(new_n777), .B2(new_n693), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n693), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n714), .A2(new_n711), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n700), .B1(G77), .B2(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G150), .A2(new_n730), .B1(new_n720), .B2(G137), .ZN(new_n783));
  INV_X1    g0583(.A(G143), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n783), .B1(new_n727), .B2(new_n741), .C1(new_n750), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT34), .Z(new_n786));
  INV_X1    g0586(.A(new_n743), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n283), .B1(new_n787), .B2(new_n202), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G132), .B2(new_n765), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n738), .A2(G68), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n789), .B(new_n790), .C1(new_n400), .C2(new_n755), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n730), .B(KEYINPUT102), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n283), .B(new_n794), .C1(G303), .C2(new_n720), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n738), .A2(G87), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n765), .A2(G311), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n742), .A2(new_n484), .B1(new_n743), .B2(G107), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G294), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n750), .A2(new_n800), .B1(new_n528), .B2(new_n755), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT103), .Z(new_n802));
  OAI22_X1  g0602(.A1(new_n786), .A2(new_n791), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n782), .B1(new_n803), .B2(new_n714), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n776), .B2(new_n712), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n779), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT104), .ZN(G384));
  NOR2_X1   g0607(.A1(new_n697), .A2(new_n206), .ZN(new_n808));
  INV_X1    g0608(.A(G330), .ZN(new_n809));
  INV_X1    g0609(.A(new_n776), .ZN(new_n810));
  INV_X1    g0610(.A(new_n307), .ZN(new_n811));
  INV_X1    g0611(.A(new_n309), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n275), .B(new_n631), .C1(new_n813), .C2(new_n317), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n275), .A2(new_n631), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n600), .A2(new_n310), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n810), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n691), .A2(new_n682), .A3(new_n687), .ZN(new_n818));
  INV_X1    g0618(.A(new_n629), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n410), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n419), .B2(new_n423), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n412), .A2(new_n422), .A3(new_n820), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT37), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n822), .B(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT38), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n820), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n598), .B2(new_n603), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n822), .B(KEYINPUT37), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT38), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n817), .B(new_n818), .C1(new_n826), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT40), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n424), .A2(new_n827), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n833), .A2(KEYINPUT38), .A3(new_n829), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n825), .B1(new_n821), .B2(new_n824), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT40), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(new_n818), .A4(new_n817), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n425), .A2(new_n818), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n809), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT106), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n669), .A2(new_n776), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n774), .B(KEYINPUT105), .Z(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n814), .A2(new_n816), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n849), .A3(new_n836), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n834), .A2(KEYINPUT39), .A3(new_n835), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n311), .A2(new_n632), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n826), .A2(new_n830), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n851), .B(new_n853), .C1(new_n854), .C2(KEYINPUT39), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n598), .A2(new_n629), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n606), .B1(new_n671), .B2(new_n607), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n859), .B(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n808), .B1(new_n844), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n844), .B2(new_n861), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n864), .A2(G116), .A3(new_n217), .A4(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n214), .A2(new_n226), .A3(new_n401), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n220), .A2(G50), .ZN(new_n869));
  OAI211_X1 g0669(.A(G1), .B(new_n254), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n863), .A2(new_n867), .A3(new_n870), .ZN(G367));
  OR2_X1    g0671(.A1(new_n536), .A2(new_n632), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n534), .A2(new_n631), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n533), .A2(new_n536), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n638), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT42), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n608), .A2(new_n874), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n631), .B1(new_n879), .B2(new_n536), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n877), .B2(KEYINPUT42), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n545), .A2(new_n562), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n631), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n560), .A2(new_n564), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n560), .B2(new_n883), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n878), .A2(new_n881), .B1(KEYINPUT43), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(KEYINPUT43), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n652), .A2(new_n875), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n888), .B(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n655), .B(KEYINPUT41), .Z(new_n891));
  XOR2_X1   g0691(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT108), .B1(new_n643), .B2(new_n876), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT108), .ZN(new_n894));
  NOR4_X1   g0694(.A1(new_n641), .A2(new_n642), .A3(new_n894), .A4(new_n875), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n643), .A2(KEYINPUT108), .A3(new_n876), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n638), .A2(new_n640), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT90), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(new_n876), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n894), .ZN(new_n902));
  INV_X1    g0702(.A(new_n892), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n897), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT45), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n643), .B2(new_n876), .ZN(new_n906));
  OAI211_X1 g0706(.A(KEYINPUT45), .B(new_n875), .C1(new_n641), .C2(new_n642), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n896), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n652), .ZN(new_n910));
  INV_X1    g0710(.A(new_n652), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n896), .A2(new_n911), .A3(new_n904), .A4(new_n908), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n638), .B1(new_n646), .B2(new_n637), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(KEYINPUT109), .B2(new_n651), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n651), .B(KEYINPUT109), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n916), .B2(new_n913), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n694), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n912), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n891), .B1(new_n919), .B2(new_n695), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n890), .B1(new_n920), .B2(new_n699), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT110), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT110), .B(new_n890), .C1(new_n920), .C2(new_n699), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n737), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n741), .A2(new_n202), .B1(new_n926), .B2(new_n226), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(G58), .B2(new_n743), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n756), .A2(G68), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n751), .A2(G150), .ZN(new_n930));
  INV_X1    g0730(.A(G137), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n283), .B1(new_n726), .B2(new_n931), .C1(new_n721), .C2(new_n784), .ZN(new_n932));
  INV_X1    g0732(.A(new_n792), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n932), .B1(new_n933), .B2(G159), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n742), .A2(G283), .B1(new_n756), .B2(G107), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(G317), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n321), .B1(new_n726), .B2(new_n939), .C1(new_n721), .C2(new_n761), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G97), .B2(new_n737), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT46), .B1(new_n743), .B2(new_n484), .ZN(new_n942));
  INV_X1    g0742(.A(new_n569), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n751), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(KEYINPUT46), .A2(G116), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n933), .A2(G294), .B1(new_n743), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n938), .A2(new_n941), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n936), .A2(new_n937), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n935), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT112), .Z(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT47), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT47), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n714), .A3(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n700), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n237), .A2(new_n707), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n716), .B1(new_n654), .B2(new_n374), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n953), .B(new_n957), .C1(new_n770), .C2(new_n885), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT113), .Z(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n925), .A2(new_n960), .ZN(G387));
  INV_X1    g0761(.A(new_n917), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n647), .A2(new_n713), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n706), .B1(new_n241), .B2(new_n294), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n658), .B2(new_n703), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n966));
  OR3_X1    g0766(.A1(new_n966), .A2(G50), .A3(new_n338), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n966), .B1(G50), .B2(new_n338), .ZN(new_n968));
  AOI21_X1  g0768(.A(G45), .B1(G68), .B2(G77), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n658), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n965), .A2(new_n970), .B1(new_n228), .B2(new_n654), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n700), .B1(new_n971), .B2(new_n716), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n738), .A2(G97), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n283), .B1(new_n740), .B2(new_n220), .ZN(new_n974));
  INV_X1    g0774(.A(G150), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n731), .A2(new_n338), .B1(new_n726), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(G159), .C2(new_n720), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n755), .A2(new_n375), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n751), .B2(G50), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n743), .A2(G77), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n973), .A2(new_n977), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(KEYINPUT115), .B(G322), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n792), .A2(new_n761), .B1(new_n721), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT116), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(KEYINPUT116), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n751), .A2(G317), .B1(new_n943), .B2(new_n742), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT48), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n787), .A2(new_n800), .B1(new_n793), .B2(new_n755), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n987), .B2(new_n988), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n737), .A2(new_n484), .ZN(new_n993));
  INV_X1    g0793(.A(new_n726), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n283), .B1(new_n994), .B2(G326), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT49), .B1(new_n989), .B2(new_n991), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n981), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n972), .B1(new_n998), .B2(new_n714), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n962), .A2(new_n699), .B1(new_n963), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n918), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n655), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n962), .A2(new_n695), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(G393));
  NAND3_X1  g0804(.A1(new_n910), .A2(new_n699), .A3(new_n912), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n715), .B1(new_n528), .B2(new_n210), .C1(new_n707), .C2(new_n245), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n700), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n283), .B1(new_n726), .B2(new_n784), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n787), .A2(new_n220), .B1(new_n741), .B2(new_n338), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G50), .C2(new_n933), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n796), .C1(new_n226), .C2(new_n755), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n750), .A2(new_n727), .B1(new_n975), .B2(new_n721), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT51), .Z(new_n1013));
  OAI22_X1  g0813(.A1(new_n750), .A2(new_n761), .B1(new_n939), .B2(new_n721), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT52), .Z(new_n1015));
  OAI221_X1 g0815(.A(new_n321), .B1(new_n726), .B2(new_n982), .C1(new_n740), .C2(new_n800), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n787), .A2(new_n793), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n943), .C2(new_n933), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n756), .A2(new_n484), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n739), .A3(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1011), .A2(new_n1013), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1007), .B1(new_n1021), .B2(new_n714), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n875), .B2(new_n770), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1005), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n919), .A2(new_n655), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n910), .A2(new_n912), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n1001), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(G390));
  AOI21_X1  g0829(.A(new_n846), .B1(new_n669), .B2(new_n776), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n849), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n852), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n851), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT117), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n664), .A2(new_n776), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1031), .B1(new_n1036), .B2(new_n847), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n852), .B1(new_n826), .B2(new_n830), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1035), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1038), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n846), .B1(new_n664), .B2(new_n776), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(KEYINPUT117), .C1(new_n1041), .C2(new_n1031), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n692), .A2(G330), .A3(new_n776), .A4(new_n849), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1034), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1032), .A2(new_n1033), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n817), .A2(G330), .A3(new_n818), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1045), .B(new_n699), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1033), .A2(new_n711), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n700), .B1(new_n339), .B2(new_n781), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n755), .A2(new_n226), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n321), .B1(new_n721), .B2(new_n793), .C1(new_n787), .C2(new_n222), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G116), .C2(new_n751), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n765), .A2(G294), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n933), .A2(G107), .B1(new_n742), .B2(G97), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1053), .A2(new_n790), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n743), .A2(G150), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT53), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n933), .A2(G137), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT54), .B(G143), .Z(new_n1060));
  AOI22_X1  g0860(.A1(new_n742), .A2(new_n1060), .B1(G128), .B2(new_n720), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n751), .A2(G132), .B1(G159), .B2(new_n756), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n765), .ZN(new_n1064));
  INV_X1    g0864(.A(G125), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n283), .B1(new_n926), .B2(new_n202), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT118), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1056), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1050), .B1(new_n1068), .B2(new_n714), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1049), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1048), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n818), .A2(G330), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n425), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n606), .B(new_n1074), .C1(new_n671), .C2(new_n607), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n776), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1031), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1044), .A2(new_n1041), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n809), .B(new_n810), .C1(new_n690), .C2(new_n691), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1047), .B1(new_n1080), .B2(new_n849), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1078), .A2(new_n1079), .B1(new_n848), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1076), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n656), .B1(new_n1072), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1086), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1071), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(G378));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1076), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n819), .B1(new_n346), .B2(new_n347), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT119), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n362), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n362), .A2(new_n1094), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1092), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n362), .A2(new_n1094), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1092), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n1095), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n817), .A2(new_n837), .A3(new_n818), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1103), .A2(new_n836), .B1(new_n831), .B2(KEYINPUT40), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(new_n809), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1102), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n839), .A2(G330), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT122), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n836), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1030), .A2(new_n1031), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1111), .B2(new_n857), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n850), .A2(new_n858), .A3(KEYINPUT122), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1108), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n859), .A2(new_n1105), .A3(new_n1109), .A4(new_n1107), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1114), .A2(KEYINPUT57), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1090), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT120), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1106), .B1(new_n839), .B2(G330), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n809), .B(new_n1102), .C1(new_n832), .C2(new_n838), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n859), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n859), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1087), .A2(new_n1076), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1117), .B(new_n655), .C1(KEYINPUT57), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT121), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n698), .B1(new_n1124), .B2(new_n1121), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1102), .A2(new_n711), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n730), .A2(G132), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n931), .B2(new_n740), .C1(new_n721), .C2(new_n1065), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n743), .B2(new_n1060), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n750), .C1(new_n975), .C2(new_n755), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n737), .A2(G159), .ZN(new_n1137));
  AOI211_X1 g0937(.A(G33), .B(G41), .C1(new_n994), .C2(G124), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n980), .B1(new_n926), .B2(new_n400), .C1(new_n1064), .C2(new_n793), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n321), .A2(new_n293), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n375), .A2(new_n740), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(G97), .C2(new_n730), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n720), .A2(G116), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n929), .A3(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1140), .B(new_n1145), .C1(G107), .C2(new_n751), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT58), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1141), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1146), .A2(KEYINPUT58), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1139), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n714), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n954), .B1(new_n202), .B2(new_n780), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1129), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1127), .B1(new_n1128), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1121), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n859), .B1(new_n1108), .B2(new_n1118), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n699), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(KEYINPUT121), .A3(new_n1153), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1126), .A2(new_n1160), .ZN(G375));
  INV_X1    g0961(.A(new_n891), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1084), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1031), .A2(new_n711), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n700), .B1(G68), .B2(new_n781), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n933), .A2(new_n484), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n228), .B2(new_n741), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G97), .B2(new_n743), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n751), .A2(G283), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n321), .B1(new_n721), .B2(new_n800), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n978), .C1(G303), .C2(new_n765), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n738), .A2(G77), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n933), .A2(new_n1060), .B1(G132), .B2(new_n720), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n750), .B2(new_n931), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT123), .Z(new_n1177));
  OAI221_X1 g0977(.A(new_n283), .B1(new_n975), .B2(new_n740), .C1(new_n926), .C2(new_n400), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n787), .A2(new_n727), .B1(new_n1064), .B2(new_n1133), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n202), .B2(new_n755), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1174), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1166), .B1(new_n1182), .B2(new_n714), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1083), .A2(new_n699), .B1(new_n1165), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1164), .A2(new_n1184), .ZN(G381));
  XOR2_X1   g0985(.A(G375), .B(KEYINPUT124), .Z(new_n1186));
  AOI21_X1  g0986(.A(new_n959), .B1(new_n923), .B2(new_n924), .ZN(new_n1187));
  OR2_X1    g0987(.A1(G393), .A2(G396), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(G378), .A2(new_n1188), .A3(G384), .A4(G381), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1028), .A4(new_n1189), .ZN(G407));
  NAND4_X1  g0990(.A1(new_n1186), .A2(G213), .A3(new_n630), .A4(new_n1088), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(G407), .A2(new_n1191), .A3(G213), .ZN(G409));
  INV_X1    g0992(.A(KEYINPUT126), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1187), .B2(G390), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(G393), .B(new_n772), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G390), .B1(new_n925), .B2(new_n960), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n959), .B(new_n1028), .C1(new_n923), .C2(new_n924), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n1194), .A2(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(G387), .A2(new_n1028), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1187), .A2(G390), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1195), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1199), .A2(new_n1193), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1126), .A2(G378), .A3(new_n1160), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1125), .A2(new_n1162), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1114), .A2(new_n699), .A3(new_n1115), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1153), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1088), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n630), .A2(G213), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1084), .A2(KEYINPUT60), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1211), .A2(new_n1163), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n655), .B1(new_n1211), .B2(new_n1163), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1184), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(G384), .ZN(new_n1215));
  AND4_X1   g1015(.A1(KEYINPUT62), .A2(new_n1209), .A3(new_n1210), .A4(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1209), .A2(KEYINPUT125), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1204), .A2(new_n1208), .A3(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1217), .A2(new_n1210), .A3(new_n1215), .A4(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT62), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1216), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT61), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n630), .A2(G213), .A3(G2897), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1215), .B(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1203), .B1(new_n1222), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT63), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1220), .A2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1215), .A2(KEYINPUT63), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT61), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1217), .A2(new_n1210), .A3(new_n1219), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1230), .B(new_n1232), .C1(new_n1233), .C2(new_n1225), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1228), .B1(new_n1234), .B2(new_n1203), .ZN(G405));
  INV_X1    g1035(.A(new_n1204), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G378), .B1(new_n1126), .B2(new_n1160), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1238), .A2(new_n1215), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1215), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1198), .A2(new_n1202), .A3(KEYINPUT127), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT127), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT127), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1198), .A2(new_n1202), .A3(KEYINPUT127), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1241), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(new_n1250), .ZN(G402));
endmodule


