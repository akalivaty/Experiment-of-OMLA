//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT78), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT29), .ZN(new_n208));
  XOR2_X1   g007(.A(G141gat), .B(G148gat), .Z(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n212), .C1(new_n217), .C2(KEYINPUT2), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n208), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n220));
  XNOR2_X1  g019(.A(G197gat), .B(G204gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222));
  INV_X1    g021(.A(G211gat), .ZN(new_n223));
  INV_X1    g022(.A(G218gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n220), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT78), .B1(new_n202), .B2(new_n203), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n216), .A2(new_n218), .ZN(new_n232));
  INV_X1    g031(.A(new_n227), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n226), .B(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n208), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n207), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n228), .A2(KEYINPUT29), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n219), .B1(new_n239), .B2(KEYINPUT3), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n240), .A2(new_n206), .A3(new_n230), .A4(new_n229), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT79), .B(G22gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n238), .B2(new_n241), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n238), .A2(new_n241), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT80), .A3(new_n243), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT31), .B(G50gat), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n251), .B(new_n252), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n245), .A2(new_n253), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(G22gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n219), .B(new_n236), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  INV_X1    g061(.A(G120gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(G113gat), .B2(G120gat), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT69), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n268), .B(KEYINPUT69), .C1(new_n264), .C2(new_n266), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT74), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n260), .B1(new_n261), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n271), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n232), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT4), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n232), .A2(new_n280), .A3(new_n277), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT5), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(KEYINPUT75), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n232), .A2(new_n285), .A3(new_n277), .A4(new_n280), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n286), .A3(new_n279), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n276), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n277), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(new_n219), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n275), .B2(new_n219), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT5), .B1(new_n291), .B2(new_n259), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n283), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G1gat), .B(G29gat), .Z(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G57gat), .B(G85gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n283), .B(new_n298), .C1(new_n288), .C2(new_n292), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(new_n272), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n278), .B1(new_n306), .B2(new_n232), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n307), .B2(new_n260), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n276), .A2(new_n287), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n308), .A2(new_n309), .B1(new_n276), .B2(new_n282), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n310), .A2(new_n301), .A3(new_n298), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G8gat), .B(G36gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT66), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n321), .A2(new_n327), .A3(new_n324), .A4(new_n322), .ZN(new_n328));
  INV_X1    g127(.A(G183gat), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT64), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT64), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n333), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n326), .B(new_n328), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n331), .A2(new_n332), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n336), .A2(new_n337), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n339), .A2(KEYINPUT64), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n344), .B(new_n342), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n319), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  AOI211_X1 g148(.A(new_n319), .B(new_n325), .C1(new_n344), .C2(new_n336), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n320), .A2(KEYINPUT26), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n334), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n322), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(new_n320), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n329), .A2(KEYINPUT27), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G183gat), .ZN(new_n361));
  AND4_X1   g160(.A1(KEYINPUT28), .A2(new_n359), .A3(new_n361), .A4(new_n330), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT67), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n360), .B2(G183gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT27), .B(G183gat), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n330), .B(new_n364), .C1(new_n365), .C2(new_n363), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n358), .B1(new_n368), .B2(KEYINPUT68), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n359), .B2(new_n361), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n330), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n362), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT68), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n349), .A2(new_n351), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n318), .B1(new_n376), .B2(KEYINPUT29), .ZN(new_n377));
  INV_X1    g176(.A(new_n318), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT65), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n380), .A2(new_n347), .A3(new_n326), .A4(new_n328), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n350), .B1(new_n381), .B2(new_n319), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT68), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n357), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(new_n374), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n378), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n377), .A2(new_n234), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT72), .B1(new_n376), .B2(new_n318), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT72), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n378), .C1(new_n382), .C2(new_n385), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n208), .B1(new_n382), .B2(new_n385), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n388), .A2(new_n390), .B1(new_n318), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT73), .B(new_n387), .C1(new_n392), .C2(new_n234), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n377), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n228), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n317), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n313), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n393), .A2(new_n397), .A3(new_n317), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n317), .A2(KEYINPUT37), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n234), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n228), .A3(new_n386), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n403), .A2(KEYINPUT83), .A3(KEYINPUT37), .A4(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n392), .A2(new_n228), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(KEYINPUT37), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT38), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n399), .B1(new_n402), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n401), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n393), .A2(new_n397), .A3(KEYINPUT37), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n258), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n261), .A2(new_n275), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n279), .A2(new_n281), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n259), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT39), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n307), .A2(new_n260), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n298), .B(new_n421), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT40), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n300), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n421), .A2(new_n298), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n419), .A2(new_n423), .A3(new_n420), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n429), .A2(KEYINPUT81), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(KEYINPUT81), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n234), .B1(new_n394), .B2(new_n377), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n387), .A2(KEYINPUT73), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n392), .A2(KEYINPUT73), .A3(new_n234), .ZN(new_n436));
  OAI211_X1 g235(.A(KEYINPUT30), .B(new_n316), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n400), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n398), .A2(KEYINPUT30), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT82), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n432), .B(new_n442), .C1(new_n438), .C2(new_n439), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n416), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n316), .B1(new_n435), .B2(new_n436), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n447), .A2(new_n313), .A3(new_n400), .A4(new_n437), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT77), .ZN(new_n449));
  INV_X1    g248(.A(new_n258), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n393), .A2(new_n397), .A3(new_n317), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(KEYINPUT30), .B2(new_n398), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT77), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n313), .A4(new_n447), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT36), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n277), .B1(new_n382), .B2(new_n385), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n349), .A2(new_n351), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n369), .A2(new_n375), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n289), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(G71gat), .B(G99gat), .Z(new_n464));
  XNOR2_X1  g263(.A(G15gat), .B(G43gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT33), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(KEYINPUT32), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n463), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n461), .B2(KEYINPUT71), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n461), .ZN(new_n477));
  AOI211_X1 g276(.A(new_n462), .B(new_n474), .C1(new_n457), .C2(new_n460), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n463), .A2(KEYINPUT32), .ZN(new_n480));
  INV_X1    g279(.A(new_n463), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n480), .B(new_n466), .C1(new_n481), .C2(KEYINPUT33), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n472), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n479), .B1(new_n472), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n456), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n472), .A2(new_n482), .ZN(new_n486));
  INV_X1    g285(.A(new_n479), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n479), .A3(new_n482), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT36), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n455), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n444), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(new_n258), .A3(new_n489), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n448), .A2(KEYINPUT35), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n488), .A2(new_n258), .A3(KEYINPUT84), .A4(new_n489), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n438), .A2(new_n439), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n453), .B1(new_n500), .B2(new_n313), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n448), .A2(KEYINPUT77), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n495), .B1(new_n503), .B2(KEYINPUT35), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT85), .B1(new_n493), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n495), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n449), .A2(new_n454), .B1(new_n497), .B2(new_n498), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n510), .C1(new_n444), .C2(new_n492), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT88), .B(G36gat), .Z(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G29gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(G29gat), .A2(G36gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n513), .A2(KEYINPUT90), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(KEYINPUT90), .B2(new_n513), .ZN(new_n519));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n522), .B(new_n523), .C1(new_n517), .C2(new_n516), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n513), .A2(new_n516), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n519), .A2(new_n524), .B1(new_n525), .B2(new_n522), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n529), .B1(new_n532), .B2(KEYINPUT91), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(G1gat), .B2(new_n530), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n526), .B2(new_n527), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n528), .A2(new_n538), .B1(new_n537), .B2(new_n526), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(KEYINPUT18), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(KEYINPUT18), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n526), .B(new_n537), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n540), .B(KEYINPUT13), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G169gat), .B(G197gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT12), .Z(new_n554));
  AND2_X1   g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n548), .A2(new_n554), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n505), .A2(new_n511), .A3(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G57gat), .B(G64gat), .Z(new_n559));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  INV_X1    g360(.A(G71gat), .ZN(new_n562));
  INV_X1    g361(.A(G78gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G71gat), .B(G78gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G127gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT21), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n535), .B(new_n536), .C1(new_n567), .C2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n572), .B(new_n574), .Z(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n210), .ZN(new_n577));
  XOR2_X1   g376(.A(G183gat), .B(G211gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n526), .A2(new_n527), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT95), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G99gat), .B(G106gat), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n592), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n588), .A2(new_n594), .A3(new_n590), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n528), .A2(new_n583), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  AND2_X1   g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n598), .A2(new_n526), .B1(KEYINPUT41), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT96), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n601), .B(new_n603), .Z(new_n604));
  XOR2_X1   g403(.A(G134gat), .B(G162gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT94), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n603), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(KEYINPUT97), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n582), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n596), .A2(new_n616), .A3(new_n567), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n567), .B1(new_n595), .B2(KEYINPUT98), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n596), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n619), .B2(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT99), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n622), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT100), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n622), .B(KEYINPUT101), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(new_n620), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n626), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n615), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n558), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(new_n313), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT102), .B(G1gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1324gat));
  INV_X1    g439(.A(KEYINPUT42), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n637), .A2(new_n500), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT16), .B(G8gat), .Z(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(G8gat), .B1(new_n637), .B2(new_n500), .ZN(new_n645));
  NOR2_X1   g444(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n646));
  MUX2_X1   g445(.A(KEYINPUT103), .B(new_n646), .S(new_n643), .Z(new_n647));
  AOI22_X1  g446(.A1(new_n644), .A2(new_n645), .B1(new_n642), .B2(new_n647), .ZN(G1325gat));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n485), .A2(new_n490), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n485), .B2(new_n490), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(G15gat), .B1(new_n637), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n488), .A2(new_n489), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(G15gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n637), .B2(new_n655), .ZN(G1326gat));
  NOR2_X1   g455(.A1(new_n637), .A2(new_n258), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT105), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT43), .B(G22gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  INV_X1    g459(.A(new_n614), .ZN(new_n661));
  INV_X1    g460(.A(new_n582), .ZN(new_n662));
  INV_X1    g461(.A(new_n635), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n558), .A2(new_n661), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n664), .A2(G29gat), .A3(new_n313), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT45), .Z(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n614), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n505), .A2(new_n511), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n455), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n444), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n661), .B1(new_n671), .B2(new_n504), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n667), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n557), .ZN(new_n675));
  NOR4_X1   g474(.A1(new_n674), .A2(new_n675), .A3(new_n582), .A4(new_n635), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G29gat), .B1(new_n677), .B2(new_n313), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n666), .A2(new_n678), .ZN(G1328gat));
  NOR3_X1   g478(.A1(new_n664), .A2(new_n500), .A3(new_n512), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT46), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n512), .B1(new_n677), .B2(new_n500), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(G1329gat));
  OAI21_X1  g482(.A(G43gat), .B1(new_n677), .B2(new_n652), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n654), .A2(G43gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n664), .B2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g486(.A(KEYINPUT48), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n664), .A2(G50gat), .A3(new_n258), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT106), .Z(new_n690));
  INV_X1    g489(.A(G50gat), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n676), .B2(new_n450), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n692), .A2(new_n688), .A3(new_n689), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(G1331gat));
  AND2_X1   g496(.A1(new_n441), .A2(new_n443), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n455), .B(new_n652), .C1(new_n698), .C2(new_n416), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n509), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n557), .A2(new_n663), .A3(new_n615), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(KEYINPUT108), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n303), .A2(new_n312), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g508(.A1(new_n705), .A2(new_n500), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n711));
  AND2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(G1333gat));
  OAI21_X1  g513(.A(new_n562), .B1(new_n705), .B2(new_n654), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n652), .A2(new_n562), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n706), .A2(KEYINPUT109), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT109), .B1(new_n706), .B2(new_n716), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n258), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(new_n563), .ZN(G1335gat));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  OAI211_X1 g522(.A(KEYINPUT111), .B(new_n661), .C1(new_n671), .C2(new_n504), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n557), .A2(new_n582), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n614), .B1(new_n699), .B2(new_n509), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(KEYINPUT111), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n723), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n672), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n731), .A2(KEYINPUT51), .A3(new_n725), .A4(new_n724), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n663), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n585), .A3(new_n707), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n725), .A2(new_n635), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n669), .A2(new_n673), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT110), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n669), .A2(new_n673), .A3(new_n739), .A4(new_n736), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n738), .A2(new_n707), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n734), .B1(new_n741), .B2(new_n585), .ZN(G1336gat));
  NOR2_X1   g541(.A1(new_n500), .A2(G92gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745));
  OAI21_X1  g544(.A(G92gat), .B1(new_n737), .B2(new_n500), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748));
  INV_X1    g547(.A(new_n500), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n738), .A2(new_n749), .A3(new_n740), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G92gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n744), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n748), .B1(new_n752), .B2(KEYINPUT52), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n750), .A2(G92gat), .B1(new_n733), .B2(new_n743), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n754), .A2(KEYINPUT112), .A3(new_n745), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n747), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g557(.A(KEYINPUT113), .B(new_n747), .C1(new_n753), .C2(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1337gat));
  INV_X1    g559(.A(new_n733), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(G99gat), .A3(new_n654), .ZN(new_n762));
  INV_X1    g561(.A(new_n652), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n738), .A2(new_n763), .A3(new_n740), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(G99gat), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT114), .ZN(G1338gat));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  OAI21_X1  g566(.A(G106gat), .B1(new_n737), .B2(new_n258), .ZN(new_n768));
  INV_X1    g567(.A(G106gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n450), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n767), .B(new_n768), .C1(new_n761), .C2(new_n770), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n738), .A2(new_n450), .A3(new_n740), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n772), .A2(new_n769), .B1(new_n761), .B2(new_n770), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n773), .A2(KEYINPUT115), .A3(KEYINPUT53), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT115), .B1(new_n773), .B2(KEYINPUT53), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(G1339gat));
  NOR2_X1   g575(.A1(new_n749), .A2(new_n313), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n620), .A2(new_n631), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n623), .A2(KEYINPUT54), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n620), .A2(new_n631), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n626), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT55), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n630), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n784), .A2(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n539), .A2(new_n540), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n544), .A2(new_n545), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n553), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n547), .A2(new_n554), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n661), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT116), .Z(new_n795));
  NAND3_X1  g594(.A1(new_n557), .A2(new_n787), .A3(new_n786), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n635), .A2(new_n791), .A3(new_n792), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n661), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n662), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n675), .A2(new_n636), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n778), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n499), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n262), .A3(new_n557), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n494), .B1(new_n799), .B2(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n777), .ZN(new_n805));
  OAI21_X1  g604(.A(G113gat), .B1(new_n805), .B2(new_n675), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(G1340gat));
  NAND3_X1  g608(.A1(new_n802), .A2(new_n263), .A3(new_n635), .ZN(new_n810));
  OAI21_X1  g609(.A(G120gat), .B1(new_n805), .B2(new_n663), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(G1341gat));
  INV_X1    g614(.A(G127gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n802), .A2(new_n816), .A3(new_n582), .ZN(new_n817));
  OAI21_X1  g616(.A(G127gat), .B1(new_n805), .B2(new_n662), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1342gat));
  INV_X1    g618(.A(G134gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n820), .A3(new_n661), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT56), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n802), .A2(new_n823), .A3(new_n820), .A4(new_n661), .ZN(new_n824));
  OAI21_X1  g623(.A(G134gat), .B1(new_n805), .B2(new_n614), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT119), .ZN(G1343gat));
  NOR2_X1   g626(.A1(new_n763), .A2(new_n258), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n801), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(G141gat), .B1(new_n829), .B2(new_n557), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n799), .A2(new_n800), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n450), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(KEYINPUT57), .A3(new_n450), .ZN(new_n835));
  AOI211_X1 g634(.A(new_n763), .B(new_n778), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n557), .A2(G141gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n830), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g638(.A(G148gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n829), .A2(new_n840), .A3(new_n635), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT59), .B(new_n840), .C1(new_n836), .C2(new_n635), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n662), .B1(new_n798), .B2(new_n794), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n800), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT57), .B1(new_n845), .B2(new_n450), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n835), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(new_n635), .A3(new_n652), .A4(new_n777), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n843), .B1(new_n849), .B2(G148gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n841), .B1(new_n842), .B2(new_n850), .ZN(G1345gat));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n210), .A3(new_n582), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n836), .A2(new_n582), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n210), .ZN(G1346gat));
  AOI21_X1  g653(.A(G162gat), .B1(new_n829), .B2(new_n661), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n614), .A2(new_n211), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n836), .B2(new_n856), .ZN(G1347gat));
  AOI21_X1  g656(.A(new_n707), .B1(new_n799), .B2(new_n800), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n499), .A2(KEYINPUT120), .A3(new_n749), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n499), .A2(new_n749), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(G169gat), .B1(new_n864), .B2(new_n557), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n749), .A2(new_n313), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT121), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n804), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n557), .A2(G169gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(G1348gat));
  INV_X1    g669(.A(new_n868), .ZN(new_n871));
  OAI21_X1  g670(.A(G176gat), .B1(new_n871), .B2(new_n663), .ZN(new_n872));
  INV_X1    g671(.A(G176gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n864), .A2(new_n873), .A3(new_n635), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1349gat));
  AOI21_X1  g674(.A(new_n329), .B1(new_n868), .B2(new_n582), .ZN(new_n876));
  INV_X1    g675(.A(new_n365), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n863), .A2(new_n877), .A3(new_n662), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(KEYINPUT122), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n879), .B(new_n881), .Z(G1350gat));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n330), .A3(new_n661), .ZN(new_n883));
  OAI21_X1  g682(.A(G190gat), .B1(new_n871), .B2(new_n614), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(KEYINPUT61), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(KEYINPUT61), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(G1351gat));
  AND2_X1   g686(.A1(new_n867), .A2(new_n652), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n833), .B(new_n258), .C1(new_n799), .C2(new_n800), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n557), .B(new_n888), .C1(new_n889), .C2(new_n846), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n848), .A2(KEYINPUT123), .A3(new_n557), .A4(new_n888), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(G197gat), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n858), .A2(new_n749), .A3(new_n828), .ZN(new_n895));
  INV_X1    g694(.A(G197gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n896), .A3(new_n557), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT124), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1352gat));
  INV_X1    g701(.A(G204gat), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n848), .A2(new_n888), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n635), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n663), .A2(G204gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n895), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n906), .A2(new_n907), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n911), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT126), .B1(new_n914), .B2(new_n905), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1353gat));
  NAND3_X1  g715(.A1(new_n895), .A2(new_n223), .A3(new_n582), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n904), .A2(new_n582), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT63), .B1(new_n918), .B2(G211gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n904), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n661), .B1(new_n904), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g723(.A(G218gat), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n895), .A2(new_n224), .A3(new_n661), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1355gat));
endmodule


